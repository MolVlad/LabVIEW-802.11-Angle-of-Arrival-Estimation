`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JZhOsrTFLyLkfKlyZ3K62Yf7O4Nz6Uvpi9yrHfQjx6OH6cAMnNPVLeNi6kVpzQPtJtt958fpBkBR
EpJFeGPk6Q==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KFJwGmX6/09xYSekA/Gg2c3H6r+B2yt9pcXhhTAaS1hX5UlBk5/uWKuSDvk4m9JwNSq86xnb1ucu
A8uTOA6HyZjdFQSfQdUHHnV5upQJ0tGvzyGCpuyNhaWqZ5H7TdWboorPhSGOujUIHp7udeknl8kc
KNTlW1cmdhzcHKTZFgM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qXXsf+JUiCBd7O0DLBq54sTG+bFjaTFdrSZuEfA5r/TLPzvZG3HpmHlmfn2/3dQAb+CgC0nUCvqG
+sEMIEEYiVWFp9yxLbIB9TWyvmsWC7wB94hFrlaGnULm46wtldy8G0W40vZG5oLFvUJ3tsurEgwr
U6zfXChZCT6fXts/doyY6HgHXWBHhInaiWU7zfRt9d5hMczekZ9ulWXgGQyu7O3qEgPKTgYiY5dC
lch5vYAOGvj+gwbiMbvhYMZxWtCsySlDBNKNWcpd0i6KLl1pOojdrUS1CtGrsxOwTXOPYyM1GqGh
3OG+xBcWHqZLALLj683y4PtjYMzjE/HTbMzxIg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gwEBzBiArlnmssU81jPGrNg8ORvA6bEpMaXvEHPgHNWqMF+EConzmJMDay20BA5u0UXglin7xA3/
X3JzNTS7AHZmTdGwR0loWQ6cmNP80ixJzX05PY0YoI/O6NxnNelR9lCj9dJXgC1nGkRJckAPFQ3I
GoOfLO0yaRG80NioVU5N1LWXLLUp2fw4gr5KnsHUl9RJOnTeuCzBhWMfDYt4PmE5TsY7+zBHaq0v
i06mDT03IYqXTCDgW9EvjImUoFyEESTMQXEibqHPfTQWNINtCU3mDnNu8PepRFHqUPsV4guR1oFB
+H7ZAIODlJCR2d5kGH2wwK2ACt037de8BYgzgQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Le7hg8IYsU8S818FN2SF9arBIIs6ZtoPuSbpQNlxOf2uNp5xfjkAasaOgLstEqit3TkaPGyYYLUS
yqBV7mgIFiopNOkgEtUYNmKDG5Q+owdbHsC0GD9parKzO634ZGUHrCAznBQ9GqBHp9q8qGLPT1TH
NCceCnqI65PLDfhlVPlv7xCu7c7f8KvqNGIy12hikQrbKpf4EYw2GFTdXma50Dj90MpBQpFdhIKk
wlZ3fRwbodN7qmZuH1vOnfpkDT+1V96B6zrajuo3e+j1QctslR8+uMUU8nATLS8GIYCxyfKNSDzr
qj4A80RqaNp7gSqekF5U8I7r7/QBHF2KZj47cQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dlA6S4LJnZ8SAIayp76Lenf24FfZqNdir0trQ/N/m+U8IUUxbAsRnB/3sPESnvXJN1CMsGTGvdvp
fo8k/i4ds/+pwzf0N3BWhbOgQ6wCmE9edMU3jFTuiDLDdfbKdHbWvhTk/r3prEslrFwG3Gk7+8YO
ekVojNEfgIv+0dF6M24=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
orJ8OGcpFqDg+Kz8pot9VmTSng1uovp4yzV3b9VvRkIg4UN5cyXGqqvCdJewDjq9Nk6qbobxGLNd
eR9/Cuco8uZXfSiO3W2X+Z2ZMeIoC6PQRaqoMY8iENuwgt/KCm2xv6j94s/FNsNok0Pcf0Ld1lQJ
ZHpu/MyYgcOQW6BnWliecrfU9lBVw7dMB0ozU6rKDwZwCl3yWT2h7nuayk977HTAxAgxWqjPqvcp
1Wdm0cilkUk+ifH9ie0wyZA/VDmvzmNbuBffsGYKFwa0BK8xmcj/YKwWyp0JSgXT6ky5VWp6Ia1z
YRyqs8XldNyDG0nEKvtJn5OZItBJrbJb1w3ZVw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23056)
`protect data_block
TA34/xCIuB0XZg4Rj7XN743N7isGOyac+EJoa2E/Vi8hvxqrFT5A9ZlfOdImDcH/M1Dvj+wTnYLs
xjDQh44y5MsLipWbQEvcFU/d12tBeIr28O041B0C+Jv6dG1FPIeS3Y6aD5mfM4ODVS3Pg6bXwkQM
rciDpkfTKLgGICOAs3dJm6kIJCTJb7hGqmFk5EZwOLx+emDhGfJa6bXUvZy/zkm+uVL1xgsqpON3
ul+KR/1ld7Adj7jcseLgAhKIeV3EsQ2OAmA8ytcaPtVrAHzNeOLkQ2cohqR30biyiJwe3C8b6r3D
LNORFOevbxCNXHV0JQ1LZbo2NJn947iwbgW6TisMrfuEvb24jpb73GVE6DKZTyJ1c/TR9DXe3L0a
aZiWt9vihqD8N/+R+hLiZAS7u4GFoDu5EouYjOWOqgAkVWu1GN9aHx9BY8hEb133HYj+YBxK5Rhn
K2WQEfCHmB9qStruIzZgsHe8b3zU3QkjcRcVc4BirRB0Z6ApkO568YG04d4B+VhaX5/756l1gCZP
mJksZEHW7WaXLOIhyMSUOSVoDMuEaRmPn1ro/wDPdH3Li3vazWbAvCxOEQmKbHSYg1tb60dm4Euh
T85qKd+KDuzgPqK3X4onZfCW1lon1z8W4dA40Sg7GdcDdUkPEWX2WEuAP0R2mF0guKZOmCxxUNoJ
Bzmb34QV0iYG5pz3IQQD6wKE1EzvKmP1xVnc4erXD2IN4O9Lkfaen/oo+NKG6fyNgYFBpyxotSas
INJ6BSC+9tRG01jrX7kzRDV9Q0rbzErrBMA0997SZG6lfX3mKGqO3f3hBqjPEhkNcEtXPdyRrUGd
CIkBQ8TeBgoZPsjw4RSh1kTpw6AniRrpvsI7tUod+uUkF/h/VYDM9RQEpIKrpG9P1vG5VLzH7NiI
F4grYRBzMMb42/5ROej37WAQ6rv0P7U3bMZuS6KO0aD4gj/mn0tVe/iBNV2xOixgOcIa2wiLt/hh
1BabBaClbfnzL4F2wWSsFb3U1TajVK7FqDjHqVJz8ziYMaBRVRCe2VsSLFtgPiHggqrWED7jH6d3
+vQw/VPHxxyKg/GQwnvhLKrKbZESNQcoZIAGxxMeA3xvUkMAEZEicegkSkmePCrpOXBjOt0k36IV
6KQVt0ama4nxkP2aB8bg5CIctQbm187UDxZ5ESNmljz2v9AIH1UaWEQ0tYRCiqDkHxjY4zd0yNtl
vZMdQfSqPr4/qAim+/SZIQg9/pub+R5FxKbNSTlKTNje5oHaOrpQLxAzzV/s95Rq2mNve5M4tnId
LHxmVujVNN1pAzrN7OFbwSErLnifDqwvY9v0HZmemWEDloAMLHp0s6/kAglnlry8YW+NeoDW1Teh
ivugS1BgWxK+2h50jbGECpDWkrIYr/hY+3dqKqm+jlN4Ai4u+ysOzV13M5TKxYpnoHDkaKfsAN5P
7pwvl6YcSd6XEMXI3J2N1ENrI0Eqo1YpaFvWHrPD+C29FVJ+iMWGqJSlOmBYAuTMA0xNPJlYLPwU
vk20TnpCRH95TczmCpn+Bxp4c2MsHdsP2cc25xCGE5gUyFj659tEsHR2iop/Lnxq3fxvzefivVfq
iLJTe1ZmptpXatmIrHMcEwUS1RiSDy7E2sZcg9K3qdWaDcwyCge8MCyumd7S/cPytuAWrPTANOtN
2zVrVNk9T2AIbShjp86yi74Q+iHnEFw9+DcJrcnEDNuhuqNNS5UGTPldTuN+NEuM5cmtM9rt3Vfw
SF5o/JH3hEHo2xDRvfV9MAxLQ5rdDct/jqCrVQcgqXjs2ueLeGeczwrbunbVO9klB5AzYc9DRMe0
NK8UbFuYyofcy2RCQYYyhDdLGAhBWB5me9rQCw0mk+s4HgYDry0i5t/mOEJB+22kriWZVPkaNMHo
/m6AZ+jpziiWdqFVITt8FNfEHhxcHhl4qh9Rrt9CoSdPIilRLqERwnHJZ2gM86l0NOh21ZPMBi0x
8/tWyZBuWrXQO4YjOT7quW121744hOPfEzg+fdXM+VndtHMTZwCinO1soiJnFdKUK4bFxyyhMdCE
7hzk+kkSAZeLfEopTa1t+NldPOBsdvjzo0u6NFVr668Kodr93NxQRgrUbOfJ6xu3Xf2Iqd7BOEr0
oxzRKCV7SAJHAq9M7PBjuXtidtQSUvL0NpnYhUUfQsBgLq+3K9IEtSknQsrR/sPDW+hA1ZzKjK1X
Hl67elL0Km0TUH4lftOnNQKVaNXduqqEyayiyhjQvUf89qQB9G6FvBV/Lz08BdlgcNFd2chrXMqt
XMPT/zbGIavBI8mDroEvqYYbRkZfRdrygriNuo6bkB/eKqAlt9ZXtln3T1XdTP0XAVLyu/jIXwtD
et2B2AmqyClWJyGH2W1sgX5hmd+CUKjE3USVYLWwgBc5sSnPc/EvlOt7pktsv+usogVihB+Kfgo8
pwDsMbqlTO5kj7i/8aUi7CkIhgZxxnL9mQA6uPPOldaapkwGVV+FduEreTVbbgbRh77lmNm8zusF
UuL+qNPxmZ6z6ZOO80TtdMNqENfX0Obudt2YJaqlK/bC1Y04sRXSmKTs38BiPRT96Pago4Jsmczq
a+rf2zcwT7Zz2GIonLyiFIaUB8tmuOhQH0obgIX9LBd8DpcJdHTYid76ga5EtMlwdXqSqNBbV/mY
F1yC7RjrKewWWzwEJHIyGrck178u9Rk9VCa4/idyX8Zd1zPSBCYr6z8fyhBqHp0TgW6/tblK9MJv
ZUka9yL8ynJw33Qak0oU8XtDngiXQzgP7TSPsRVDHUBXOn0jTmFxvPTZDLoqPf4OXVPNQbrT8ml8
RC8772qhtxLCR0RM6V7uDzjh57WFO63xY2+oO0Ls/dqX6xlos699n0Es4BVeeyZrrQLk9C0fhwXR
klUfoI/vT+dHHTS55PN8G53i7Y3xUBQkr/JpuRCbASLF8TYP97k3dX67JiIPovTMaBcRrGT7HZdQ
xlM66YqgZVLcvaxI621/s6yFzKChxSBD1VaNG1syOjnT5M3r3yjiHQ5IOHHmWTd5ozT+kWcySVE8
3QKQbfGl/FwRkHwnrh0YI0RPtDp4rlJzSOEsBlVqoahAcRTq1YJqSpFMnNqI/qpRZdg813E4x9ai
hMLWNZqi4wF8S8sIhb5SJ6nWTDodL52eH/Zhz7BV5JkWbT1Esf24sbQ2GBiWKqD2a9WdPHzMV5RN
r60JR35N9cTfwDhKSUO/AAUJdZsvks9LjOxWqShck3vbjWg8yUcwuazTifTXmvtealZkKAbRUb2Z
jKK9xp2UrXMR2KqdXW2IHaAtkVwzk8tI0zId0U9Pig99AYPYVd+4Cu2snMlBiyyTo09btsV8ItJ/
uhsqt0I9bYiE3l3477KwLaa0hcMyCuCNNUr7kJC97HWCvASUG1J/wKjIHLSd7d9uI9eeuQvcN6en
orwyp2qKdnT+BFXwMYdU4UsJ+Usdwf7xMZIUFr+mpLyoJ0QV8yYuHS95HzkGe2+iGu+K/Kqc9YNw
vS79kT4fMivt7vNnFIgoz19l1SL1aBCzJiUpah9j/jJJUrceSulHe6huekWbSGyQBB9dT/D0CgWv
qInBkseljPozQfsbTYcSs8BWmBXjtWEAcwoE60Z02XMsAOf4eZsyrslpGoMGFr9X1BrZLlyT/fcG
b0yby0zvhqhZsDfrOeuXOwvGIBVUobYi+b9ys4lcXtlN9vmeqsgh972Rhq0wnJZuXTM3v5bYmA9u
SMeqiB+77HIH5aW7NW6mEJ6S/vhpgNcmP/o3XSmLOK71hv/zqKodf6kZJs6e8NzUH5nHmRJzaP4e
PHh3pvx28/bWURlhVOkb4LIj/CgFsyt3W5PTu4H19PuOVtVGS3hwHXw/r1d3oZ2VrmgyHH0LA2A4
b/qEO2NzS9qvrLJD9CTJgbiovbn3YkFS2rh6CsOks7I1jj8Q/ljDwsVki+H/9gMy/Pehs2pZrqPv
cz83Y+siMCNK4p11kdhPcs4QLxjnwFXs4jSf68FJOJ3dCXAC4sdYFvv+Q0i/9RuVT5REeg0RlE3c
mWzucvNCN7VGAuG5KFRbb9188GLdDEH20t4WdUSdNmnVaFP7F7ibvl2QcZsA6JAfCnwgqS75Finl
Tev0pXIavVRwufG3NkUScYrkKfCDVmE/PLZVkDsFdOP2xOglMg82tLv9zWuAPakIk8kZGdIyarw0
vfO9ilMtmXLNSNwIZ2caKNI+03wFxw2uBU2V70piA8AVVZ68MFcUNXozJLF3jxiG4QVwrrlbJuCB
3xndyMPJ7yUCyhVSI9p356A0MaYxL9urDMKPdXdgjY5xHUSBjGBg4ATUSM/vLTqWz+/qmYh0s/jt
93PpO4t3oOZKRERBk5aahSaeBdVoy0MG2qljd/kczPf3dsvgDpK2e2mb/rvYn0oovikdg4CWojrX
oPyLBQY//ShCjB9kjk4vPWK21w9FnbL0FPG839mXaPAcozxL5PgMkWLxns8FO5nbCSZKNf+cHgoR
ELrArWAXVvmwGiJ3rHtHAMmq89Qlk6iBpPfFgs20c5+nS6Mcx7zOXF3J+8Jh3ipa764SfQDcN6dD
ZltyIRKoQJrzgURZRVPo6IzqGt7KNSPzy1Z5WBnBYUIkAVa0fcNFyEdMiBHl6su64X68z0rV0F9b
HnepSyFuLB14rbUYSf2EKJpzAUzxQIjqCJ+8hRAiN3JmRysn3U95bE9snVi0xfMdR5Jx7kkPYaZC
AVGk7nhFGtXTADkD2yPgzut/f/g2iF+Y/03k4UqJKidPcD6q8z3T/EOUqD/pfPBU+B8DvoDa6PDg
ZCxPU6rl/qR/ejy7np36v47VIEg26knTczCYjKG7lmw9tRxbfd+KDA44SZGMHDlaKj5vPJZ/sk1f
wPTi0+YCkjJNebN3GBaYSaGUTZCGPfbScom2R+Ds4yxOtnjOrAHrh7rI22gDTGP0UaeRQi5i5CrJ
CZ3nIlXSTGgmsmnlsJY1YLtYja7Cz3EW6Pgy46wVLL/TMcqRVoN7oAAKyDX0g4c8NwnIaW1QRX5L
/k+zrXsaXl8OZOmGkVGRRXn/BBi15xdk78rKV3047OCWUlaxej1FHHwACsdJYDZX7rIcC7Pn3xvT
lepQ5Gj6mqWGzV9OY9oSpj9Ec5KSx0jFYK7QBgYmgqR2ceuP6zEM4QbfadLu6zlTT793XDwNRy3O
YJWtRQ/hEViGZseMKRjjVB+eW3a1qAVJ/qF58aeqiHFFfK9ZZlkxZtbgyRmcWrIqQkUBb8mFDea0
ojHpBLQ3w6xmZw4+4IxvLM2u807gUKLy822NlcDXWSf9eMR16TY6Gyao/QE2tniLu8DU0frgfQqM
BKnwY8fPvaZW+xgDz3KU2hG2QiUvmoqyJDQd6ZUNamT65d24tI3RMcHrw9+CXxzDUbZqRJdYyv1f
fP1a6AmRDcVUHXB/JAtZO6aSZluQuIoKhipV1Cu3e7Ua/Z53xgvsN/5um0V6jowcXgnzqTB5szFP
+ZfoOl2XXUovXWp+ZxnP8ypLZvtYY+g5UrOzjUG7v2O5PCb+BZ+/fugrEcwL6mA8AAM1lVLPF4M/
zFaEgvC4xKCdAIzs90axwv1MZnQHgw5Op11C8fmkd2Cqm2xG6/YpH31XoPlcPIpCJ6lhB5LnZDBH
j0582StPNWcqNz61x1jav0F1O7aqCKwMVsaIq5lkAsXTBWZ18xmj2xKAmX3GEDelQjZ7rP9KgmlU
M0hlg8nVEOauBa6fjATlmM4InUJZvtz3bKhHnMCHQdz/ksf3XKKZ/rUobTrwVDaeCjJxQv6vd4t4
nXiKB5N0TTDi2RZ8ii0vu7jqIyTFFnmPOTAOysXN8e4E1L/c9oXQIyi9Fi1RHfpbqD+Xsq+HlTcn
L03CiDxv+S9M0m0GpMTg5zpYynpHI/8DaFaOeXt+MXYvdMpL2b60AhP5gK1LW7m4C5KcB7qXg9aH
GwKMCuf1Fo8kHJRTgXlK89U+fyjB12NA+XQzCodJRHDm4JPx3fsDifZjDJ+KRWP21HLeZkd7Pwfh
nWFMYSqQFO1wLPX+Sqgbd314ssyDotvmPjIrcWdUeTJaP39QYZRk9mtY9j18d+DXWTuqq+dSkceI
Ik0h+uO2VCbHTS9BP+tASoic83qhwD9C3qz7cKAUtdlQx7Fa4gxYA+1vAiS7UdsfPV8lMMu+G0/Z
r7o4qlSA57tY7v36UvNk9u4F6CXFDEpyxfn7zQEEJ57b4EFGZCzqVkfhWZX8zxQjkSUPDv37Wfti
VYCT+99DbEKN+ddRRAopyWqJRt3QZoHXb4uvts+zTOwbCKRF/DI4by48iwFvCmvELHLYX/nGNu81
592867g7odLFL4DmWeEvPFJ/HzlfYj2hPRY/bLTH9qzIzZLSlynONaKZ1xxtTusrqAfxdG/RA8wr
wzYkU6c67bhUqZrV0BbnQVU1k+5hXjXDkfg0eJwbwvP/rxzS2M+Z4XTo2JkIzpcRjrNXkBNcyhSC
/z208u0xz+2xqZ+eAjar4OwtYmToq01yyNm/ChXz2xQ+V4lsJqkLltAZfbgHk5ZJT/fJueLBYYQ1
b9q46Jq97pTAPzSHnQiwJ7M/Ia5BH/0zweAwHYm3vKPUyuR4ag9eVX864lTxiCR6GEFRIzePp+QA
2btX5+pCDwwHU/ElM9Jze+fu3ZB8OvO5pwF2HcLj1sPy4q7aTAMgxim7HjcgvBdHR0ZEhcpTM32w
+0JCl1ehlIDsPpUZr7UMMIvm5zfzfNSKe8kz7BmIXCcsBOEktHpXZcAxjI+yE0xvfQNCerqRts+T
NCgsj6HJJCWdm3uGHZeLbtikrASHN1iiq5kuZ5o1mt4qb27VQ8kmSp5Bayia4r/QtUxzxU1lyTIg
3OcUCmiVzDt2HmpHBnfHWrrKR5KbtgHo+QipuSrezcXEPgU3BrqY+h40/plllG8Ltnlhe0xLrlLc
8T/PXM1d9u9D+2Zy3lqJ5cDwtpGT/rj2t4GNBNJ00OBGW2d2wWSzuDNQUHgs/euu62fPYyH5lr+t
R+KCFghDDPJvtw5Qti5YXhkUsTcY1UO7gS26YJufBYYNJZlGdzSfYVFzNCA6nsc2oF6j8ftlrUfz
F5fnpJGVcr+keCML/TgxNoGLkUfxwgCOZGdsnrKfUIFwmntJDm6pecsclEPBdX6HVn6ZL6SQkfHu
clT0c4o7pIcm7pYqHviUQwn37gpvuIzqfByGyP5/P62JpTqRsxHHCNb3+Ff/Vomq7+tajIKUjnbQ
pnSRXg0wXTHKIZ9luttpfxvvUkx9GYpW+Bm8DAYWfa49WO/QgWTZzOFmrlaZuF3TsoYZl4bNp0qw
y31pRyZl0Y9niSrwoA94Mj+MhBcgpG9Tr8pqxmXIamKVWctlu2Xk8UC5j7WefrzE790yUDK53IjR
DvwYz0dcquXX3kxsmZrBPPhsLaNYQPhReZSiq/ALgni4ZK07Q4e8CywTKQrtgbLfT19EttdG+K39
SaukGCX4gPaUwGDIHT7I6t5W1t+O7Qyl7McimaFhu5qMylrPRqFCJwWNh6FV3STV5JlXQ+MwcSeJ
oQB/EEwWaoHaumZsVD0TSCVzzCbJXmJCSsvidTifdAhMaOKlCWRBIJ9xUNQYxHmm8T7i2m5QQSkV
Xcr4fs7tq2EosyUJGzEjf0VnOenEmm779eigDLqgHxl+cn3a5ke2OTPEfIcB+SzTzDkfErc3yfRp
TNqlEjI3HMnyemfuPjcBB9FGe1ME5OHVFdZba9B+J85NBplbRzqvXm9z5QTLuvb+8btr5s+VHbh6
YJBhZ3UdU5Pht3YPA1WIx6yCd0Entn4/8V4nZA2ukmgv+CPnhlD0lhsbj7BGXdzNF5y3MMTUAm0o
4og1+X5nW6797ghPJJwmeeSSC1sCI7uqVolgfdSzfCF+PX8C/oJb+9xSBRJkKoQRMv7T/zzSrw6/
yd1eRtp+aK9z4sMdojGAxDkz1TC781izHDsCEKoSsSy3sgYT3jMBuv65GxR1WI8c73y6oke9BqyQ
8W2/rY4Adf4zvwaulkChPOJZU+vR+BbF5YHxRkjVjgR6zRzF3f+JWJD96fxl5vq2xKHRWxLEnpYV
fMDREBO8Y/eQB6UBE10kox9eyU0hdhxQzSQvhTs9SjBT7dyMTLGS1HVN7IiU+KtsaLpZpObC9P6S
+IvYcRWGk9XvGFA074daNl7UvO7ZqC78Pg7EQJqFRrjGGkLf2yWxCkxn1hyibyUlEbrXB9TVX5gJ
VeOFWdgpIwufSgC/EtJ4SlGyOYueAao0eJJs8nG1gDYJX2OWQwISfk4YVVKVb/1NzMmJnSXBY29D
yYP6B5eg6GJAc6+iQ62BmDep7QJ7kZYBtJ4iEuiB2CkTFy11Wqc2ojFOWjHvDzaKQwNR2t1x6yAP
5l9XmBOqwiyBYk8KM9W9TRTiRw/m1bVNIsKViGU/9wrLj+mhdlNRcmmK3rW80ESzlg7rCFV3zJX6
lL4Jmr7ql3wWw8q4SSBVsQ22dr6Y59Taf+mFeFP8YFhvEARPlhIWc/beNg7FQkvSJoF0rw7Bo1K3
e7LDErjfOdyu1/+dIuCnuPVu73UVq9Kkm/ESJagk0f4fENZH6rgq1GbK2OYWEHXleXVMcQ5u5ix6
NqhENnigN+/wvoV6y3/8Py8xhns+k5l4tW41kHyDYd9Cb2npCCAWRFnDERsnP2Xp6LFYiz8WvqRw
CndMg0fqI3aewsyv8g/PtwfGlEdGyR2BQOCkQmE2BiIxNGt85N3R7vSPJ6oUabjTpuN1zXPjNEl5
SwTf2p6AQ80HMMznJrk8R7ypiE7oO83Mgm16dP/f7Pue4J/wI9UVE3sjjlrnRTT6otLfjbcRmcbb
twNDgeKddhYcqiYlKhU0KzHlX0+fT77jWll5gVJLzDTWbtSPgZs4KwSPWL08eamD7t3QBX5cKcxw
zUD6Emt4dAdnXsr1WiHQD5cTXGW3hDijqyaZLqLjkaX2h5d3Q2uBdl3S/QPWQCSbU/OfMuspZv1q
yPVecMVJWnPKKsIK/kx6l8NeIG9pZPbvjs2gy0cmKxwlJlkjMQP8jJEfI0fcHY5YoZii1jdJ6G79
bQ+Yht01ZBlzneMoMveOwetQwvAzf5znV32ck+xg+FFPztZG7wy27kWkiLv8z+zo9BQV960HOa76
IC8VL5eiY0NESak1i40+Dkf0h6zUCUdy/cil6O4w7WEWhHs7mru3a3ZZYBniz9+4ARcMiApy7afl
lGHVpC46HaS0+4ubKbZvmpr0fajOvmaSxVaLRcfquKWamC6KAxyIFGQucAwSy0f1l8Dd+w6C9k+x
L32/iyfXL2Uw8uRkBnJ0u+C647CXHJXDC+YClNQV+YIUsguKjhNYchMss41GougwCS0K/zgIKFzv
kdipZzePsN0mj17DRROmgr2xoFa0o+uCKubt5Ux8CwXruTuxUGJN9GsdJ6T4IwTpBX5XkwA/CoaW
1BhiS8zyiUO/YO7Mo1eiUcI/TOBuLPSTYrZzTSs1lHVE2ZuAK1lfIpuc6ea9PP6dl2dMSeZo3i5j
nzmVd9bv0yml6D5XqAtsUqLLXDaA6xXEjiIzT9YB88pEQDm2HucUBSr2f9J2X80SZ+bTg0GD0qhK
Bujdvl7OvxpyEZttnIuqYK5aDKFO791CqWEjVHkUhkAv+k/vlk4WSG/7fzIZyJolJAsepRFOQJjf
LZqaQ1fFnmGxitpk00xvaFaGwyeEdphRrSfDvME9RntlGvomDJ28/++hZVQgLKTCZFRnAcX0kSFg
cLrNujMbb0M09htfNZkn6WEFTrM5Gjl7nh72jYipVw4sDkwibH4D2jiKW/wvJXwYVThURsMEdieG
LC0xSuTjUzczvaapgPtCsilo+RVjDGr6REJFuyFnsWWLzbRqS7/D20z3AQxsKebuVGPnjzVTU47j
KxNzJ/A28PG3b9gS85bdnQTYq9LPXP46nKeCnTnxWnXBat2RChg7Z5w00FrHAY51r3RSOgqFGaLq
dRjUBzBJxtzg0n+QGkY0JWabvSlvuDCnc4iihBebmb3MzFiPuALexv7BeITz+7A4THDytJiuZ+DD
YRWYEZF3bDK85D3gVV1oXcKDd7jhWPJwntkxLG8S/M8Nbsxmp1HRsx9QdzbiKVFC07DSE7JcQkvV
ZW7pBzKkEfdw2fUGS5tdS5H66UkwTgVhSUDYes08GAlEJStDnPTYrnNg2Z70adGzUxlDoHGwl37J
ZYaQdF8JB4FtRuJfubIzWaMR0uXyqc4hWhSNN4sb0b5U0eV4RCO3LmTZxlU/ykZN2avbKzL968tj
feLUdqsrhVmwShcHVzzxRhYLq/gjsu/9PVzEXARKEue6UkOIJjl5iMPjM9222qKfXwWL31pZ/mAi
SW/vAhOyZm2kRlerVu03e/lIu/53zYq8v9vG73m2XftTmWXJ9mJomloD4cDBzTH2QqooYcOGfYB/
O7zm0M74zRb3w9LslZWuh3wIfTRa+0yZ0yvmf11uqT8jKXtfWrUd5qwmBtbLiG4r9/MuVVdaD5cY
r9LHRY4wO8UXCZWImoPc2yzDLsUsEXvbOYjHf1ZRdDPCoKYsRO8V9FYeg14R0bcIe5uTuWzDU3NK
QH3dJ/ED5uf01M/Ot9AlqOMAjJbcv7MlpMLKpJVbA9gnUR8i0L6GCVyJz+9OjzfRa1iNCVqxGSGa
UzdrIJcx1kat96WrNW7qCvLOaz2j+auUXnFocfbr0wPium6gNchsGa6vHgbRxMsmdsnACy6Jbjxm
5lV8qlEHfSFx4hSYt7cQRjQy2Ixw9RM9zuhDZZR+UBzcUDutD2+3Jlu1Q5ePo+0mpI9pqWwpZS7w
e6tc96Es9U8MlGiirafaU9/YwmBKFV0qV5DOZIxlst32FoIJ1ntCSJIJE7SXk+SwvdoAN1e1Ki+T
wuM5XyLcQs88zV1UNZ8GWWO/6pGcgqlzCjfVhJhQ0Sdb0LfwM8KuK0Zy+C4wFLlbOJL7GUtGoUMI
niL+YopZDcB4VvXb1leAyGGsxYbpXzoya3QB66bNcFbR2bCKBrFUob66DQsqF17yzoSTA1qGdrZT
30NDUwGSA8slSH/nOM7qZZe8w/+MNJuLzxa9H197AlBziHUrliTJNGR4f/7w27D5c3y7LQ3yMV4d
WFbyc3GG/FABjF9exvKJdzosno2drXCSalP918fNCM3tzYjzEngnRgjHogbE4T89Jn1TnFMD4BgM
3tYApP8jWEYDcUzExA2VyRmrJ4Y9weBfOrhRJVD8zKR+ouVGdaHg1UFpCJk4NTiGZflj/hljFLc7
tKiYNel5MkdzUuDInDOfCDsUCWylPL0oyZgu8mtVBlju7JC+O1F2hCGrl5srOmR6dPPvrt37zs4D
w4Nnum2+WfnPSNQZX4zLy/lEH4AuRchE4uB6Vhqs8U+fx8YgUUvyTA5NrQ9InZgUAaZWLQtL14fJ
J9wMiPG/ttUag/8U/Usp/SRrd/x6a4XLim/OmyjnHuD/lDKBouhu/hgCAQnkLWWV7xiEJQ+6bRZ6
pYvL/DnvNZtqwbqL8pNqsNL7xRT4Tl9fz+vt03wMt/lTy3gALVSXhvDxM132SxNBGePr9IiR82Z3
RX2iObPHERqakplydWQGyOJwUOMjT+PT+sdcxsK9tkc2WiBVhWx2oO8Spuv6aDgVFjAoHSpLAPNG
84ucIT2xnQ4+c3sPlGG9hxw4CfL+ZNG+u8lR6EwYKoOBogW/fhVcBsVCIp8OOl2cgCTKKMgwJmsK
wYIRLXPxnN4chXj52u6MtuACqmRzuy6KpW6eCMsLucnxiZKMMkE5OcUZBS1zariIuwA02jGJS3NZ
7kKLXjyqh8bRFbcPLD2qBoTuUm/BJOnB4LJG0gKuhX2tnc7mdyG3mMy+I40NuJlCpX1PpK5w74tQ
qj97GtA35bJ9TkGn1FN9Ax+DBHo/l59oI1L3DvC0zd0zONTvdGsdPaCyCJ0iyms0iqx5hVXs6d4p
CSE4XbYO96JcwE+gYhEkA7ZLsYBlfvk8eT1fk70iXuJuRLZ5/Ol6rl0PrHQMPVIv0d4F9K2i1Rdt
pm3+NiWG+JpIxHfgj1v/BExEuU5q0Od8dHolFStx2gQdSlmvDhxf9GQOpzlewyZDrpa7z0XvJorb
MynzOOOAeHeH+0tjIJtzxEcEVReBmx/Wh0AZrFQ7oVr6HX80uD4Yd9iPqONv9CpAwpbSKBzol1yT
S1ReYdksgM+HQErbZ5XDNcqbzGHkpRP4h4hxlj3iRYPRw0bqRZOxx0pXZO0OCG7o8Ytd5mc7ACMO
8v2/8c0iSFvfZIOWWZqu9uRyJlC8jILkdiCST6xYEUNVsejLcULHV0xGwcQDoAjB7mZK47lxLKcB
jhVyBIMVo4qmIcNrg6v7hJGP51qm3bCEpl1m5g9wo9MpWm30vOh+oZSIUtTRH881cAg4DLpUfeE8
/9u7a6oBchbAe1/17ksupurGbC9Fm+wYbIJk8RIu5EW9/+ckZKrhOmoiy+0bbD4vnWeNLBZTc0eq
063WXrJPktX2eMThlzp8gZDr074ZrDCzMesPQ/gRAALdpZwIiBrjqW69Rv5IESKSU11DPspj/Meo
XGj5t3YRgNFKoOgJLS18VKKUbvhCh9mbcb4lWTFJXabMHRM68p1nKK9++VXdEuUxlETgbUYA2dNg
Q9wHBu/XuGv7J3l6xwAH5pEy5IPil6GvnZrFcxhbpmFOg0o/SBUpnBl8/lfOnzpRIZofmcoVStQP
qPK89ljsRK5H5PgDOwIBZeg1cES+HxTsUi2JWIKsp+MIZOoKuv8xGVLDfASIBuZ9wYWAIx9Tcqsr
u9K9nz7uXxTTJoEi5I4jfbb/PtvmT2Cl/+r6wR5yc+lc3jBPkIXLObdmKNVwC1+JeTg9EkbNdtnX
v1W3mRkbQidHTeQxt+oCRx2xbB0Jmjj/sjQyJ8cBFVOqh1gluMCqjMt0POtctl8W3smdwG7/wpoS
aGkSKX6cOFQevOfTBeSq2APU7iPCtzx2qU42LkhdIafXxpk7kM3WRauVnA6lzJgewxU+lBfm1oaU
3H7dgRJDi4lq3zmEHgOaismZRAmFwrUuB8pvaGy+w8s+uF9GFO/Cp7/laP5dFFF7fMoTwuZZmPnP
d+acAh1ZIuBfoik0KQXwy6xdAPvdjMSAZYSa+jUu8/zQ0BiMO0xbjw0NknwEk9C3WWSyhlmaBFF/
1iyzpmGNiT/hebj0VrcE6OiYJMEC0R01YiwxdUFbtm7W+wbPA+iyzNnjeYzEtNblllLAIvsjDukT
Ji86CsfKqeG1/ZiIalKwYfjm4ntMTyzrl/xpY4YyMuf6+UVZp1qz9rI4UST32RledRhtin2Xl66Q
C9hEYc7l36YysxYUscj4ZMr8V1/Nva28ecEWG2nvm4QlMcm+78nRQXhYQeeWJbrT15vIfrPz9Slb
Gm0GYC/jxoEL1qwO+8cE1ha1MKXDsh/qbCKo4WRk2mUyyLsBH7tnL6eHz70ut4GFGIPWrUNnTrqW
8GZaoFJjxUeKRhVKXft9KVmNnS6YG6yTd1vrwLCUoCXr9XIOw45oSO6+32xVppuJ/CZ8Sj31ls+U
1VwRESayCpuxRfVIjYZoDD0HNWT0i4AcZoZFlC+S9ltTFCbyyw/mrQ+JM4aY1fIkMAbQevWK2UVS
aBRhDNL9ArMdUbuBx5p+c9/kOP7p/esi1t4+B1IAF9F7+LQSoZFfOmfS9Kw2ylzVETj6O/867ZH/
12E1fniPzWwB1brn8WLJBJZI9kkPOzwDw2DJKrm3Xde2qJy27nlll+GKYyCULzssDD4vU9rOLLpk
uKVWpVS8og+YJCZh1JfnJOMhHRO7V+QffzwOd4ioLcbqndNOVcCHKVpoRtUjzhwWq62/QpTbc/BI
OKNfsICYtGqiqZXJb5t4n/PzLQnwuTvh7i+sn+Q3QA2QkEDm0/yB9w9pBAYEhKwGpQrK4zJIGlpd
z3mENJub/NqsoAWIb+DIL5ViM0SNJGVMId6T93WfLzkXWpSYUC0FPT4eTEG6JAO4ifzu3MtCBgq8
vI08+VgI/AG7NGCQne/nMPEZYDrbtY8z3MPwOjqLNF0sbZtTVf1mSQ8kz8n1DS9E/Tmj3CZkEzoQ
7crFNvUEJHFI/KEZDWhkeoPssYmV5gNOPWLsVHTv9Y/T8Dg2bb4tYbx6N7vDRuD9AqGLERu4HinJ
7ARS1RkJ+CX1I7HaSpHWmzlvQAewgEXjsxAQk39oqk7FbRDkK2hdEfhEr5UsWELy5+foNgNIzDyk
Q63pAPSOmXZWb0q9oWTc4/mWLzFyv+v/BfMyZlNurbvDc38Wmx6jlokZQYL7+4GudiqDpvEKEm8F
8dy6M2yWkA/hKW7bMYzPMGJRV2ANPGUhl6ubA3380Gd3DzY6KmCD0UpxHoe6oO+JASWyY0lSX5Pz
QWfOosuBZn/8nAQsYrdU+wVREiI4sM0aBdgAxBsGtF+i2PqbnXi9C4mbdZGOCrEzKUMaKGqWVIyC
aF0PnT7QzWm0ZLwtWRsL0SeUfMTJBqN+vT6X4fVUGYRZZF85mikmgTh3LpKyv+pXbhpReqA3vFr6
5xcScnUC993O95o9Sz2d+z0V3JQ8/RLPSzKVrflJsYllJgWnAP59+ZyRhZnyqVcI1jVDpkkUM+pL
AxEhKi65bgvlpjieh/A2t/FsPfChOIEwvju8d2EkpWUO9BFgGcdM5FJKvje9D+rB2hz2DLh+L0IB
d1y/3yWBAr0RWYb4xdZ/DdyLZBHuOsna0UE+N30jgxh1lDLRlShHIAX/wkSas1hsmLEorzoTPid9
OhC7hqNvZJLWQv2tQQbpjMkDFMzQ9NwY1hI3KCUantK4m/ML05wIbyzWZQFL+KHCRn2B1l53N/yx
yxwD5Nv0JMn5WeSjT5c49V/dIsFfMYQ/99QbvXtxP9lad+Z4XdjxRY9PgUjvhc0OwxU3oU7qCICs
Vrp8UsOk7/oRF1mDFpYSAo4QhIR4mUOSuCEomRUf1NlRbIPYeBV7JLuz1nZIcScbldiTjJVjH8vS
7qs4XSQ6Avr+ZQ7BFNLEAzGhW9O8M9R7uPwVem8JoFpsu+tnSHwXAMYyjR0sNppU5xFhYyFCpNrT
2QuFlaqZxvSvXAo+S+0MJiK1WGpwrgrlwnuu5/cLomKaPJVkF+Sbo8YR+eZGfgDl/PPKWVJc5ytH
G+Kd7GPGCBfr+KHYxggK6PLBdelXPlY++QUW5gAlTlBOHq8uCpUFyyiL4my0kf3WnA3DYJNrasNT
uYkwYzAEYHdaKyP1uLyoDvpbOZSZysy0csGezB/QSbmTzq18XEqZz3X2Oru7OfjnjpTLa/ZXcfX2
7ciCTbcBi6gXivVxceSvw3jbs4Jgn6tYlrB3Tag6OskgeGev1xcAVEABeNzvHtDosxj4RPslWnV2
zVj/5Yr/ZkBc4P3VFvrr9D6Xd5ADYqTyjpV/RWdpxe4dh4XV1ny4+PdB/IYc4oRFS1Ez+DTs0huo
M99mjginMJWRNL+IPuSS/Y+ZFW8QnHbOvTPKTfRWmgJvgIvGsmbjbvPDy7l6uh0rppBqZFc+e8so
mNeUOqF13T+GKSnFvojz83snJ4vRRW5R+RrLVEr5MiTpa5uACNUWgeTTZkBYazGbJ6QBd7q5Ks3r
eWSIPvEOl4ZHCUZNk4GF4adpY0fz9zZSZK6UbgPwCTdD02Gl8Y3ANv9BOPtgrx7wJavYC4OCXx77
Heyp0A7Ba6Gov35epgFZXNBQ5Q//16XOp++VYQ7LvF+wnvYcvEFexNFpwaf2hTE9WWrFZ/Uh+9K2
x5cLBH9pzzhc2bga+hM+uvOJ2ZODGWUL8doL4PS9LZdktHCckUhuq21C8wFQ1I0ChUhmhl6YIYX2
vb0c3zICmL8cybAl7jlZnzMIMmAlETY36X8s/12IW3rSTLD1d7o3rb3Nsya9h8MPfwmaM1M3zDbZ
5IdNtKNyM1wrBSTSwesanDtpK6hYdy9+6dPSrazQH5C/sg6HKPfKmtygX/WoFZKOhK+wWkWPntd3
l/Wm+jkBGUBGf2DFPo4+shRWznGy3XmGzOjNb5BtwFrr/BWbCbWW31XlnGzoCWFh4HDaZ5MrYrsT
BNHS3lv/7INCGdbcOvOP1+ylof5Dzl/EiO291q2qPQ2JTUWwfFXcqA9zkS8hjyc0yHAQcsvrlwAt
U/pImU3vXKhsDXaGjbah/nPJGw8bDsC0c0DGqnyzinMwnWpBmhmjIRUiTYtR2tcLYSh5zocKgekU
E+XLh4MVlV5d/hub+fpJPxRMU9vmLFHLnoeIRzqukCh4D/NfGMCXwh8ehWUDyAru/Zus50fzcDzP
DIyJc8nnkmTkYfCYrJOfSs6qftqKMWVC5dYLm/iba98yo2ChkvZfV4T66zukyvcHu2TE4neC/G/Q
L2JKcuXWNxMwHNEi1DB4WO4JeobBk21N5l1g3aw6GO6dZktfdOoWikpAG5hjLd+RtgOWSU/NYi0J
HpwH6YxFyiPQ2NN4O47AWMRNSK1PjUdnLuQnKa7Ss8MCDDB1mS3i4t/wYbQrqBnOGRt+ns1g8lIn
BplSZOUddK34bCYvSnm1taUXn2kVnnS5AgQNbPd7U6/MDrDY+xVPa+/VDx2QGNn/3D+tURGfhfI1
932mTCKBRhL2OR3d3/5Xce+T4BZ8uG+bJoBiK6KxCJB+omwTFsvz53WytExJCSrK8L2d7UCvfLse
LdmsnV/hCNwdTJ1yiNM+xiDvlKLXRsWBZw8usIEFZ1IND39cSIP9IoJiWdoaPpdLQDxLvCfRCOUY
XyodVH9Q1KEdfsBqVhviX0YpquIQcEoqpn77bOpySZAy5jqe4ZpmxsEsNv0PCh9uEmE2HukS5qGN
FlonBOWNUmhYpedSVOOz2cMMTV7j0ROUTGCqo+anxguHHh3svN/A9OxubhgSUobbgSLQRdontX/x
w9TE8v1p8Jm5G43huZrrMseHIAf+nkWhW4ERm/yjktaRb7e/Ic0wblqQ5OzEEQUniVFVxIfvxwAB
qKY4Mz5ahkFBUBXD4ljVEcucz+4g6bMcv2c90O8FZB1Fh0yve2WdpBcNdiykpUKPKviM6WBpiNGu
XZenvKIYYlLngcFVSBACoGBnUCT21L1oxOGM+9dUzZOHmygIAPn0ECyrNm/otkN7VYOL05wWAEVv
Pdj00ELceBy+3Qoq/gzM/fgtj5KqD88088Qo+7UwQcI8ZNLS40+zJhPEmujdgNZpDkiQxCSh4//M
cyX+Pc9PJqdHUYQ83pljloTghUbhtE0s+5JHxEk3NooVcOpU3DO9XSQb6shru9ZrUZXWklMtxFg6
7YFL7SI542QIo5TBgYlylSFdIdMaifUTHXwSrPlAvDaa78Sw0dNFKJg4DFHsK1kq8//Xmsvg+9zL
tdJ72W+A9sQM8v7qqLN448Sh6nWsm0oHS8TWEtrAIWTfvIZWpvLBQQ6DrgXIZcgBlXD+koCl+Sh+
WjUBjQ6Mrk107b3IE57N9YO+Gqg8j45cm1BgAWz+TpUYLPKqYEqWFlxk0DW5GRjf2QrSnRZzFu9n
ts+l9fuvqaQwtTOHlNzgv7HcBHY/WXVOvKLst/rLnKo5xaMLHIiOTCF1ZjIOhn4dIQAf2TUZwKDV
MvvcAGHzllaBQRdYgF3+kdXCumhxv3Kl+WTJTSp9YGT4LM2RV88ipKNQA58Bdr6qaHbQJ9dWlAh3
VIwiVUo0iQr/4CIwE/muxOiMGup8cgg1TUJyiHC0WboPeCMGGWmH265oJO4UDrOrzYuWby+MDT3h
LD4kg3vPjt/R59jQqVKmImyCLVBpj51iWKbZYiBm5iKhPFD4grd6NGeZf+B0IpGHXdFYeMWeqQyP
KLAF1bshOTgpz2KRTzSXDu3HdugXjwWtdAylACs8zAKPRwCieR+fETjMSwIHu0iyYC8Fdd6pCbMS
ZKQ9oGkMlZKO5DSbwjec9GqDZGoqZyTLWK4ygLyocc5siUhUklZn9nfxR7aVkixwGg03YNvo/yB9
kyt8FsMgKtJYceJUz/V9JtAiCJOsD/CPSzpUYrKDkqmWbNl6KSJEjdRZjD3aml2hto4b7JDGC7nN
VA2tewZPo1NpapzOkN4t3stOS8pHOCfEiSaFIj1OaXk9NIdr6OixqQHQO8g1A7oDlF0h+UI7F8Kx
Ftkvnrl+uC8tfIzi6DNlGLJs23DdGu3WsCoWcZ1GWyuP9K+mhzt+JGMjUwb9Sa/1Kn1m2bwUrD4Y
WLqw9zQXmB+Sz0F3cXrkcwgX43Q7fWqJ46xXs1zmpqWljmvtn7TUK+kXQLs3oEkItqQWLWngalcP
9uJyL0ELeScuS+RZ+kWNF8cHWI/f3nyakr9iGFk+QfOdQgRRVyM6gtgy22sFSt9HZyDQlPol3jq9
1Z2goQCJFl13VLWfzhyHBdGPA7/DPVoWUBCG0Yl/ECKY+42KlcoPFa6wMhyCqxt20U09yhUyjnJU
sgTOXC6KWQpNSf+WyqPI/pLA4ifMrGUpQW2QLU9gcJrEBRzCUPkn6Fk5heVDWO1cymqpi/9gkeMg
KsTZ0j22Y2FzrPTcUjPSuypNbf6fiOQNw/sI/OLUzVWl/ZMcJsHmQhcwal7NL3txVrPEqwI+yHC3
BX+aefEBw+WlfGUqzNncyoZWCer5TNIH5s4Kl3tH76+op8AXBOKjsgWPbIkTnEUB6F4uk4XlvGmU
ozmahvAJjOcjo+YNL+c3ZIT8l7M5q62djQY5NnIJ0eSQ+wuwXOVl2hqhyAtEi4ku8FeCfKERJWd2
EN05swpewKe3d4JWyKJFSa+u2oDX/U9eFyJ6W6Ywt+cTkCOll278NPO8UiP5WWwrN9MhYPCsSIKP
3dpPwfsDvBeApKplvELDyLJkkoZB0cBFKcUJEZe8qPfjqav+J1OR4IH8NGZJC+L2waNl/ofZR2EC
/5Xp1nrOPBATzhRgjo2cjHQkZv7EDwz4DoN7zI1+4DAap90ye7NLfmDtkGOjGKXVAVLsT/zVjd+Y
U/F4vMHUhcxbWtaS659YEETe0Alq/Fyh+zq/HaYcrv1Jy1Mjta8lmgoWr9gP+1IliI8SOmiB784y
/Shfvq0t/NIIclNHHS+hyk8umXJ2aVWdC+c/Qt6FNAztnZEYlOllPfY/SU7xwUwqSg/8v4bCbFuk
3hSMAHr8gQTVafV1r+l97KifZTmv652w5oeL8ppEN9v+svoI77M2ta7vadZP0jDPmew4XipKEquk
Jxc2G/ah5UgpmhOrG7BpYFTIg2KFQr285rKLQbzd7s/ymoC4oFVpxHyj6lyrrYFza9fS2sPHhNTl
UDX1f/eoVaMdTzLcp8UYVgrzctfwK80cPTZ3PjgcMJgPqusaLH0QP7yH/2uwHSMTuS5TpsSkssAv
Pkv95rKcVy+eowXxNNER9YT2IyeGdxxe1NxBrPkGQAWUPVb0crSQ/EpFnZbjdCZydX6K5Sug1aC3
E4wIelb/Xg3DIsprpe5JwV85eXuznB+Zaht109PSSI2gqyrQz6p1iuqGOggJ+RGb4B4qXkH+66vn
BoEnQ+rSuBoQNWH+GhOdizJVjKx32eYsiwNvMjbMVe9VXJDOLYpz2Ziy+b5P6GCnxAVx+bUF2BQ+
GIce6P+7hnxF4bmfLbMlkipBG2OSWcp6nEbKFBuEyaQvcy96bPhheVPGzPtGM13V76q8V9nndypi
rjHoheF3O96mFDcRJ8yszwnl4W4aUjyuayA/4V/L3/MEkrdc7CHl4pPhPRCjIEZn69UDFgqsKM+X
BI6GiIwaqeT8Qa9m99Pg+eNDRV/08QXMEwtc61E3b9YvPtx3GOYU59B1ekJ/bI7ozAPR8CGoOcyW
v+BFtsKqT0n/GgYJn1LxBTxAuMp5mTB6MRUJyWHInGFQHMqHjo7EjzQzV7B9MNsykDHZ8A6GiirT
8OTCYeg66TBCzQs6UFRlmPgmsqAlpkcDUhTf18ZJ+je/9K8dj3TyRE5/7pm0KhDnLrT0Ntoi/bM7
zDO5/NiiY+utKf7D7qAPc9Wf0cKXqA6j2h4GjjEWr7+wJ83RhhwYXSwmJtIp+OZCKPrV/H7TGgSd
bCPUqfRbrx131pzxwu7PZY7F1sjLeJpRToSvueLsg07rDkvip41gsz5QIzi0TpCeNZbem/xcCNmS
sm4wjutyBMp0v/6oTEaUXV7IuYUFT2WPZKNX8htROcjfMS45xoIWyU4wH7TNnXsDqbcx0iNK//A4
paK6ppjFSZty6ixycd/X6gebyBxvjxuV8uRKVw4k6Lf5W5jYFB6VSEiOXrfJhxxlBf8wI2KJT4br
RduptE7m4KuG9cKjM+LabxvhlZmL6vXO+K8sxyo3ITxlfQwFmsCgoE6IZ0I0KWbvhP8WBLuiBHVv
kJqqOcw4utPbb/zINRHeUzZPkWUYijB+x9JbjNuRxCBm1R8q0N2GcqMdweaT3x+Wbn5BvQZBSZxz
4Z0NV8zgYOSpsa4Q8PaLjW1vBdQJtdgLgsqHmcv0/rcY/nnvg42G3P48A7bc7EvydLv5n+7AEnqu
/YC51F4hWA0/rZnN5MtWepHqIpOs0NQESNfRzjzTK93nShk/siETr4aA2qb4TJ+mWRYUyWe2k4BT
hSxLk+cFdjB6pMEcHu1KJ0gsBhRJZkGizIc3vzlUXSlvzyk75RMQyqqWm8vm9sst+Rrn7aJrKzi+
C94MZla3ASE57cg8UTLT9y/Fy3LVQp4J5JVFymoqzQXfqINp5hQJbpeYwN3xNJmqX2MrQPmoJAPU
wMKvMf2g4IQg0jupM0OV4z9cacvJ0whXmFUqL+HxOfJUukGMAI5GqM69pycgGeobSfuSix8H1uO6
e3yHoO+UsVA6VmQDbr6n9zmgcFwTepeYmaDlNz9MyAH1F45C3UduOTNNmepsgk0SpExEZsc8UhUt
eVZF0mduNsdGa0nv9izY8fIn4Q+SkJRErcF7T3Ub73rhN0z1/qjuR22HZOVBzXuLdo2hgSH6Zwy+
gV5z+eK0xU8K3mubJOgATVgZ+1aoDv5eKR09M85J2CFxXvo+M7+R2pNCs3GK1a7i2roGWxIAMWtd
QjoHeEqBjwtIl2ys/dlD+5y2KsLv74tjQf7ZngmEzsYaQ2QH/MYIFEEjhRV+XZHTktgRPwo9Uvbd
7AD+kagCa8RjKZiGhHh/8retz7UIQN0Lt4P3kNQQRbsvHprOV7l28k/8Q1K96iNOVQa5jhAaZIx1
QlWPpeNk8sAtQtwSMpRjwDk6JAhI8XZk74EJ3qqyx+Aa8HiqBN3XZTdFc15p4QYHqxoL/gtGEBz/
hNsNujfOTEfeDJP6YuqOXstHoVRJAdG5O6x/GaCo0EvrP6Kv43hjwOxWYEb1xV9bCFR9vC7+893S
lQxtWA6GWFvtJbTXABcRQNCMquljhQgiERpzF1Z19xiiryxx2vnsAsAtLjzoDZPUUc1HsrvNUUyH
G+mDR4c1lTR2NxhUscY6tuBQ7jVUseZdWSOzeToof2DSWY0o4PtFl1diHk9i5wvTCPP9HC19pPkD
QvRqKcqct4wDqEoKVeAaKgWSpp2V7eQJD65JH2+WsJv4vRPkn1yGdIBVuLeyymBu59HlmNsMdRgT
yEY7IF38KQbho1dYo3ZI8wapLdmfviywyTV2JHXFLL4ThMV7WUu4yWj9nLJmGpGcTC5RpjKbgYwO
mPUne49NUviH/Ud0OA5w/ok4An5E0yucdowAmx0mkt5J1458Dko8U2LVQHseKXkSgfBZl4jq6ffD
jznTtYHzWFn6fYjEAQzIvRSw7k/rzM/feneHSGLn9E93qXxnsxA/nznpOa4i0YXznK48H6qwd4Ev
ig4Poc6mD2za4uRs6mqLk6CgLz6qsYupcCyv8vuUQI8CxTF/WsGbv1pMLCiWslIs+SbUCxxcJ3Cl
Un/vJXn/9vHJAv8Kha3q5qLrpM7qyfGK4ryD70mc1uBY3Y607ePzOaUxCHxnE0nr7u+QBeVBqqrv
DOJcYt2MkC3mrTy6FOPyKQsGrnwkj9YkkzBL/ksM77bS4cikkiyNAMtFfEZBPP+iBoDiEoHljsY2
wfnds/9yqw2HxdUm7z0QIXvM9GXqzGZc9u9O6mqHdR8n8N6XohB0GFKYrXM0YatvJ8yUT5QDAKtD
tctE9U/eBo+XDnIKpjQrcqXS5bIV1qju1tJJFoFmob+WNQ6Vax0SGHXnnBDzY22Q0vXJs4q7Ojfv
ahUnxBKH4zaK8u5dCUBQk7EvsYDZ8B02S5AycFRIPEn14ysZOPbvIkQWxgafbxTBHjq2gXSVQJ42
K2JIo9ARi37pI94+uG1tWfxYbg9kzPR8+Dl++EmXYv/h3QHI43Ga4tafDN/RxkKuLwf6NjpC0cYx
3lUoZW49o/U0OMy1O97frrHx0mFV/HbkJPEkOMDMr3AVmJ3hPCEyMdfd/xNCGqRyD19RnQW20bx3
zQlGAYdXebv6xDdPDznXKOpJypS88rstENUS7xKgp7XX9GJAFX0AYgfDpHV3Fovn3/9E64ZZPz1J
zeKdPXwdRCJdAnZtK10f32bzUdO+vGuk3Lvah/H7rTMnOAuB1futKthz5TSY408tv2k2ExKC1RqK
nhaSIxw89dYM28eA2h/8zEaAP0mGHeetPE1mxFspDLwJu6ts81LpGoLA9NU8gGqOX7RB8UPGbsFo
Ijjqc63G7RHAPAUebOO/R5JVDTx1UpHupZpX5yDE6+abKgQIr6MoB23VgXUg9GVgIjgZl9Ap/9dM
SytHUZwu6epfC9v9zU95u9NVopJnzcKKL9zX5YyXwHg+s/DlC4ctYRHOMlO1jv+1UBc80aSrUMeC
BQeWJyi136L47GZHCRuEiLO6dPaS/cli2CbB41j5ZjnPEYRRb/m5XvCsLl6OlHxbSVn3q+bHsF3T
u90B1e/s2yGgU3buJyT28a5c9F7tMMMLlgcQXlpeyNWMGtS5TYKH291ZsxmOdnYKPZ8fkmpopnfh
58zs2jpQSXlnurl/Vph09aSmSzXhHqQUqT2emeHPRwQrckhD0KeRSRwT+zqj57Bwh38fAxzAm4y5
bccNvgDqKNWhHuXCdHBx4PtwbJQmKm337v8nzG+xJTVJDY3RmrzEcB6Z5Fq8EI2NKd23rMacQwMi
CyeFr1TS8PGnkI/wLiMVnzDyINz/+0MJ+GS4yMFkbB2Xb8HYT4Htk/wJRitHkffRzJQVuEku4AJi
rw9EGyhMeAtWOI8xAU/bJERrP7da3Ai0Uocl4BEZ+fcuehH2yauQQPhegL9m441xLkBDWOgSuM98
tR7e/xNu04l4nfyaUQogRrwAsQ8NijB1/kd9zHS+JA5KX3zUb62GrAlcuW+Zt0F6HKZWZXlZmRTQ
m16jorknSVg9fGDmTixPAfBiYKsfnLwVuB9DyPWTA7SaUmT9tBHgG/GCJQL3MIDiHjfpJP3Tdx8G
qXMAB+qSuwJqVeLMog/hI4uvCH/27PGVbe/OyTNl29PVlIMbpbSIOBIsnLEeZzbIZl5rGz+V0eu9
NJ9NCNLElLq2o6t+/MwTIyptWBUH49hWlBPkhcDKCi49JzUWyjGcUhBDhTSQZms6ZGJ1rmcF+2a7
zvGcFYaHacuisA4ZKIM+FQTR/QombBcK7xCN6rc2Yt3ERdc/sEoQPb+MM35nxZZHNnuIpQEIJ8tH
XTq3uRTI7SQI6u036KKYL+lzge2X6emBNowa99jOQfNtVPSulwZVCKuQbSsmXUIncpDy+lo0JB3a
GkZcC7kkphAlY2YClipaDkU8BYmMnB7Y0G+pSa4ZwFr3prkGK2s35kvJBrURdS1AD1X8bh2JHVH1
uzFupYPvH2I3ErhGC0DvfbLmZi/JbipyWOX8yGFprMZ3vni2MC99Q49bVmOz6yDxiccmUZJPQaQ0
UYW2ROUN0tHGt1pyf3LKwhJ235CX8+Td0TVoG95iOX5BYfwDOcIarHefOerF+puxnSL3S5ExZfRe
HXZPThw/G16ck8TjGI0rrm4rDrhBnaLjVzKfDq7bBWXj0k3JL95yd2TLrE+aTLHkIYWvD0Xq+rYz
ItKugSGWL6aAlsMW6RaCC2V9pWNWssTD9Gx9eysvrH9wbf0EUA0uV6f1HaEXTjgdoaeAWt5zd7L0
eDFuwY9wwhQwZIvkNgZvgBI1azCsmfMq02iDa0NH4dEjNiABh1pf9VElECpFd1iSv1Z+ZyKczsAI
eGiJbIvbv3fJmDTBrDvqxOxibBETVHEcWTA/OhWxwEUFEVsKPPyLFhF72JeJXh+q4hBjE/MhDsQA
G6K8wlzr8O1LaiUUKnuNWcnKKsx12wmmK5dSc+HkiqfmVKtjvTmVwd716bkxQmWrxUQF3wCxTeVb
+LoafgcVKiIu0a/O7vhHSzJMYjWKW0Enu+5LPl2K5HRCbxV1czD+SpW6MpEbhYG2WOKJ5pVehfaZ
tTA1/1RC5b3R5/XSfAw21TW6i/bHeexMv29g6J/zXFckVsMAGttil7SuLcbfL8HRIES7xBliYF0M
9xsPAfkYG/HeE0w5x/XGX+FmcadlK7kzN4y61qzo7B+xGDqOELWsOPt1BX7cQpmKtLtxV4qOCUen
Nx42vmpR5sIbNULtWWQyPlkFO11wkRkckyiuYLV8UpkeK9EeWpYw6qsqMYXYjHsbsh5RQYT7NiXf
ok+d287KEDlGgMxsq9agHDfZcmCukLS0QesIZMI03TVZiAhPOB3eAW19rDeYhK4gX/h5V/b1HH+T
WxyTlCdJpN9/Mh1MGytegmYG+yEPDnR0h9ClWjiciMgsm6rHAtROeYdbxSDfusxSMfq8JiGSyF9U
tqgcdWhMl+JroncQWscOdln6eowi/ZNdTNfg3zyCoh9/U6R9mDDJAdSDBhK6gwpEgRfldBwN71tQ
6kX70KWs6pxfhbfBYA3Snn/gaoDYAhrynb5VxTjmp7wN+SH/L6rsUhRy/tewgMbl3UUMC+BI1k3p
HKqcYPGteD8nE5/T1RCIfy6UKFPn+R2bqzxGW4kSGU76c5uaKTwvjMdGuoJ2lr+uxDAf79DpAqWJ
OXg8DfOG6bFHhBrNyw65WcIDtPPo61kcSYi4xP6AtYapRj6S3B7x1xL01d4NVy+UXOQH3svS5j9D
8sfzMz3l7sd3pznjon1mHafzpsQCp9xDQlxKeS7O8CiNdnKt9ipE7ft4NSZJeniGgFvcYJ+9Ztqf
64eULLJtV8sf2ILIBkRxAptNkntpF0iBL96+LVSN06om2WvX6YyIp2CrnnpIw2tARTHc6EjQ5wKP
cb+ov7ngw/8/z+IOfIvnGn/5Qpd/AnjCaHZ0MqrQUSlNbHpCz15NZviZhQQiv2S79X3mCD2c5BDI
ze03uYrlYYF8iBc66HqbDJ9OEdJJbw5mrrXK2cCLfLBfA9T8uBS/TsBgPLkD/2f2nAt3MECI1u3o
oGlYFArHTLkO2cEmyi26W2bPBwJIUlTQXwTji7qikrDCOPR4KPnYcGuHpDt8Ht05IQGMJUvLPTNZ
cYWzGPbQO670zoRMxyHXxqZvYZ2eqfN+Z4vJzk3BI1yI2n1FvGf2Ju9kTUm2cYBJrenq3uWSaiMr
qGGLqLB+2mGNNZmBUpvz4qoPQCCEW9nhU7amhWEP7DunkHR6oQuZOfRJdnYLqaaCH1KZKlyqh6yC
cg1HT/iBixZaTF7WLXFSi68v8aWzWwy9iFDQWd5lUR0Km78/6yencJ9k99REzPKzjwLjbROLLLDM
s8pH/UYiIG5fs6XesFDF5hkuFZ+AVzkEEhTPo0y32s45oPV2XDk5W6Cj0j9lz9IuniDBuGscILGb
p236FNXRMaiq1IV1vRbqFv1VmIXEqdNqMsN++2ugj8Ts/RlipOqZMP+XtC+KbkcO52vbrFZXSEPA
uNna+0HCIVZawWPBH4G94Z8CVD0aISDQS2ZnRO6c0XMIMeLe7TvetUJzUPzCPv6RJMx/SfpMMQzr
ThJeU8xzJQRtxC/pmJEgb4bNOGpdgI2wPeK0Q0vzm5CXXSQFEOCwbD1LDp0Oeo6IK9G/Y5BFxQ8F
N7sBtF47XLYZl1zytB1W/3qiwFDmi75nx0KWEJLVsTZrJEM2S2Yld2qbHRSXu4hiD3YtaJdPNzOw
5l7Yf3pqtiQ77GJjQb3Vy0Y8nVxHx6ARWOpX4kNVLE5kUmivBiSod3VSG8SLmg8GySEgPYWdZwq1
3mFPX7061dziYI/2/52dJ2uDPTZ5EnCG3IqKvFRoGrAqa82id8jneEV2vt7uRbQpsD2uR2blw9tR
bsqsWN9Is+ipFv8BMM+BWgXYGtOZQ9EtOK10UQiP2TvTz8z+TUi3g9ummNuKgLpKV4tEduf/WymM
xlGLICCqtiQO+TTqJ/7tc+dBc0DbYo5J5DBjz6ZMuo3wxRbkLGlEX+rpDbtbA5tNmM8QNs8OM74V
FUn2Fa7wayR9gDF3v+Lx9KOu5qRulqELkUnfil9k4DKLvgCdvB9dYb6Rym8g5Nqkv/7lohmiCudP
fukp0aofKmDHwdP2XpAPAf2kZNb2aIjsKG6Vs5ryHMKSPn6+dh/DIyYlVwwpV7OTAQfrNvMAQUo/
vQy5brMp+rM3NQ/ZhRP4ciLZ1k+Hvv1Lugk4BHb2f/o4qrM3DxdIllP88/MjRUXmWp3K6Bt7XIC5
vqlljy42eJvd2jRFnmfjiDdTB7TSmahOwdWsdDfBMVcp8hcaMvoqInKZ7PzBy58rcb8Nb8KIdnaa
p6ytHznIAe5AjkERLxhMbOMBagx/A2vWlsmsjsrIFpLCjTa7/ptFeFFQ0OTmPYBHiBdlG1u00Vu/
3/ltz7PY+V/MfO9IXBa/V03ZnTiABbOIqMsP20gZXXKNY+2qkUSdYbRb4fuqVJwC5M5iPUHM4+yb
bzPHu7ogs8v3k4AM9rFWeldLWocsAqkmoDL4wdOBar6FoIUsXgvMWlNaTIHVHf7WA+yyg74xUdqx
a7IVJeYrtcYInyvf7S9wmoOBE9+LEKSjyYYKQ8sfZB94vF+NOl8PqQ1MLUkVOpS+h7WeWDusIpzB
JTKROXYcaPDWXbM2tqoHjaXsDOx7QXVsFH/maT8qA6RNszBwEdWOhJCX8tvBr5ZzFL+bv5K76epz
+iimC6tNm0yqrfafmSGluJHvf9ZnMp50bXt5pctxUbl9YNWVU9V3nWA4HvwgcZn/LOFuAd865X4n
Cw5hBzjLWev+pF2Q/INef2520xS717KuTR+D/RjdQUsKZlNwohDb16NerMEhgTLehCWfcGlZINTs
jrRe7nytgR0Tpibq2lLim8DaIk9tKSPxLTR5LYIxRDbaimb5mPB5MFMh5zvpWcq+JaMkP529j6AC
deHE02jBgN5XRztmfTVdDfiPZbgW+CeLNX0B4KFVnlpGhdT2fLXyB0NDCUY/snYA8iiTSn+EABxU
m0XA+JiuQaBVln44rWHaEe+sSjcKzJQ0/av2yeP3MAiZ8ff66DRcn8DmHUC0lIbFSESwRoXCy9Hq
vhuEvzYaGqCCATFM0/Abwfrnnna49yzUVX2EeX9S71j0Bo89pC3HLcoJreD/X445SslZvJvtfN3m
IH2hCwoPnB3ZBUWGgeK1cusjae4Li9LzwQpVoZJ7gQ84/e0aAHlmDLKjTkdQ3SaCiqu8b8GECQGq
DRL5ALXDoT0Wb8q/qu+HsVf4deB2+XzVy1L1/zsh/gyVbQwsgXYeeTUSaoLQtIkRLKWBzXcHVMD6
z39ZytJon4jPRVwbdDx4jFfZ9imd8P7MC9I2UaQmXmtEp5dLtzrqUBOlO7fm6x+qcIhZj+zIoWlS
CvE5rekl33DN1aqdt0SmTPMMMudFjkIwzRcI/bg0Hyggo3tM4gfznA5qTjA0i5hpSMTgUK+HMHlj
W4Hw58X8jLEAj63JrPonA/uAGlpg2XfcLZHuiu5Bt11hLXvw3YdcGMAVTHeUpXQjFB5xbCq5X6Fb
cNTArbIAdWFnocyKI8kR3KIgFsEDKt259I3wP3TaLZyQq3kT5QgrI5xaxVxuUf72nDMsjPtyAa7j
BE0/ZUl2IBLs9DHVQ+XQ0eSxzGSfjSz8XRHMbX12Zfv/2HhRsZIygb6622zldth4DCm20uQby3qX
q1SYPCq9IfTNqB7Sca1LL9Z9OSk3O+2yLzqEQC1d8oTK/ml5aKMUfnye35me/2ivnslUKFy51hQ2
3jzMMac8KvfgxXesQD17BZjyZtGfYPubSq20/V82UKlNnMZAY52+ukD8FiGbHWc8y4y/5BJcSNML
K8bXXK/YLsEgOHeGk6/a6KE5fSsTxC37ieBNdZDveOpZTI86IyJod6zrVHNiQeQy2h9afnJd5T3C
ehZRKe77LFUBYPpcG6jZHnmdNheDdSkNyqV2rpMthyY+yi4CUUgB2zBB+3fEHYulcwwiMN7794tA
o7DqF4ptS33kZK2NRAjYjK99EzrR89TwnRxtPpJggFHgsc2fapLzR0bOYFk15caM2PUGmLwn/T3/
AWnWBF9Z9TdkH4MHbX2QhB9toU4TrZGjms6whuhINohLgIpPbnT03GmgwJYhBaspxEiO/mqJm4oC
Opu5h1PCkQg4pj9GvHTGtyexVUFpmixWBTeIoMp63Ge8YI31jjOGj4jFTH/C+cvcRJQxwAOhu4Vz
lPPMTG+AynjFe7X56pZw7l4CYKWf0ZDt7jJwqHbWsPmRGppuGHv/QjXeiMnazO11DZXgCY4DoUGV
vPHjh056/JLTFfOKhHMOwwR+pVaNQCdJbpi+ytHInMFPFSElirIii4FR9/Saw8jmCl44q+r0mlEP
JSZnXuaL6X4Y1uieovAeHDIFZ1GzdK2jM71VxkqC3OMo3CVqvVbXUuxMEjNFBSYkaDqqR1kzDnDS
41OH98N6+Q83GyHiPiEo0kbxPpHIFj08E89CqnA7fw8+8H8c8qx6eoCJUGEjdviAlzSU+JiUIDLx
XcRhsHlxnz82HCb6d9wXVwVaqieLM34YOA+W1K4jFF1h45ggsABebHJA3XrXSJ7qmArVajDNYDOm
aiWAnTCIy6JU5c3zRyv35Bq66zRXqfKPc/duTa7/t2zurtwBSNVy7zfJ7dDoT1cdut3AQsQIe+im
GcW0VgzdAtDoiJYFC+2JpgKj15aO8AsQlKFGhkcLNKdj92NXVa3N9Up+QJZAev7jmJfow/kmH4Fy
f1TlSKb9PZiNztNazZiuw7PWbbUs7UyhJEOZkaYVdZ7B/9RX7TjxUi/8fMVXF5dAJsjIQsVZ6m5f
qOWbvjH+BAHyZWEMMGlXpzU0cqZaJL5fpLqXF3aW4o4iuV2K+TjomCK7XNR5fcAypBEAmFnfJDf5
Rl5kdwPoJiNHVwPgvaHQIF3LJn2yIfGQ3GJBKKXzSfgtsgMv7D5Yef9+9Lh8jaMpTCUc+R4u1Lf+
bkzqAn1VE3wkiKJ07azT1uituamQZcuYdV0glPgdtlFYIajJvEwKnpfzaoZJsYYwYvNfNeyqbp5V
Gp45yuwPIWJCtx4s3HTYt/umNOu9qvI6F3QLlw/oZ0KMenAdkNKuvaYqDFBJRD6AFUJFp2fv33pL
T3huTk6kylyTmofnxJvjELRjCzXb/9idg5uCsXw6Quq/425VqQDIQwOKZgVNkLyxh6hDlMnmXtbt
LwpSZ9ayT0Mve8PQ8u64V8OiSR8u3VSkfxBI6e+xAG6wLT15uWfG3Q+E768s4z8vO9QnMKTQKHQK
vGQIEJhwkLZj4CXro9mazK004aX8SObdo5Q5UT7iitOoc2xcCYjTN6Qj6g+kPbf/9zBAZkwq9OCx
CJiU7Oksmga/ljXbHuBiGpQ1RTwaCfx0vTQ/lwHHTD/aUPM3Ua7OZQGIKfc0dGiXzynqWSr4sH/u
Rr1ORH9qOR51EUsGUQyZ8x6agBAEWGksvC9KLxCT62oKsie5kxY2Gh8phYffKWWqs073Z5gzKPYm
YuLXi0WYSWwBD9ZGCvISvvcb0EjaTkzbioYPbErKH3Qn3OZRJY8QakG0oF08IX/GQNdDRKjO1rhW
N/vGuNKs18TEHDBelQegV/SoP/ftefk2iHYyII/Q+Wa2EcYKvPmSKXnslMPC/V/Z1TmkZeuPz+sl
tT5RbRQo0jyZ9RKdBQhNRZKITrGyCYqBrauI0wK5Se3oqBsdZo3muzPXpIIDxjAbRsMNGgjdhdIe
wmnVNNb9ZL6LX36K5Lb/q5+fFyqRdomorsKycaEUHPcJMdDxnfszibfi9yzpWwHxA89GjtH8hgDy
pQVgyFf9+MjQbktiFJCbkCkBfbe13XfP1R+MGLh3eOgITQdL4VP5qpgT7w3r8Lvqah+oyi4JBbjS
y/rzJzpb6F+cMAf4CTm/pSVhYzvTFvSwZMZnCw+mbnG68FM8lAJQ0pSFyhD4Ky+BZ27C3nOkm/sN
TrTxFqz7sv7v1jzKYOj6yk5cP7D7X94bpioaofnntqe506YQ5A7jBf5tp5LDmTqQS6azQn3nA9w7
2AOO1FHgUJTvP4Xb50zTpP/tVEZkYmGuUIkANEtWyIaDjUOkOU7fBzJUYoidd4V2TUFuYPiBjJFn
OVQlfy0IoR6pxX0Ah8M7YCraLxPoP62OPRjKxD8dscz2DIJhSaSpGdwWBfwFb58n6zQ2D+CiBTOE
zYMxtxk87VbYMtRtvyW3lJ3EiFade39dD3iRNPyLjw79MSkR3Ajaz6p15KmgFepZWuegHlfebsIp
zniDCmmAoOaZHLJdNUSDynMCfz5kLuKWk82pJK1oob/1/j+MeYGtqC0ScW6swu0VnVNC6mJ4nhdm
JG7AzVBKWsOUs90zei7YLOVDvaDxCNrzB5GonJAkc9KoCZ5WOm3MesFP985gp2ogvls075N2NsMK
+wuCKPqVh1s90K1Vai9xzd8hHiANiMXHqO9tKw==
`protect end_protected
