`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GG1VZpLieZht8VL79iE5Jm/UmSXf9KuxUah1MkxT1HMot8/Hz66cEGOOx8pGU/3bmpzDQjlWuAKF
wKacAmh0wA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e8aj10Z/Qr6aEWhOutFhtfBmGt8kzLtFD5y/4YqbQWY8D+zD+JO89I0mDMr69bykHcl3rulon78z
aCjJzFyzI5NSGqgqaJtvKvO3xqtETaihGpGY+1DHVViok/V9uWuSuCUmk0qzQZd0I6yTLAOJ0szY
Xo6eso8MG0q47MT9ASA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nxVIHzRqMnwWtoU7bk2TS9BMEABZ5Y3qiV9C5qokFKvn8QmRnszHXOxNKn1mIPZmabW/MxhPIMoN
V3mL6hwYdacDV9+ZJv8zXRW7q3eJHEPgelvClVCaSgSkLfWzZI4+J/BqRfKljtSa+7ogSFcKzfLH
M9bkn6YSNqLTJKC8ewoY1QYjAH+wIGuMjWqRjvLCsKwswimKTwXlowseR7NiStoLZbOfQ3QvZcmZ
+sypm2HiwsDdYB4tzYZeNnatAmy+ST3bbJH2GzMeFKEiUbN2tmUBzjOxQQCcknBYtZ78izEdeIc5
yYVlV4FAa7yt+ZUaPkwwkSblVO4NW4Fl007IlQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
piuJCaSpkwpor+sHjjlNdxoKJctAQywR0aQOLip/4h7SSoHWemyg8YD414QPr9TwulXnkuiq8TYK
OSzlYsqTwXGZFOJVUg24KShFyIjbKGSpiYdjwDJanNkeyxER1Iqh3+IMvE2aC2J6mk0wbrlsrA5Q
JISy3WmDxxB2frvqR4yQUM5mq7LBOCOgiRR5/gQTkl1aD3cbUsfuxUYVnslEsPVVCBqyYwzJKQmi
1fxZjbyv8nlEOtnFS901ybow/gsfHFGGq9S+yS5aaWnmdz486RfxEBlULnj5F9h/Vji6GVqLxOvp
r6DvFLstei0Qs3Atk+HJZfiS5sAtfb8XCJ9Dqw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QvkWJTPB0IrTVJAfKpulQlyJFHjxGZu3qHwO9L3qF+kdTVs9wR0eKtZ4Zy0Kj0Ek/Lj0Df2Cn1wk
OL7liiL2WnLM/NYoh/sNkYbATYmnG4Zig3B7gXv8xoNe8GGjN/2hUDCrLsoAXU6UPXtXoH4a67oE
HkrHPERSAitMTMbuvYBUENrJaF6yzLDUvJPt1jo/QgbBE/IdvEgX4dGgddO2uERpXGRqzPnXBx8j
pdS4eJliVAtztSoaxInXYxvMaMfTJnl+DWkopIX67HgweHH9sNfqCLHemvDqO4NteeQ5HXF6l4G+
2ThgcmkfBiskutO/koT583nZfO6SUDK+eEG+0g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q1h5f91FzREswT6Dif0jspBp/rntaZX90s50dY8bIQapHuSA82tO0ZRvmHokEgDKfBGvOYRe60DF
2l1CRSq/W8Wub65YZyeqKMRUodGd0CkTQnmUC3C4yqIc7RA8gWzBxO7JBowC4gSxCxGchC5gDL93
ZjcOVMoBmZ8cnRx9VmU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MwPaGRne66TjIy8zIiMryKoIeYPjNLzijwDATq2+bieKAZItFKPycG4aYVvIJmcrpdPn2eLSwwNL
lJT8LKv8z0+5H6pngIMq366V2hqMM2I6H+wjIgZnGeRfiPiPUF8TttfaxriDkfdh3GngTgOJu+bc
0x3Qob/BQZOKgrAzqIGHYRXO2uoq1FCmjNrXXgXEmXUOrvf4xS9dc5IZznRGCRTxBy4qQh6WRlS4
BUzI6hE5x4RBbhIQ/2h2wyhuNnfR1OuOKowaXxVX8EcuM0DptXKJPlnZeWKfXtmjMuMhlM2NeiVS
k5A0eEgzSUBiLHZfufeMRmJELxkOPNNrWNaekA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133280)
`protect data_block
fbmHNJSxzBRphQKMV7XF70fL69iM7wUcBteQtajMntBm1b+BlKxuNLZDWCl+PqpV4Bdc5v1yFkwj
4RN66ASLjhTmBni2sru2RaBO/clKtYXxXcMQWPbGE/PMN8s+u6z2F/kAWeeeyTkFXCttMgwNbAw1
+fAzrivvFwf6gyndKg/Z6OCHoWk3h0NgRF5HlH0vxmaXmEz+5qi99jELyaF7ITtLGMV37EkLaiR2
Q9yvdNm3Hc6GqdUYxXWYpgyydIdai7EdVKVyXp/1FFlmZF/1Sux2buYkrfo1a0ZvrwZPH4EXzCYF
XSxMruogihaKtjl6zKpHsqldFG1uZNxuNnqLudgQsuob4fkWOTYDWqXtu0tciK9vETG9/k2x4MUN
GhpK4xVjml+U4y+Q2d/e2612cXQ0YW5KmsIKPkdXzFUp70m6RI2Nky+OyGY2rTydPLY2TvUjwPtg
0rXbIQNUKLbCsQyqW/B36UZBtkGw16GMDYEYDSAam6XDbpYIQt4xR9J07bTCOR2r/+wb2UfmCtkF
eQBkEvdnfNapezFWXbKy4dvCd2fcNtm74it+IMPubKhfkXIgD6lYA9AJIdjiZP6QQtC547Pl+G4u
7kDRDujrhp5OZUuIA/2uRGDuzSVsM2oxGRBttmqSbSCw2LMgqs/LAot337Oph/FOQpEEEYyBdwEr
0MkWWkoUqKMC0JibZrZjvUtCGkOaLkt9ZL2A1HtHI4rd6CMXeItX5uNiAl4PKaDsTQCiW9N2UJz0
6qZzaUfmYtqw0iutKZur3I8u/1m3LTF3ej3yipe4weXpZuaseqKgbWlAEWqpJ81WpksAefN+saWf
EhwYNo19v4MKyPczprBdsXvDbnGcO0u1M0coJXPZtTqzLfyAqkyzgmQ2kZV3oOpTkpMFVlAzsLYq
teHDRHcqEbWHD85Ai5MBeUluiKY3fMFyKoSnbkpoCQnc5lPXz3JVYJtmF7vWkDFy5o8DMN67smUq
hTpt5pHDCJgmRuJk8LNePi4wHNE8cTPLiEpc4tYrzYl0TYhRBE7OQDNm6YdG40XL4HZz3YBfpnDL
7sLTo1JoD4RhmsIa//ZHyo1dgoGes1fZ6KhQk8sHiYr1wtxZkziO8LZ4MU6alW+0JoBT4JFDyWyX
kqDMhHTO8S7WYo6czZp6NIglqnXPBp9nnVAQzbM0WiTWDY9dfJ1pgqhymYns0/SX2CFYI/NsTAXp
QsuaFHRhf7IO417EW6ABqNNWiS+QWuw24ZIgSHeWho7c1m2Rtm+CWJSs9uVVT3DbaYjZQhDNlCHG
brSiRgjZHctiYnxCpRAsnvl/cFsSJLGRBwwNJfvxlJ6tEAj9CEOFpkgPtPzUww9EkvKRyFQEH7gV
HtnvMDwi88GZkxyUl7qVSx/n5hIn8+mxtDHcXB9x9fbBoOWvkWXFcR8Fj42MR5ZJi92kemFdtal0
sRbEFOUmjEcBy3ecrbfZSVZGNTgEzI4r9NaQfNr+L7BUds2tAd57ohS9O+vU1kdXEk7BgwxQEPnh
WirveEVd5d4HNHUp32VhAGu8+pPRZDoRYeU7K8RHsjmCcSqd4mu3lDQZVo/QPZks+i5TVt4bg3JM
KRPoVPycqkcvZKPAGxNhj0D9EQ81tf4/KIok2gbLlg6ClNwdnRjx2caARk+Ypvr+lyJy3xmzCI+u
gNmci0EWIchVNOvzcOvvQdEvLnbAqS8e0t9YIpqjceAGLZ6dF49RotbREHEMGySMcRCAGZ6furnb
SViwdr2Ib63h9WxTMedWQ3/DJszRfxyojmJsjjSdN1p7T1gSiTVFwNAZkJPZ1CZObhBE7MN6A059
3c+ui2GAjLq1LflGkw7nT4OAPcwl1jCI7JtNHG9ELabz8z/V8jYzDaeVUhY5cECKxQMgZ4Os5qf0
ylJ24pGuM238oi+ThOEqhCsH3L+2zZZb2h235yIjAWS+HaQ6qNOG17QHeYZogc2BUQ6egIuFPF5h
ej1lL87WZ/URwhlH0SWh/f4y6s2w/f301aOyWVEc99DBcP23oRvZwq/OgdNVB5yrvsaySMulqVsz
otYAMpPwwE6RRYZcTlXw2gLFxX3Z2554+Qyxkm3LgxGo8/EJm6Ra3niwo37qKrC3UCvW3fCZfOsL
rNr2N1STzuSXIqQcrrMsxdIEsenzsre4bmMWcK0PJXUvMHhbJW1gPcRWii6iBx5/FqIRl5uzegc9
xbCZIjc14BhdnnZWifSZytBVeflw+mkuv+NNL4IQLhQkojO6/JhF/kfMWr7UcoE3sqMspUJjUggF
uplCo6FJvAEkNnz6qZwS4qqgCgYHVXIk3M7dhAmT1dqT/EGoYZaL9mMPeRpqmkE06pQLLqKUv2s6
EuNEbkq2rtm87mJsKb0jWkUHYfhGA1qNErqmBLZLxOaeIn/L8Xmf57YJJv5q0r79VbmcD53t5owi
1dRTssmRjDBgewLyrTTpPbVdQSfnwv8FO2o2MmlE8go9RDGfIGa1gBT0mSYARUzlzqKiRk6n6ne4
JpSOyYrHI2EfWI13YwXDcQ86gVkiirrmVx9sYRA8cYkcdl+p+scLSbVTZgkknCsP2YKsy8POCVhO
R+4xEoNhg/eoB3HAhoyi0dov4y1lFzDR6/QTCEsBXtLEZ5ZGLM0bWIsRbqN15xh+MWUPPmdBQU7s
uKNkLlqKUzhGOw499/yl4miAdrr+Cv4OvIfwrzauTvBuNwLpscriHH5ttCbQUEpi1GYcUFfcj0BP
2ekfZzBlhW8gHUaBFtCf+Ar4zylw0TO1t5dL8cDEOv7dU4igO7kgIXa4sulzZF600ynv+jUvoSCf
lOwA0DSgHdGSHPDEdn7DewBATCaz9mDqkgrk8HP7mwgQqZyUj+vuC7AGQGb+GfYU1HJzw1aPyOaH
sSo0Nb5vlglSgWdblI4oh8eZN+XH5RSTOp0TLE0Z8GXabYVsoPK+YO66jXtZLBQMwMw7bec08Min
KmHXRqud6RF3qf0X/ISoIluIBg8x18dkzePbs0Ot4rAvg94dz7NXEDijW4Evp3vdFezM00P4iSJY
2eKNOMdeGA1YKoEvdenQXtVHdUctS5xOtKIWj34idgYldRvitNWAjqZZCfCwUIq0CHRISxibLBlj
0SGn5HEn1QLK2548Ko9boMd6zTAxj92mK/ufE8b8NohspMZb0HAqmHjSMhxWeHKq3R4neQy+fu5j
4XNNR+KnnslrSn2B8pf01PG6USQZPjOFchHbre8uZH+K81DKAKXYoDBUPao1Buwn5Ykm64Dj6jh5
9mPDC10ANpBqyCXEflm0x/lUC0syx8WKql04bUg7ekgE2XaM6NOoEzDErwKZvaDTHyMR4D3yq2mX
/FfoKBTbXEfNwt9NEh8jerpToMmyygfSGVSeYZjXia8ka5yz5K182Lp57rmwqecMIF/oFqms6lwF
+9dEqXs9v/VBGOm7u8LJMbnsNtUDNwvREK1/MXYAE5WzkEqb9nK8xT7632dOCLAOBDNvPp93qL9c
PerkghjymJpJG7Y8PdbPyUDWeWnzHnx9khc5yKb2fZuNxcSWeERF7uhc7mEFO0U3+eLXACedgT2c
xZ+FtLWn9T6HOYZxTqDyWG3YW3/BzhiXkzC6Rer0VJ3YBBICeNw8TxNsYZMEF0ZRvbzfKk21kfx1
juAmEetbTCG9J/V71K75d4W8P0jR1WF+yd0+MUBe8fZ+9mr8PWcgb9os9BFIMNavcuQodfPjpshG
qb5CvHb5UNiYWAY+IkWcY+7nQ+MijRlZtQn/wyjDFWq6UrfgRKK7TS/8gGz2g28O14e5RS0tglQM
Uf1+LinhwaTNao/Aq+eHiHMEmnTzVze5MJVOYJLqAgWDdD6UvYcWbBTHbXJdGbamSQfG+n7lNICL
JzdW+HVtHFTyz4PcZumEnGmOABj8R1mOatI6llFGiLDYAhUqvt+xLS4DnuVmKPP28OpFW4lJVAcD
+wn355z79Dxki4cPmD7sfHE3za0pUmhAXaeRnswUKn8ZsozzufG78xN2BovfIfEozDz84212s2PG
0Ze9s/8p/Hadkv/Y4x3CPiNfcfnA2vA9ILagjS1j6QDS5tDfkea9m900U7PbpTK9X7cu8pIPiglR
dcdFFbJijJNAW4ii9/Fi7SQ5TXDLGm2IYQvjJJL8gUXr767y9dekPI8VM7fg6KAnNLBFHfNsdi1e
T+hfDBNcqqlIpZ6xDy1rtorSipMy2/BNVRyVbtQlDhiCuRXGzYIUvojT0gz6U8be02Ylw2me8fEA
K2h5tSplCZKZmFd/RQ1UdKtbea6jEY5A/KgUZDZ6lkjJFlW2kDJJb1YAANS5MocC0wifYbk6I3s6
sMJSElTJVsPYXg1EYeXRKZNZKqxxknuGJ6L9JpORLIlGARLKvwt7JXY4e1O1rq61qis0gXN7rCa2
cFf4zvk10gzqoTcZ+tkXtWK7ky5mFSXN0VbAM9KxQ20isLPa+1vu2Ufdh5kTMSxs7a7m+E4bXQ+I
Lskbymp7DpvB46O8FTxtkMpCdNhO4OMzY34cOM5WXN4SnGhb43YK61sjpc2C+GMA4xERED7faSYt
Z4II8HEsDha9ynNG1wipmlwxGkPBn0p7+Ku2YmLeLeqLQS94wF+9PZb+gROmn81EvKO33wSCHbxJ
lIHUhLOSxMnBTYJuqYthmi99WwRSyfOScW4rbdasAQbqnGEoIzL6lEuKB8ubNeUSFSnBWNnQKK4c
dy2PiM743dIfRVAsHXWTVWkFmTeGBqQSXCmesiShD32H6EZ93qPKHLZH0yZFziZMAWXSburuYeoe
jI8FZ8vwGwOLRAZho5Gu4pA0SCCqMFVtJqFjuQrYxmJ9iGq7LrZioF05MOQVFJC4ZLkvvXHEmlgy
bmt0oocCy/CuqzXoHknYYPrVEoSzxhDxyxTfvLURxt1nFLrhH+xCkIOmbIuwmcYNfhRQD4g4Sfh9
c0s7P2eBc6nHx4SCzxOPfQ6MJX4MvzKEV37N3Y24P5FJ7O69XjJgQq6aIdFkli0jemBZ2Sv2hLAv
ZLKfqlUMd1D6mOoxdePLb+uEFtN226ZDbnwwBoYfOlIZZniwJJLXa5LTQf63QXjxILpdDcZMwY8C
ksWXRI9TClC0ZHxNrLMXsIbMrqSrnEcbUObwgmHXYB9Rcq04h2h1sgn2oHox3OJfJc/zcPfhwrOp
q7lYukm45A+h6FIJOkIxFBypwdpdu070RN+SKKwJK56+6IGsdOOng3gTlr7rwUp0tfUa/zXsOsDh
OTbKRoxu1WGL7iQruIXfABm0HCN0fuv1EPT9jdyXFvf1jG+FE7MTIve0UXJfub4MzLlXjL6kbGHq
6eMGOnEejQTVuouHKagdI/A8dZB4T7XfgCD0KxthW8mLHFODlYbPQ8QI6POzotJZKalDntLPD/wN
mnlUW1MQlhn6KhBV9VXcY4Tj7NarH+TYSWoDVE1BxOEri6Kx1+vzO4FK/eBrDOEsAIX8k9TXxdhy
aJTCGIjvJ2IilEdlruvU/Tf1+BJc1z5OPYVP5onJCc92ZSeVHYdtRDi19JmyT+gcFweKhw7Ht0Ae
NTRHLb8u9aiLaAKjJDSRP/BGU2CUlH0/L/UMtRi7vV/gh21iyToT3aV7JjUoRGv6xWSa0ZW+yxE2
oo9Vc/JQvQphwSGOoHcarEh5ya+CUK3qU6CKLyrXI3RLxf5UPQnx6qTXRdLeSsCBIOvsG1vB3GKw
BDLVVGzhCMAmpAPB2XW3SCSSykOlaW2UJdd7EeWLXxb9zFG6Zcpkp/s5FLgRlGzadMvNGTvuqu6X
1r2ulviczyvCJ7x3xtk94IM7F4y6T2ndk6ClSOIPwMcwLLLSPeLxc5iMun8p+tv87IynH4HIk0ru
4ZiIwDJ2iQzr2lYy20C8kj7TB73qp35XVamO2f6KtYx5tda4s94+/5Uy95DqvCHGGUghPaQinGWa
O63BQX0jG3A0W3BYhPj8epi6qQ6cEYgCcum49XFJP3Not57RALnn7MVWIjJPyIOcG+VDwLdfSW8A
gPLldN5wYGX9G5caVW29VrXa0ud/iFvsdCFVBvLTl0JmbvStVMboJDXJFIBOBm69kBntL1/uohqw
wpxydLijjhdOo96VJGI2TRnLaZyVr5akhPphDLLH+6Jglc89525dQ4pIdM2MqotWVh34QjVg9LLp
zlg5bRXkQ+iq0b+MiEvMx6E+vTmylgFbDxMreigH5CPLAlS5EOSKxH/uyDtITKFvIqYdGEloxUtf
yqNZoPpD+Vovv0PcWnfVyyRFndS4IYts+PJ9vWybePWh51hJSXeDrOdBAyMe8xWy8xLozAuxUd9V
gwnEmwmIFsVqvmgXD4ZHAHLwHkMJzYWl+AEFmwSh0+/af0WzSWvxi6SQoYWI445Dj3fEo/oFXi/0
AOim9fp6yTDtFc1RHnXaDBC0lOqEcchImQDinHQLwx+ZCz25XszIgkjq45Xygt83UU9DHIzc9HOd
wFa4jr9LD8Lbr937Pc96YKxp+JuVCPduFWaG/FILxLQIRXT7u9+Pb+hcYN2Hb3tjZsbXIkB85HUQ
odCU+Q6bSbsMhBt7rOYh/SdF6AQPyT9/wRrsHCkTR+572IompDypx8vUeyyPHKB3AHGEvRScmxZK
ccyyKM6kwYwI2wAVf+mCcF85T/O+gNk7jWm60T5Zx4h58OYp+E7L5VdzHwfHf656s1l9Iq6m/hk1
Pvo7SMnW2nGyCm4c8iZHmeSRUCjbmft2GdcYE0qIfywRbql6QqmFctXaR6WYN5af2B/gt2o1T30Z
lyUdZYkRCsXYCXITu0NEpfJ6hrtjdNFsBQ3jnnN/ZjUldTIQ4DISV6Fp5GPQP+qFizJ99SgXrarB
BElSIfumsLDUdwGKf8Lpu0OXCxe8hpGjNb0sb86OEoY/MfXObOprdsia6NqKOkzSzCjZDMaa1neD
rdDCi+fiPAW1ApewZcbopQmYpOdyJa2asCltblTvQUOU07zOyx6AdfIK+mfHJen8cX08GZsES6UU
Gw5U/t1IqUiAMf+Hu3PY9ZLYv4dOc8q13D1pVVAapiUsuoqtbmOqjQAEFgP8cIfhlaNxPZyE7WvG
Dp80tsJGMoRO1PIJS9UuKD4GH1Ww9ezs0ZMeW8oelLTEV5DbhC50BKitk8uQE48pPs2wbprYqcno
k4yarFixI8WHSV7QGRpfF/vsDpWWzpEbbz7zff49CHmd6tMOIVgHmkrdzDKFybtdyh0gPtTPzJy8
+LdlX3ZoeU5UKUg5rVAoYmmhj5Bsvn+5j0EB1wKqdtqsXvc358xpfOv27uK8pgA03oMTDEEAht74
UM7vz+RVQMtyfeKLyoTE4f4STKmVAoaVBJtwtdhl6nrsklYcBhU2wn2lMmAFXtLslwxd83KYGnTZ
pvw/wfzir/doNgnFnxCsrY9bqb8SQcDckgs+JvmA767jK0OF+ujE1e89EJC5zi+Q0ghXcW4hO/c5
PTb141ml1CIkZ+Xpu2A0XDSHzunfVQ+QgqJqQ0S7C0tj7DDn0yT0z2a8+6ppiLvYGj7pvuR7GkeH
AeLJbNbzjIPPJQ552H1/JglQUmswtDoFMXjlSLcujTNF5Ro8r2SY01iJHG29utKBcxMT8fhuoM5D
TTRX6G+hbni7H/nnpLcFP7Vbwy7xx8+3vkGpwpCJJFMDanlqI4CeOmJjyJ3eXBNwHxeR0vztVLEH
hO1rDL/N5r5WtJBzFsNZdSoX3rRd0imZ+2pnn79V2f/kQ5LTfiuiXdMfqPORrUdm4LjYFUj/6uUi
VhMYfmGFQzuhU+q9CFT2AZ5EblTkMfhIe4or/n+9PUSN6fnISD8o2kAMkik5D7zoZjPafukrik+7
Gorz4gLDHpG6sR5hH8PnA6XcL7kJ/L49LJtn5ARdMARPMV+nQjDtntDDz20kphMLkRGFxdXZuzv0
rYo7CBpGf5ED4T3wrCNkiWk+VBFaGKZKgJBEK3Zt1+2E60O3Nh+/p3OLa5Norx7x8Fi7TgbPqr88
geqFRUj/BH+D1MEgQEpcefLbqgmbxnLhFTvMs0Uvu68s61nMtEapnXLWF8f/AkCBnPJFd8u6jt0p
0wZh0/vsIcA12MtpNAReWvkR5Drt7flyjqkXp6It2JBTgnYU3oZCj4yNGCNo+IOy42AmGzVwyviK
7LP7rPrMzY2pFMQyWBD3hcCEpb9SsYk2HjxOYmLYIhMsoPQp+MuRZztblimz2EOTB+xdmcMF93pk
gShJRKU2z/51hhnZegkufRBGbA7+Y12jVQSKMUJHJPGeQpr9h17ba+JMudehGi81ADvOGgrRMV5Q
RnJLVa/Enr/cq7U8cCC/5eqjoKMSs1EmCqc5zxjAhkk4Mtwkz/o7t0Y2uu3eu69TSyIxp380G6Ak
aE8EkGJuZkWPXEhDrOT05Hgl+1ZAgor8CcsOMH5c5uYsf7K9BevHWPA0e8zGm4Wh/BAwO4FmBON2
0yFARrB6/rkpEeX5xhw9JOldLARdCwNZOAWnBRCKRl9wEgy78vBpbx10nB33Belkt6T8+z36iQQe
rLlTSnrq97Fpy/uA1Db8dZvKMZUwwo/WkE2V9kLGP7redSVu3X4HxZtLlhzrLH6DbQ59YDEVvVT+
7EY/PKapCqkR+2T1UUWDMEqcoCP4Kr+fCq2zfv/Pou6CYNCjoKWQt5nNiiU8tJrqfsje5CA44rGo
SzQDG2VvVaU6WQC6XwF7H4XrE/qFFmF+7bDQhMUOupkmrGlTclptVGBD/C+F6HT7HsVvh72l9z23
RfnCxTuGRuu8h9sybTYAEUHEwabnUmelxv/QCvQ36IdvaY6dM/l7AcgTb84asvpZe6da6EjT6FUy
0bNsDe0B2gpj1e394HZPSaFm2fiz3rnTiQBa3QdDhUqRj4AixdzjRW1mC6f7LJ4pnUJSabtyFlUg
/b18ClyDus4yoPjIKnB2l5vRw86d1AGy0nJ0Oa7ZTylIEF5+D6FJ1gZyvh9pmKNiMTr+Sg1kZeee
6N7Hmbatt2Eu91D2ndf4Ov25HcFGrlKkfPswBlITp/oYPsNlybJB1V0bGZT/2t734fMMROI1S9WJ
4k2hTz0UZcCR0k9bFpqtP+BaddQ1xU+E4gSBK8RC4vbzeE59nFIFZ2aQc2IYhnGT+YZAeSGsnuUK
5jtZSPPnOaXDusJB5Q1Pszp9dRdtw9BQtRITzxYWj2zMgQWi5X3rQi45qL2wRwpNfQ5LiieZ9N//
nWukyCCk7lAWDdbq8apKGyhoV0qjvPKk2+drgu2UVucgV4AxFZI5wJDIa6bVKWQt1mMD82n8e59A
XpKH8vx84mMFTYPJvdGq1rWddbT4EFxx1f2h8Pp92TMkuCzNuwH04WtP8LePYIIzacLseaPcZUHa
aiXODEspLzNZi70ACmGADy8nd6/YsVo+TB332ko9HscmNujCw5EKfX2uKY047VtTrtnS85aG5fZ5
UloVv4Q9jA17aCKEqMlRzZVCiiEDlOWTvanBgqUy97o39LqoNIn+ojL/Kx8R/2zgLyHYxizNcfK+
7rdWh2TgK/MP54brQFx7TsbcfgA6+l2sbjJ/BFTpGi2nxFUmQZ5vnKgTI3p/a1lt9VR/8cQHcm/Q
EuYLNnXFvSCNZAMxvEzwxejKSHVz5rhr0leu1xQzYukn+thlHCjON9oBiVgZGsl+7xZJuA3HarPs
6Y5YHAbx8LuQvZqe1cp1QqVu7Dgdk8kEwKMKrwjMRc1FEeMdlmtcjFvXQ0iW0xMRPofYncGtX8EQ
MNFaa7MCU8cUXZMrKTTxjyyIPKj+ajfB9/vw8YbtMGmMpqjkEYdVBLwSY6zFLYi90ijh68ZC3c6o
cH3J4W/TAqR6ITbuyBNTQVaTUEpm8zNgINjbAdyR3VQSnUMstmnp2LDFK9ibPCt60Nqp92xTSDQ4
ImLqte/oGB7CA12rs3hUO78lIjOiPMoz3vfHcfUyLuLmjjMkJPdLqxB1APvsyNdshvDnNhn2lvbZ
NBne9z8s44qa5Xzkmm1q+yMTdAyEMGJBzd1JhUTvTn5NgXyFrfMxkObh8ABCb9IYXbgxyZ6Na5Pp
xsOsROkat6DYEwJXSczRSxMvqzljIUf2uQ8RuUws0HHv4l3ZZ+aPV0U2dLrhUwsgsklYCF8uoz8k
DdWyIk0hr0IIBU+rgW3FVwEPq8SnZKpT8wQWCmycbZ4SVxuvgSVK9deasLpkQO4h6XCSm2E7BYu0
FxXbO/Jzdfi3n3H6pNdLwGcy+msLS7MRiSBVFXaytxAkIgVfbGs4B7FzB/SkD1t4fyWxGGqcOl3I
dqqZfBsxor+o52wZc4csJACO9WV+/PCIStbSkZy7JT5sXVzDdppOzJ/YtDzFndLXVZ34yPUkTYHZ
hEoUv6yTMHkF8x7yMg0Acr8FYCw5aCKdcQhk5A9go3bZuh+zq7YTkBM8qi6HGRVhY2fgmkKpTSwx
sNU0ifvuUP6wHrxfsMqSb+P+REzcTqZ9CwRLImrjMTXaYlEkMIeRI+VnM3COtxehH1f67vQ5znYr
DA/3a7poz1XqXwC9pzmItiTrMgCWIOTlmDGE5vl53qHuntLFZDh3y02SuxTzjGBqsnYRcRS1tLDg
J3QM9shNFAFnwgcuIdyOuWQ8XKnskWGBIQ+qoyZ99iE2gLTLFrAcvDirofkPr+ahxKHLgZTp7G88
PKo71aSQXSMZPtJpkzy1dnEOvjhxEafD6uQuEEVE16rNKRUrU8dDJN1FPh3FL13+vZk9WUPsUtD0
s/Xchfou8HvHT7tulmkKt40ld9yOEA2/odIljnckE/kLHbWnn+xFdAdVcr2asDc5t45hLk120tf7
HzTWRTckr5ImN/4JB6Q6Ar/s7LHveJg9F5Vh9sYJHgMJDVHKuoD7fRt1gZIXQsBTqN2GMs70jcZX
E0ELrcxiR/5pjevXH1/kTmWoKb3lMQ0Q+k7TjLB/QiMtX8oCTTp/pSmT0E+43MhrRJufHIqPT0py
w3GjFFwk4iS9eBI8F1crVImqftp4SOa0UN9ULa6kg4eJ0czTssehIsAdiaLrZmsHgtLGp5aVozx7
eri7ZIHz9bLe7OYpsFORWQ7/JGqa4Sd2k4QMXmKO+FOGPVpWfJ0MPfNXlV6qLOr04V9+eogRmt5w
tUWMUd4N37X8tARRbs65iEEQJ+jA/k0r3V/2D1tazehJFtNhGLGTfU//NxVqjW4iSU56P8pN/rSf
2PlSQ0KLn8EKmo+A9t1qXpFHVmEFLsMQDrA31gYEp9wcmEWpdkt5IWni3IiVv+/WPrNCWAbMAq6p
dpV6WkCcfWm7m/SKtara8pt31sv+SiWQIEyj+gCW3L83oSaSjPlThrVveGg/KDWcYH4TgIVLv4h5
32xqusuvH73dRQ/dlIsPeexPwpgeGdbAYUwufB2Ksp/WC46M4d7WwCk9cQw6X9oWd8WoQ/LaJNRr
9sJtMHEQFOVPDwmbQcSq/dHDVCY6p4NM+3rSZc91o0R4FrGbf9dF4qpisd+E4e/S0m5fB5uZNK2x
Gb4sVxH0oGiYzSm8byrjqgdVjzSXZri4QIdtJDVOPF2cQFh6n9OK4oxAzD3LHvnae6YMRGSF3OoU
WYRal83v23V6pO9jOU6hq7kokBrA4VDPLCkVIVLq85dsO7C46Net6dKXP/vl/+IwVl84CBEcKUMC
4DNn7GvvFSHkYxnOGB9nXUq7gQFajb7hffDc1yggVPNeIjamP4A1kp4ilH/omx9BwzCYTcBnvSuz
BAuSZeIGSHg7cMikbBJyS4PEOhILpO5tf+cIBdQb75V8IQ+bKHShkoaJ2Fz5OHDudmk6BWkKJoVr
4NqRgd9fHY24gWdoEacGpMSvOkXXjBEJYQVZB6OqZe5jZOUmXQdDNWxbdFvlSGEn5cHo7J7RuyNQ
d3UBtv0r38uZoGfrIvglvPUJDiNb9zwn94a68qWh+LmV54+i56NoFohrdggHSv3aF4QL3GNgKbym
Ys4qS1v+8dpBa0ZftIOo1cjO3g5NlCB3KuMKZYqZkrWs1ZSy8LakEkXI86+46qc5jl8En8oZzu8q
XMCMpU3Dri2Ty6HWKQUs4paQ+brt6QtdAoW36lWrnHMXVcW+h/ycMRpEptfcAECzesaEDqHc8Dqa
HObo8ic8lPyV5sqd+5u89CVVn2mfDcC4dqGAAIJAGNpyZ9TyRPyOnkVyVjyFtx/RrMtWj+Iaafjl
sSGb/VLM0yPDShzc6BAM9B/6ibbSk6ohLkO3Yy493c/BgcYtuDX7LXwHCxzcmV9cX6BBRzTUuuIG
gA2lVp/4thT5BBuxf//byPRRDi32Zg+zhoRBZkOU2cUyaPoo3O97h5zWTU60tWBtUxcTXVJC9PE2
Sx1fkPQj8J9D+PuYmay/Hb1hURqyMCusGVC9hLPMukExI94RpmEVinURb3abS+ibzd2wyrHo4ymB
cNhlX3Ea6IT889HnWNzBIjoPy27wW1RpnykMvgzB/xlF5SbbpiLSjXEAb7e0emtoWQYwo0k0Fv76
tdqVKWdCKh8v2CD0aKPq60sAe3byVJG6sXZ/wF4fu0X2Z5AotDjjkgDzCdYzZ/LCvL0RLfC0o1mQ
L1PrpCZ5RkkF0lvGEM6a7HyceNzG7hnmrJFCyJGpd9IIkGiMK273nZvm/GaVAPwZzHWHc5CE+Rp5
EoFmI7+cwGwZuN1yq1CPRHYFFlTbzIHok+Lm/wKUv/1T6CX+dupncQTh2zkqAuBpELCDic3D0eIz
SWT6yo5AgddWXMBard3cHgU8a2NBun1bJ/BL5lNhZSzEx6HwcKqMunG5qC8ei0PUYuJ9snYrQdRq
wPe1fpXgGDXgh3eTukrgiGmwFINjc4UUU4hCVm/3w89Kjcsfz36KKD7T90jTER+KWUhEFAEGbzAn
A/3Bk8AAMTh+16T9t3YToswHEg5oxJI6UboZK3Y2itrhWcibs03daCQqNIuWOShUPr8s6Fd7JTbL
hdr/2IkQEZnCJSYQNe0odjtlFebvj7SE0j66s4rgjTOsGIakB52osR3GaWUZDDazJBWhBnlIaW/i
qw8jAcw5KyxunGjOfZ9Kxj/a8VbYUect//meF2AflBPaeB/sFBkGpMGxluvZII71NuXgqDsMgffo
8zhAGrklQ4hrsmFSrDWCgst4AKeuMSqKJfw8Au8zHTgEIe6MewArSFHjf9SjvHhBP/YO1CTrFJbY
9pjP6BXlD21KPsNaMt40PFlfG+zJ79AtI+hq18SjrQ2jyh8syBsxbZqD4kjX1WODXkD8nqGuqbuZ
pemk4JRWg2FdgzpFMVAOeHne7OUqnmxbULpTH0H08oGEkOCV1RFvW1ARLOrVkXWofzEFpL+io7vL
grvfVsMQmhbCh9+1QJEEAAn0u/Ev2ikFwmSSYAi7b6/piX6VjotOXobhDoV3rbC6uKwLebjRBCcS
qGxSUXdb622VHc0hzq6gPQVUBeSqR2Kj56df8VBl16KekgD6yHE1tNmQK+Yu5a3IcgJPej4aZUd9
bqpDrVP1vGFNJU0zRHLIde6O0juneLuaIiHeMthy6mC2TpArY+zew5lr1sf4XyeyWgPnt5+vJG1u
dV5BB1pt5lb2ePN3w9Le1NamwyfbY9qmeZp+nWdAcPYjVuWSSblbD74xVSkeml5cKK06urN6+8q0
YbjR/FUz87nUqjzUUnPkSQwxka/iBEgbYBVi0iZqmo9O/msf7Y5u/RoFPIkDzp2avBUumwB1K5Dc
HBwuYjEVt71pATSdjUUYmCoFwoHZCXh3UyR3+m1GKYu8qGw5lRO8By938W/T+6W+6PfEdjNx4dYm
Fte5JMq0NniqajU7YlWwd+qIn1M15+Gbw1OeOtyPAsmHcTx33PAHCcoO5sLZlDE0PCDDZtbs61vb
R0yVhGNXexAppFENUipSlCSd+ZPnZ4GkW71t0e7LjfpSgKrJIP8T1uPJTN5tjOlDWAOK1SHMKgA9
41lyeHE0zWvcpRFeCbBEVezm4fcmfnISK3Owl/p2BWzFZuVTr0Y72xLug6wNAsT5jQrf0m6h+y06
G8vtqu9dvcsJuJw9Moe6qGU3Z8wECEUMVVDpn9LnhSs56Ia0zanvjR4W8ruotoT0/+X30sNt56Wv
FBeOY74D0Y/8BapCa68g6fWBM9roeDSHhZqbMsctsa69GrB1mWcfnJm7uRk6siZGQ2CTAPk72rpb
hs5IfwcWCQDCpsuqGGmNU0QhDy46JCfEjMWzKZSUESzOJCJ+ufcYGbzwSNKCW9kUW7251ICTt9vm
xHBuLbK+IMEPnQNEhoz/L518fcDXhnB1EDvgfKPtFKKVe+vMm31LEoKP+wJnXa0ClkxoLkyYh3hU
xgeLQycDqpHGOPs+p/dCsO80RJsEcs4qp+DwLp351MiHUgBH9WAeei4X+YFQuk8/nFH9MYVUVgH7
USpgyMo2a8847V6dseSVPZeEP70bZ/Y29veuhiI1h9xSU5eqfb9yQaRoB3M3owpOZOMSOcR0grEl
RO+Y52oKgkl3lwP5jE57t5q39v/vVEo4cs7uowvwFVdt8nW1QXt1491LXkV/Mekdtc5NfRap1J9g
Exe90cRgcMs6MhgW+CvQudFVqYWTp96ARkoUiKSQdWfcs0L0/gqfGhi/zXovx+zjgJXDbV6iPWxS
wDPOL4gtB8z+oyhNg9sUhxLNQ1qIpj5Fzj4XIurYgHLher226XrWAobWKBYvtzjcP+NtsuUHHtDo
GeayK+7Kjw0NBOkdO2TmRbu0JRdy0fZqHy3a8COSBTTsWESzLOO5PaiIilUeZF084KLuKhXkCPTk
Yg9IyO+SC/ieVSyyUG+91X+APpuu2i0/ocdmoIGIONiW2sK09Sp2IVx2ZqtKglGxdZSua8ti3dN0
ge3cQylpOIUZHSxXET2G6CXl2DMkLCrcn+TLfcTGz5q6dVp5u6lFwed4xJF34wCnuF7hjdgpiBSi
0F5jyxseOGuwl7v1XgCMMgLZrs2i0KeH4pEtXJk0hndhF2V9/Oz8KKJ3gCu/RZxIOOe9RywNP3I5
sxwXxaATZpE6n1ozFxRKKFGUEZfK74Gj3nTl0pKEj2MIHNfazyFQWmX9Rl0voUqGxX7VVnUYYDyu
WSvjftFx5LQ7FRvvaD3YklJvydAfKj6Y9bSMqTOseUQEO4G2ijXM4gwDvb/g0d+MceW0gngPfNkD
yQbOsPce7w7KuBJidQbnd9Gy2VShTz8DWbr/MXtUz1Np9hKbzA4rUthlJfA+EXfulqXKY88kYtSV
9N8L9KmJfL++c+5mjxi/oHldmhlgm6e/TVI49p0X78p5N0t5T9OoCl0jBY8shdBokr2zRA8gQ7Ii
nAVEbFdYxF77zE9aXQK6fbIJekQqxbT6O/QZI+gJo2aSkHugYQiC3xc4BehtWjHw8Kuv9v4HlB2Y
jyrvqbNqYoJowjmQTbkcHYx7OsW59j696faUrUeVwIVyNEnywgwZNisQcxNK+XKX1lSVyD2X9Cbc
dQsRtQxe58vJ5XW7+ZOrSfe1o1cX7kAYpIqN1RSwIEybfmFsiNxBSpRg6cspstxPofjJWsr3snoJ
K5hMESTFAR7FMsx6L4miP055hG4Fpc/cmtbFE/CeW8GArqKb3YwSsg9hXWW2Lx59nTFzbTPbwNzt
6xRp070kWslNXbVg9mX0MpQFvJLLkw7tG1XOMVeozIEwH7c9ZixCO7ePlUe60iQuC/Jqqf2DzSqE
i9z5q1OmPpwl+RY2fME1HazhOAbUfOorzLfHL0Ns2eJlH5f7Zt66RB98UAnp726hCxiasFWPxZ39
LiWy8HDUGL0Qw5Fmh4d2SAckd6bWWU1DBiM4j9m1BxiZeEwwHvyqyoOvyVLeMykuiWGsUORvUp8W
RDT7sVwBvw7wntGADzwEaO45ZCb98tQL+2MKzUG9Zoj4icSg4ImbIn4E69B3o/4hVRGixI+dCvzO
aaeMaALa8t5IJcyKxin10nozZHmw5ExH9M5CS4xDxjYSc2gbR4VyMUj6/vxfHPJ6Rukv4JauNdQC
/yP9RYKzqeJ48/mgaKEeg49MNolcpJmxytstdPWtMjUrsgZZj3iFboJtIr+QLfp0+R8iWMpBaKhw
XDnV8aaAAHA2r3sIGpmqVNTGQr3RrOZis0ckVPAJZUDTvfx4DJ6YIOfSxncf8Fi2mgw4UgJ9nonv
UcmndKlIP+DU/AW7wqyqB/6S0Kw5I8Mcx8o2Je/YRf5WXX7LPjtoRzFcENgIFS+4QQH7EMJGHcCB
tLyL3l3yrkggJAH/JYeezkYa2Fz4bOUD1oEEPzcBQ6eBsT5OK6cA0MCLMcxzhCXJCPtDyTnHxdvb
0EhOoPjSr0vhwjnYlgERURbqG7wCFnaaFusQp1fuy2wZrKq4xddSs4J25rLCrEuhsaRm7YWh7FiY
iz5MA/ffWOdufMf3amnnFbSiC4s2t574kDiz3KV+dE7ZKMCx/OQQnDj4p0DqgSNNUgtImRUWxuR7
Mw/13A7UDCmVLOScnmPrdyc0oNCVJP6l5OHkqZMVGR0TTi8wUqCrHUZj29zOoHPJ0z8TOZtIpIqv
o/Qdrlp87mROHQfUlWZnTdyH77DRBIjD/75FBiNeRRIa1KgrrlLFDXZbz731D39nZqSAtJfYXTtB
lIor7ZTByxh9YRZMeMyZWLPN6Wv/M1Ph72WSDTjRYhytTltrrok6E4zHYFUc8+J098VVVoFJO/Hl
X1vEQu7G+LWAy85XpcDcRGFYNb32UW1APm4NqkylOYbP0oKlFx3DyiJRi7RfJTOuBa7OQ6xpcN6r
tY2cR7zDLl3Eg0niDstOl5DdgctC1ZSLHYOl5HBjp2qpdTCRaWdtl9i+KYuIR03FH9jEaXqPm/g9
x+78EZZ+PxuLRotWx8LbG4oSRUOfdv+5aqEl8WFza+OICfK0g/+e0LOCeE6HKYPb1iRa8HWtiUZM
DTERqokK+BYrDzlw+EzHNHCBlKaBsmJqJhAwk/sD2p0pXBXx0D6fGSrLJnlH1uOmA8wwC9frCQna
/Pk7KdNFUQ0QfW4T7r3XMH/WkjyBSZzJ6SaBRZun5CAB2M4oQHKsVBSfAPIiWLDp6Byzvrs0vn1E
bg4OopIlAUsLeW5PjPnlTekkIjfWwqT/Q3/dBRQMRbGwZjm/trbDL4J+e2AMppN5TX9ZS0D7hcHp
AsQr10zZ2tscKlUA58zwaPS4+cpwEtar+u7sbx7W6tVlicZeUWw8+1XYCikVnmnicSSHHGwmSEKq
h0Zu/cc4B6KAxixb7trNPHYZAgatrIu//B+oHg2dT9Hk3KrTwRf7JEeRwflUqyEvkp/kZV6wS74q
SR3qyT0ZXNVtCPq2/QT9OS7lr4gcvy+v/6d302z/UD9dteJc2bhLSU3W/aa6Drat1LI3oG3Bpidl
Ate4bX6PEiTcrutFlGp7XDH+SYFJoE1ywtXvG6cph6JddiS+CwAYP13gIhXqlVVNsvJL1zz2VEhh
NpKTx7vp2TmKOUn/4c9AZeKPWWwLsNYt5Cj3ey+tM6AWv3p9i2Qilc10tJ9xbv/USN/OPk6/qVwU
e/bjG6UyvtKENvfflSpfsim9WiDWI0aUuBPWUvG/JDG3jt72YhRiB0xM47YRyokqsqRBN6uCR4+W
+q6lkVJuJgja8CgvJJC9qk3RlHnJkgojq/LFmP7a5BBhAlCI4H11mAtrg27eni1sMqDfZSWClUio
MZhCIjVE5CTQffcITCnuE576JFDui5TU/oSwLUtfThmGXe4KaCsjQaaqu14wkvdg37P4vGHA+Exq
7U3z4hH+ZBbia5mSCvS1Etww2nZspRO8U0LguTAGr6G0jUWUERL1FyzwFs917UJNConFLet2FClr
pkImlybIgdXdBaJwfvyQCNoKCc/6M59zwKFVtMNTWaVLng+EvJZtxvRfp8SPdz3zqK7r+xylKhiv
fWlOllISlP+TDzporokl9J4+huiw5RlFfvHoqOs1ULVQToCgS/61LHIsR8lAHUzjJRGT/wDZJKAx
KTPxURdZJDyxRs8HMYoJbJOCrdv5F06XWIB92qknuMAl0sAGkQCInLzptPWyJ4GVI5TWuxlfWh3w
g+KkUM7cgIfR60278OndV2Ogs1H6OONxkX5AhXih3ie1++zVGWjNpmmKARM2jUFyBrAxZJPwhB1l
e93CdGniGhr4iNWYKaJn2LBDhhZzEfjz9iMw0pqdhGoaCsRvEtSgwLNono53Yrd27HLSxUqHlrzs
9Qp8R/PcsFNR3fOsCfAEaWWVeVR1NKcwDiQ+Kf5B4QAMlI0no71EnkIawHraCuuLIkWzAFhAyXkj
KzZy/cTkCgbgxvFiIG2S6yLH8Q5Rp+TbLYjXO2SauuQc0YKTP3yVnFvLpcTJ3Lt//aiA/DuULLEu
ldXbmmHP6jxMwAZAFD32FvatLwyj2igWAt14xl/KAp4a12LEfSWBUTkFhNvMK/0JmsumfcJD7fXU
dIfms2UvorBffLKF6nmn9+JJQElH6mzH5NbvydzCRokukH6k7zsMfKIN3IXJTs2KZo/pf+tmfYsl
NFln2htqwiZumGmX+K+0Bva7gpsWxAoA4TH7SE+bZHk6TAjrYPKzYRUAoHxZZ54EC0Udx9fsJoov
AcMxhVH3uGVl4uQN0bpryxKcUauUEF4I2Nfhw6GUJpdyKxr+YqVY+Z51RKkjb52cwtigle7hLpKA
5d3KLbaYmzAGIdpOYH8+bANyLDZyhWQtEkhquhTf/UAJHlAFJq1lgNYAbJMfNuqeLHQHBHGhUU69
NNq3K7eFZrBY8d989LllISu/VlWLqhxmc3V9XBqb3XDvoIs2m03JAe1jCCV61u2BQvdS6vCDWnUK
pq++CsTfFPj27nFN5r5UzGnGIXdN0kyRhdPScKc1rHvpHuKneNfG+qMXk2jP6MCfggIcnR1xTL1J
ZvGuNS2i/kSAs3mZ3ToruT8mAk1e5HSVwc+LvHMEav3WiWj6G/8FdXeE38F0lkLFfkI7hHJ7Ys+k
BjbCKIdUqTRDyKhkTaiaW1yt17vXPhG67a72yVLQxcIOmeiIKPGGWsE5SGGYJVRUke+1YHHlQpuS
mepFI5VrjtbkKQvf4JJuw5wGeZz8jVMRWQ8XS/MzT+qlC1XBPWg+TaI6bvFrhOG+S5tfqGz/YldX
XVprV7womfKgbwe1x/lH4re+7T3DvXQmxVtzNPX8w9I2YWQACncxWl+SJuH1ORW2W3I5pxVvr+dg
y7knvvfXGh+tgAqeXDtl/FE1Ki6ZgTJofzE4jCPO4oSUThtIyGN+EHmQ/EW/e2/iZG+K1YMJtrvQ
5icUUNSnG6ATZXlkhKfnNSKixvLk67C3bSjj05NdfwmAJ+W9cn0dHQoIXUOzSxmHqyAQ4QoViDi2
giM4hMySD1YuSSscN9xAX7rWcrvM3hOhYM/2/etNOFtxjilmN1Cx5724oap3yLhgCLLkFsP6bpiB
cM/IpXcgbAGG9BSGCYGmyljrR4kj7CxlXGBB3Ha9Zv3NQ5spvdVgtq5ABx3fTv3CdgnOrN1CvFRG
dDNbirB3vgV0H17LZ1f59NQHEpBAhEkvIuOt57eVzLZTqXE13J9tCbx/Oth53IAhc2/DhjrJndqb
5Q2kMX+apyC6r3ZriTGjJFjX1RZoLk9rNG/D/jCR+AmHqlhr5FpGqwyWO+RGLuN0tc7PYzy+tXO3
FVah2xY+ubbhVf+VW2jgz10o+3/6BTqLfq6ZqZR8tNg4+g5SEn+N6zEk23OVUJDRU+kwFL8hp64o
9y1KJkhIZz9x+/i6yItOp6E3uebiBBV/4nA+iMYLTnGZGKk4u3x0H9YrgnrymefyZMx57Vd0tCdH
XbMZtYFj7wFnn1aMr9f9kaUm/K4ArFdJ4XTEzEvhmLXrfWDErEQ4Sh3FftrHVigLWqMiJj8qcUp+
OezroH10IssoMJL7OvkBTvQ+iGvG9qKMXyqp5UtztrpiKEqt5UKxWg7fF/rRrcTyb6D9liRy7zcz
0flhyX2fFJC5EZIcngAGyiP54Q2MHPYAPHbYkzJH4i+aRhqD63OVWLySu/LFxra9mJZGZ1PMe5oc
a52aq5fFPOncvrpK0+ZwWpBwDssEmN8ZzIRqj1X92HCrq08OQ12OC4PuTtIS1sEpDr08mOPshcmR
2DsBtmeCSF0Cw5kVewrFCMNd9BObz8f7jegZWUhzYqFKmxtHrSyf5BxWn03LsxjZkcaHc3j8Ijuf
3bMF94OOHf3QXTxx+02br0sPm50mqtrsIIUuRul85P6QSp0qGZPe2aR6IOXYXzG7xvHIRxUjv8uY
IYEtbIGyvF4ob96FvgC1HCj0CMzNIpRHdvreSUE2UCWCxIS4qS7D9RF9W7sCGBEPrhL1bZCiut2d
lgzXq3BQMIiWpeeBlxg32JLbMxrhZDVT51NW2D/Va41h93hf6jjgVuqHHaN7DxnXSvOv7byCsxeN
WJ9lP0azv614LUg/ZKBlQfMTUqA3HZmyW9E42r9fxo45QDwDa8ltPQQ7GQg4ycPmolqM2Cq8T6TH
Uybye5FY38N9BVgNtOlapjJn0/UHcoAFhaut7qug5Kp4axQMeHw1dEZN94bDuFQbRWLTQYeB2pTK
CGgIU3nDat81XYlP+1h3qaQQfG63D2s6dL5uVpO7NXKIsZ/UGEzCQpvcvDaImVNAw4rvYc49aYAl
05zUb9jrn1ocvWS+IpWDQRMEJOK2t+754okU7JW/q+xeMG42vHfq1s+TktDQMFLRwk5OadYZlxRc
JOi3dp55/WbHQgsC6iOyyYYSz/pWxL1Wu0l4q5t5nceot4IyQzAO+IZciJ1PRkw86xGBLwPe+Ro9
ZJ8HqlGu7qjiAUcRw1Hc8aYbUBnV1nIcv1Exg3/EGWl9MtQWLiCsJ3JNRmDlRi9k68UsTPr4hT/f
ROiJoGwJnB4bEuWw67Rpxqvih0sICzvL09aaK4FLO886qdE1a8y4BfnWgimslbm1xK6mIEklpuek
n4YB2rQTUuA6O8DK5ME9AofzynA+cHY4xorkv/MjiwuvPuXcmqjoWIedgXpqi2woGD8qzRQP9lvb
Coj6tdHpEflr3b7l6ehMv5Z+qgq/40MWyvJl5ySGCsWMpo94cDYdKx/HnV7mjEdh7UKghY9amTcK
nP1tZuiV2jy+0oo0up8J7Ere0l+R9oDgFyubP3eJcEeAcwYY4icyKgLkQbx4D1OlP2Qyj86ToDkV
c+UXwZ20Hazgc/d/e4OxQoOWddOAY+dAcJzfALBHFamH+lFEjl4cpUZXXhWQT22YSygYe9q5nZKz
1srxHSmdDObOIuBB80aciUQp+A7Rrn2HJTrG+c08Bw8WBlTMdYTGwdfpjzZLlEyL0s4axTUvgQgV
uxFuppBz8xl8wHbx4TxIAyeYBBg1nMMrBa6EZb44zmXATreh2p61e/oIUBSgUG0AsuqtNrUpbUcJ
lrqA8w+zpJWluWHNkZrVGEVCxq8+GbA9nO89EvROWlgGGLQvN6tfKyF/W8a+s+kgF/4TC8D0+leo
AgPkccjoexosa3Btw0nuMRZfvEAcn/rsJ4dp2JBC3gH9L2Kl358XEtGwdxXM3ZGXbyU5jmkn1eSm
lM79zWMTXa+880+SzgxVWHmHwDCMkNm/A2tQf3NOfLYR3H1YzfVfHvRNK/1MRENtQp62U4PNe99f
tBdXweVmEgraXfu/Ilmnw5h0QMCEWEqpNdR/DHVSd+OTGxSeXm9vfXD/jsZeqb0AbYDOJjtndKS8
MfpHO54c4A5JZ79txI5qrkyeeWQSNH+3fGH/bLg+H4hfrgtNRl8UPEcsQnwbZTxKSZSPj0+CC22s
SdyPnwyi7sEkBIJ+Ik3d2I/DJ4r/eXdOdD1k6+jos5erk4R5G8GKP+eG1I42xh8a7saf1idUCp3X
gVOSN6JyqLMFsQt2/55BEh5rhHaA7HUg5GKl1SMDdAc0eHpS/kbl9xQIIXdh33WfVAFWZ7SNOb2D
fo1euYpam7EN9lHMhDbC851xb0ClhWyCdCyVbp9QG80X6cPSCZcqrqStwHoaS/CseyFW6iMIkxPd
ovdIWT+ko3gFNm76Ut1ETP/ca8sZdoN8KchSSRpTnpwqk4YIMyuUwn3qtBd9Ya3C7AmHqzCJ2HXb
kGym3JDFgY65pkBk8+ToL4QXIOR8JD6BSpe9ZQUU777KdipYRSP34vWe8+GIHk2cU/u6Us1fNCAW
HGF8HZJlhem7EAw/z4d9WRzUJpWFeZGzn8MO9zTOvsTIH/50C/6YA/XAc2olBzXQzRr8g87XAd2w
PmEjJDrp0bhfM+MfVkxgBvQezv3MpOBiV0ykggVIS1LQoiS5PYgvRvR/B8ZIYVMQMCcvTEjRFFyM
1IaK0ZghoVhwJ7J3XeeVuKCv8dk+3t8HANVXsbyoaBIycIId6y+cf1SIGEndK+KYiuyVacQEQcLS
PyVoIyTWICwkL4otzidDddK82ruzSbSDJ3VcgUOUnpbKl0vo1ZYJzyr58KMwiAQmRaIx1UqjFGF7
D6tHZlZVIgiQg3IT9ANJ+GDdlIPK0rCnlsoFMTg91Rx79Oogh/MSkW8F8CFX78Zfp4iSfuFIcbCn
i9fIBGPPiYdVrv4RdDhCvLmt4igQb60I6vLFcoYnsLLuXdPXpWHGvipFfdqQkRFFaL8qloVdg1MA
l17CLaU/Bpvs4tzJ5nCxT39tZB4vt20H49V63P8BjXv+ymkg+ktgGWwVdQMJlLJ9tuz7j3oO8/mB
yie4Ro10iIxb2YL1d8lgWCNnFi84codpEmbGDaGiAKB4JlwcDB69zAL4H6nJu0LdxNKFZl4kCwz1
4TNgiTnR071bmqbLYV1/nlB3Dndl+6te39y2G+TYYBjvGugP62EuwWnV4O3tXaU0sTdOifPEPuMs
PlYNPY++7xjRQLyiQSGeuch4IA7c+udcSKSUqPHsQLVbVL4OzXHf4mzwwt3evKcbhLr0J7redFq3
Z4NCxw1lDd/IQ9q4nYNOjJwgrH2F9zlXFlLsFaVH/qZLTk6KA5KBe4v5GG8U8zWxI7zFqE2coRuu
uOXcbOiLDRV5bT8U38r8zaK4mk6UGH8bxD1d2Q1nkMrerLBcXJLuT4ESD+wv5DTeVFrQn+0Zltb7
rJRuF5RPm4VSL1/3Sv1Msq4TKHupqgKlKmkSZTxOSRkP3g03/GSdSp5qpLbxZkgsETxwP5amm7Wr
QU63gJoJ1e+GBL0sIJ8X7BKk8VesgRPB/TV9JQyaY5vgLdXa+De7X6gZJbCMHGE7trnuO3X+jCJh
M63oAPqyRTHk0nD4BJVD0/quSAbna2MV6Fo1BXoPZlzumGHL+S/I+V6qXzc0ODTSqmpyFvkM5EJk
1X/t/QDzKxudft55RX+Yv7gKnZn58bBG6NMxQdMqIPK5VThyF0miGFoX8Z+C1FnPPjNelo011Ns4
ij6xRfJgSQeJjKnLAq7sK1qC8Qky7vjFwv1hJmSysCG0Oe91ztv2S2ifcChjYv71Iu3WjOvq0E/E
Bn9pfFnU/UfhOHwJfppSFRGQP2GKN7fxhhhZ+lkWquir375Ya1s690K1IZfgnKH7/7+t5o+eF1j6
AYofVGiB4t9WdLs531KYvAFHFrVgym3JDjQD1qBZgTP3pk+knHO444UXFDY4AnTPAIyj3G0Yk4JQ
gOX4mJuf4uQKsBJrgQCuN49GvCg8DXJcpYAfw/XnQE0DJD1f3U2dLVcHA3ggjCQoimB5BSg26JM0
wDLeDmpMkmWnQHdoZv52k67tkHHISc9dUWBdst8nVn8IJxKoEatWeHIDTPqQrEaCArzazjNi/EIL
fYZHVyg7xEDtMYFYx6CFlFJ08SdPxydXZD35pkH5IqKvWVleUo46KqejqN5j9reTHdorkw31tK5s
Y2O558GZvJ4dHJxSMhXCPKoc5daP9m2IUqmm99B2+Wf3/uBImnqbtLKSdEHaZXbp3xyWOTvN445u
mDhgml5mby3xE3RhuJCVkpZ2LPfCQZLJjxljxG/UYClcwLfuNRzNoB2ptGSvTSIxfYmlFQFmSYpI
vBhvrBQyb3K3HH84EeHrhLLpCX6OvozPe8J3PL45vR9ql6k3HUEHuDraiAX42zc0lPUKlN7jxORa
j6RZBQKxIuetK21JAPaV8zrGTLt8Yz/pluBSV1YXZ7jin4INYMuCzGlFrUbGt6WonmftSefA8Jxo
HkKObUrlbLBoNPWr57oCNrniZfy8qH4QstelVIkCQolrIHqZtDRE9oToyR81hXIJdDyrJu8QxICE
jPtHiz3G7peBobp/n/fKNjJi98+VADc8CiCpkdHCN8VzJXlMfKeNuJwa85/zcAcz2pOX08m9ZeL0
rxMP4eQQCOHtisqBnlwKGNa8mqDZoGp8CENmq7s/ugOy02EsHvagf941TNoveM7O5NeDH2/kMk9Y
hpqNHxUFy3aY/h9MaI57wBOaC62PqnwbK0R5pk+9Zc+lD9IOZi+VEU+y2hA3Gfibo8fFCd1JAwnB
v51MsbjzGyyU70P6ZimOLjcAVAuCiFkjgnnsRqDrb/ZhtW0KK5tgM9gsm4yBmyGPfMtfKYURnis8
HqXXPseV75LYmh77Z8iDLpV8aWiV6Fg0havnlncZNlpHtyMsTeKGFIfpEB/8TwnF5F4mb94LuqUl
81pSOIoB0UxL7ch2V+0IzO7Drn2g34jJLLoxoZqanPrumZWxYbxBS5u5sOd/o9dlgrH5aQZMzkrl
MXmUaEmI4bopN5ZePmCKotb+zHdfN/ZNnZlG+HbXisWVeoSkhdcink+mBCtgI29iU0lmnVc06C7B
HnFfAFe3ajtrVFTH5DhDn37R1geiNtMAV4asnlpJW21PDoYV8MI3CGTMduts5104EKWXtYtVpO2Q
hoEqfGzUElenNyNg9ER0qMMIwsLbsaIxv6LkiJZsgyGsmrwqfHm7t9z05nTZZOia6AT99t1lc8Rl
xK4OHR4UE+edOId0DR5N34AbD3DK9Pa/rl25dXi1BKWye0lZRe7Y4px149JOWu6o6HGPLdGhdOdc
i5RuOxTLUlgrj+0P3oKA5MD8kvZO7xZscrjtDIBULtxanAcoxsKw8+zpVmY9wCmZMtEnBjmImXKR
YtwwZxmwL6O5ZvN5iejDXlJx1A6RBoq9a/g1uTFNEWoYmNjarPqRB/46jpSIqHpGd2o+yMg31s6O
4lE/Qw9Rwe9JbobOg65UJJJHG+KRcvgH91IEJUSs9Boa4GcJFcQMqqbCpJX+t9K7g08h34aeHqph
phLvqcOoyeo2tWGez/Y6SpnMJDu8pAZWjBLMRYvMcAcQmD2h//ayvJyb/v6K6q1vpL3tGfLvBuGY
5jYkamI4/pARUAkcZJOTUUSUWyw0O2cYDJ8P2IpG/7cgPFGpd+LC6UCRJnZcUIqCBpdzoChsh6pt
8t72BfH3/TKxDrLlCoEwX9hCZo4Tg9adBJqhv7BFBhw/8b9IEdOcA+ROxiRUBKqu69wn3R0h98A2
LQXx7QaHDmjPl3SUF6KOMmJnzunP4RG48nhT093GXUAQV/UR0KMzkGasAwNfq0skDMCzRpVuTHkT
HPgLAPIsgVSpl24vg9OJEwSC2b+hMeJPT0wA7sFwhMhFz24LfmHC2oPb1eb+tUg7HSWw2GZGa7no
dhIlGT6mTG9E1zV9j4g7YwOndspOv2szj2QrYyZrYMFJta+JhqvSKKQF0R+DRa+yj9PlzrgyJEhw
Oda1eO28kdngufdZ+DebqdsUJ6fIm3wMbYYFJbga2qlQXhBkz/vP0MhB/+AoKxB1CCzGK8kz0wIJ
6moE1Ej0s24cS0WzOx1lIfqOu23KULalYfwYc0/rJqvtSdcvassVY71M1JhATGo96xyAG2luqNeK
egOwdQ006wETtcknHT4m3MsNuvazzYMlF8U9u/niIniB1z8v9kjuCexRGwyVfn/OPu/veMnurlHx
OPeMfQfOJ6AJlliObQQIU/VyEuDmmHbTDiKG8i1sYeAPvlvGKTZ1Pyfg5fNkWUkY4w8v2EOkQxgr
aJ6kT2IC/lAXgGj5gv7n65MB+LiQoSvMoN8jNcahXIVyckv5H63DoNqP2cYoo+/SReqoKZbG8dfT
iCof89H00SJjNO0ZumyOnwO2Ed/ovWBFWXjV3do9NojHegejR+LhhkqGX03KMIgxTjUnMd7el3L1
3Jz9//dfyZvbGNNSsXGy9VPEWDj2Hx8ErnndVHicYhxKLdj6GfuPSMS3cmhT2stTQ+dWTPwUNP7K
6NxonKf5X+WjNhk40ccnU8Vd0lrwPc4yduqWUlyOwHumGK4OPYRphS5wgoqdZT5gidIKMqhvq/Va
3Pt8RJsWQCyEOjBC0al0fRYqFuECKia+HyY86GQf5x3nMOPlhtG5DSV/Dl3U+Iatg9bfNhh5oksh
9pQ+6+5M9wOmwnyxsJSBVFeS5zENixNGfL6H9QonkpXCIhJRqtuGJvTlzTjCkA1QjXrsEz/YjXfO
s+FzFcopju6e42ZWzASPkued6dvbXnNBJSxgoZaMtu0BWD9/aP3x4OxbF4eTG1uglYDXa9opKua1
3rTbkn9vpC/8ALFjool8vO5O+RGPalqv/bb/XCVyKkqFhMT922jM8LUck0p2StIQiGWXqgOpxqW6
npUyveGcWXxWJduStubjglmOWmoFUqDKEakQQICJ70r3znn/6qyrTN834mVc6QLyYi3UWXY/EE/S
AgfTC0o0J20iuiZ6rpBPUggqUOW6xH4Eh0M8s/Oe2TKb8S3HB8iK0054+WsTir+tvTyg3IOXi190
dnDWVmdFDJem1SusRCv/cbmtN79Pafeh2dl3E+0qfwO/6XzhwyUbx67E3R+3HXLgNZPNp4GcRQK5
yuAD9gW6mcDEdgXEWXJYdoLVEUkh/yHRMfJlPF9nRFMAt0PNMCNjPtLjSWjTbOtYX6Ip+YOt0nvD
3R+jevGq1u13M79hKsZDjimSOh04Noom4g465AVq2J1uBB9tD5i4B9TRVu45plqfHBCDzjZQnX/s
YJn0j7Uo3PjX16goSEBlTo9KHsWNG4Rwi61OGLmOJqIhD+VSzPsS24Ff/c0lqamAzVU2NTBGbtrC
/4A3RM7LaNXAZpv5VzcdIV0vFanBty1sBlWO0tzH4W0BpgplfaC/gSjA3dYSBqgioM79TDrVy5+k
3IMHgFZegKkIfvCKtDmv4kILaotRBOs0PDR57E2nkHoJrnaLjCNAqsEFCi5dDTk5DlZixPigV/OT
yLiOrh1K9EZ5Y5qOG+Qj2DcaIw2/2P62n1i82o8Tj1dWz5HE5VO3UxCmCpsnBV7BGEu8HJjP4RL0
ZJ9LQUG+5IdkefE46Bf9bT+frQmnb3V5Zs9RkuKRBsxAq5ZLOiQDL94ge/kqqIjquG0/sQsfRYJr
WsYjsnPdmu8IlsDIf49E9HAbh4yceyXRlzFv4VnZqtKltxnWWRJFRmwFeXhI4V4j7A6zjzXzODOh
OM6dIIq16Y7s9lSDGEkYE7p5yaGd6Q3IitVX4+yXtkowfpA6pIiGmFVELkpt9AcIKu7oIA0VEqPG
+kY5X9JYOsQ5ABf9d0I0wMglymizJEXR/6VMW5wTFfV2j4V7RrOJbnSR3tbQ/sNzxCDyqOPr0paC
cqiAg6jKw0vjVkwJzSu+di+Imev7GmlbXQTXdxjlZ5dfHyYrSZImHIIvFZLThXRAV5EgOKyqGiTN
gVEYJEQvrSGU6Fy7aKd5tg2NxwJJowm2awWp/mRjgjwYdtfCoxbFnGqZfxzE6ziNYImi5Yhlmy3t
+Qzda90SPuqhFDs81+EkREzlphPEyjfl/KfoPaE5aCyi8SYaFEux980scQV7DAvQdfeOwUu/aEwo
GQuBaGFuMcHup2iFyB6MxX+mdrgJel/CDiB7XO5wF7e1vhcUBqgun4fV7KfFqQQBsjbqtJrxm/3l
R3lLAlP9qgiXZPwQPPhXinSd14PUOCDAkytwNQfU0iQz1Wv+u+21oL5hnM+WXcym0TEvuv3jGLH+
EazbOznrV2+M46gKMu6YjSYtEnb5nw0NYksni4x/i9VL7PvZfaQw9VCfpcQXewa+odxFETUF6c9a
2Mq2yw81RZ2N3ZkPXBSvfr0EyJf2kB2C+fJfoOw2GCKfASFpBzBcbBAZmuHWSb+ZmYjHN8/sfRoO
GFU9u9gEYGYFdz4u3bqtdE46+EUhVJ7F+6nVXZItX4tykT1oBIolJnXC/fA0aV30nehyxRu/8Ayx
OCvDL+4F5J15qwlAkWd1AlCLq5zVpy2hF65YeHzjPczw0+U4DjC848uQ02yF70L7hfysvY3X6VAg
PDS4NHkHQMTmK6K2BzyyT/kYDhZz7QVq4QHBNfv8O45OXB0gShaDoVwT4X+poHFdfY9pNorIO/LZ
VTcpVe3+l8bsXS0vkMVGUiwxtc0ELxGMXbPvrTaR9DxkoXEH3g6LTDfibDsEJb77FSS7hwN1/pw8
+NGQx4pzavtBDLVsvR1sDY+9LWM4UBEs7DTrxhljopqv+EtGVFtZnrgzZkaSDRV7SJslcWWwLTiS
dhGdJkgDNp6IdH7/GfGhdwhZDmnndOALM5sUmXJ+zugW708GN7NxQvc3MUOaFwU/9q23dHzFze1a
OxomidgmF1AFbw2DTc2MuHQJv4qjd0B9S4aN/08ri3eKyJiVw8387GbHHqkcOUXezAMz990C8bOY
KDTjNC1ARnLoFF/Z719uLeg486hJVHJyh2+o1X1r5p+OYVHssy2GJ4AxOAgI4kBkkhSr+UT09KiY
Kmlz7TYJRiQtUHlT9Lbi6+Adoh9YuXCgmAEg5LjXKESbuapYcPNEHCtfA6YFCFyp/VU3/EXmMDF5
VuiINJxFiR6O7MmdlIiv0OTZfVIdLKg7Pzo8m+G/3I5BbpzJM2nZ4KFNGUd+SOxSpsV5/HPD7lGY
ur5DyTX3X6SnMSvKx2mH2dsZ8ZRa8nUX0CwEENw25YwUGYVu1QxF91wGOZPEiK+UPWhh6N481s7q
GC2GRd/fZQz2YVFC3RXUKs9yXVIntRudse3eFaZFzcYtxMVXGQl9W58Lowt8pSK+W0C8rvBuV9dL
vDlOw83Pt0F9F4BohUssqzDagsnpVcxEJfIXIGs1kACdSeCPebzdZWZ5uam7+gAcXuN5Clw6H7sB
Q8X6+YzBSOVkCarWYMkmVDoW6g47NrEo8MUwVL1pgPV2YTtRI6+4vLYP5qWDykUGWbq5N6H5l5G+
vO4s8H7GS9/huRSpUgJWNcy3aBAUCQLNywUKH8q0XPVTWgzfr18LNJhs2f4dsuhPVJaqusVBZCEq
RXr3LDlLPdAxSB9EqNw0lR/BYdI9O56x2IeHCyl1yR7EeCKYaTrCqLavkkFrg8F/U/KDpfuVo+13
a2XMkGCDH8So3s8vOLgEX1HqxHMG4RGNKtCmprz+gYuQ0Z26Ui2DJoSd3RuXjuGMQbfs93DaWJbZ
hH4QejnrS8xhPCrv1iuXg3acbIxxLudrTadEjx5T5dk4Go87mIl9gNUc1bPn0UEFsvrIivhFkvWQ
IDe57v7spg2/HXGLGzIm7qRVZGY9DGbv6BfJJTODQ9UjPRpkd4s7+WNte+6h6wO+HrqjCm5mTV1X
w/8kPQnMt3DCiFs0mEvnAgUzy2GwZb1smpLuiIyrOAINt86lL9Ai5wci8vR0V01azgQRNZaH9M9p
9cFa1UauxrrnMbRsjPofBphqGBnK3Bc95JaOFyOOuzF15dPi4b3NifER6kGxXCKCjwh5EbXvIMSR
uHqQtXjccAp0OphnykBJp4SahnSeoKinsB67/RxvUbPGHliILriH1H5mir7IzDqrs9+LeHELl90w
vzO4AVggT6KiB8sUG/9ia7TuBpZ+WONeH48/zVekSTzYcUS8ANp0FfugW8qThu69WUxtJhYkA41V
qrv+yL+8jWdXVe05Iz7rFRamFgnrSnCSO2CmChN4FnuoyLjZEuU4/6jq2ZtLekkQKq0qDhxjm7hJ
p31EunYx116bE/Rst6sY3xxtB6uqjqiSRGgmTRY1uoBCEggPUKajLCrT0fJRCbVBPttjfh/bZhKc
kLqLgqmknUqHLlu6n7fGYtTrgVuZkPFs6YAbTrNhBliJ1EN4VARtb+TBbPjxYK4KzEWeJDbvtJGH
OjLeYT0p1c9roulBDKqEE2GAzdUsRKX0cBh2A5gE/q6KmT+IkTjUPqjucc1i5XL8+1dfqFntq2Up
cVNPo9maR+Xiy4GzqqcQIKIfkDsoL4mSpYQI/Qb4+/kOqVJWhaVtNZX2Mm858AFtLdEIa3R0s8xT
+CGbMUW351oTqPiASq85bO5+ZtAx4q6q8ApOCEV4pC4kMQIMzyLwV5hyLPrAHYm2CR6pxXOcmlvf
hD3TO0UL9I/CLeeEyGmwR/gKKdph4qJqbqHRvqE3wLBcZMMqn6tW+sRJpEtCa/rBB/RYDxJrlhx8
02vrQuG8mtJPjF6xkLSAD6mCeJs1KwsaelgOHH3kJOEWpcOn++p0dtH8lHRYwv90LmUenB7e+Voa
S2waw6DoFysjd73yTkTA3z0BHP/L8emWKhUZUCIne3LdkZt43IAJuRLZNKXeL90fviskMC6n3ZSl
N7apBjnMhSqigb1OO9Ued48mjxcdJHVEkOJ8f9BPnkLD8Go0UkxTZvwBP/ctZ8JA9NRK9DnZsWzy
v6s2gDJLWoiaFWh/YUQKRsrQidqvwnR9sxAprBasMNGHBqOZ/KwzEijUleCarsmIMeKWBUaS0fMf
x/9EAxxWhJ3vq7iwN0GeebFcw7FzRH8Pdyp24zTL7RHM8PU/Hpb3vjQP00kwcla2A1kfNd/jiJkS
+iFN3DGYLrATfu44I2tL2OhwdvAzO6ANZJd9iMr5isylpjWkVnnryIAhfQzFG62uHwOO+XDSgzBl
EUfUQCPeTQVx/dU01YxGwK8yy/qvmxpB+rsX9qZVYQta1hp4m8dEujfgn6nxA6TOMGBs708MWGQ4
LFnL/EgmbmDVBkZv2lHAANH7J1YwNg2lAxBz6Kg4O3qi1kQbKiQoxWrDN/w/N8qqtd2naKx/oqyN
RblW4TidxrV3li6hjz25yigEyU+uZcjq9YsSW1L8o4nEaBKnDeaRdOAPxdUck0viBvr81s315iWR
RBNATflsYYKhij2WH+9BJA+50cgu/7YLsoyzC1dYFR9DKWOKutFspJRC7lTnOcU+lslL4f8SxWMs
xVc/nKZh93AwVk7HM7RiS1ZLTC4T7oU19CJuDtIb9SIRBYL8vlcS3LaISIkJe/eGc+QA1BmSy7n5
tUft93LX5rRUOFumChONidJnaUr7lnoRqSHNqDuMHbg4spfeIgN2EFKm2xrVIcEJ3TZ+FC80PcJ3
sErG9oK7Gig9zOVQeDpvJbKrherTdaHlfIHfH2pZjUvQiqwhn+ZNGbPzP4RY5T/csbJHOpHrsQq8
2WETmYYFDV5p+c7aCmgF++8O5GeDwxwybUcq4LgR3OIowfBaLSkoAH1fhjqzisACa49DvDYRix3x
bMHGSjgr3/tc3O14B0FDpSpe2jxRssGcOqv9Jv85urBWs5tiXSDqvdgpefM5RXsHzUrusfWanqI0
uqcqnJc01zv03FQKR3Z5Uo4l8szL6QlXlzTztJAZFZ0BkfSYW9eGYyDmZ6gOaafBJ4edNd4BhJQL
vnesGXhpQptdqHlq6449DlKDEkw0psBFZ/Y48CreJqeIVnN3FyJeWL3QkNHp2meGxOhcnaqJDQ0m
Iw4zBzoKukMIrmULdd4ze0ACSTTld2u2CEUQJogRtnUYOTnBaZLxqzvUrB9/DiGcaibuDRMb2Uaw
Mb+vR//gJGARzRphp98hHgJ8DAd3QFqPs42GEggEjmoStyz7tsZbbBlNzYs2GGh0zdA1FL9vfw08
Q22ZVcRDzVlHpPVwQJRiTV7SnqkVWbFMop5yuJoVKIMD7Ms/sV+g7nkwupy3qNlU4DgusADWzXWe
5KGW/9atkONE6aW5kHlnEmXJQnYhIHJ5NwlAs2j6ofXQmKnnSLSVdnoCkuyXrQEEr4IQLf5HRUB8
De13GjOQk8u2qcNCwOiG6ALk1cKV2YChVD6o8UT+YAiEk9OKwrPrpt8Z1Wyhit3drqB6pmyuLmdh
uDju9WVavMC73sO7Dd4lFHqEuNO0gOB/gNyg3r29+cD7bm8jiwDALp6ZF4jPltSTxhB6z6AKx0Sr
+F9nWbIN6FMAltK044GKA6MqNEHH1N+rxr4MbMfmD5MEvpAb4uwQqgw5dnw3WVojXHOoobRUekAH
Nkc8DUSETsaKMBFMoxEhEraKzd1XbW+f/qtxw+f71M3jkoHpldQY15JsVEQuQftgEpWiUKn5yHgu
9PkXJdAtMypDVywEVAamF7whe/eC1iE6sHqbBjOJNz6qsy0th6jpSaNUvlW3oDb7lhr2/HD43g97
xoGm3IfVRdoe83CvKQd0IpdLjWqljV5XZJ1qDMq9hAoSVznvLYY28Zy3LnUtgTDUR4s02y+Eff5z
D544MohrAbH45/laKobd6GlqslEhia2n7W0SUDD+HNZ851uu04KhqMCTCPSV3DZtaFraKGfpxpK4
Q88ewhIspgrafuJovLRV0fI8cPf5D4zEjeaSqDCibqiF7XrlKFfXEJ16lnRbfVnzqw+ckBPfTdhf
PnE/LAhNCUj7yFQNn1Z3dX4Ifn2Rz+zEjJzuUb6pdJ1lX44edaeWu1uN6JKJWvM8bgLy0+/BxXHS
oHPHqh9agD3DKZHSk3wkvWrBifIflE6seSbxFveKTKspfYRztb9GSKZvnDBNZgG2qdYvv8nZWOta
r+qW6CNNDY9AO1Tqd4DLhrtVbAt9fduq+aOe1nfJxoRFT7rQnetPxyNRJx0dREm3fVxcPfF8I84Q
HyB7i35mmuX+JMM02orff1nmIPlYhqx0VZhw1uuk12IiORfBCnnA+sozTtQXq76LcRaCgAZmX8mo
fQcoBeByveDXLbaFiPwgOTZfb5XQTAf1ADbidiWxy0Sp8ytJKaem4vHLWRAj3VDZwRD/hnGYlpav
inCLGv5vJpvzrYrfnwq9Kqs6dDme4fhDN/jeA5/4nioSZBuCjz1LbW+UdqA+avF2bV9OepytoS1c
LzsSP9WBOCWIEmfHlUOEE6A8Db0ZL1trT0+HdiceQUdkAikPDdiJDgBzU755taWN2s0YqM9/pMWs
8Dzo0eTNHPkhR0fo5r9gWrtoVazrpsKHQhe13vAqvpQqAEyTmuSpv3cgW79gBBhFt3R8GHy2wGpN
hSsn3l6srxbK+bLRB3p4IM/QuGCWZkyWHE/ybi7yiwp2q5l/d5y1YZerZKW9EbUD2vqFVhp+fj/i
gm2D2FoEERinoif/nnOyCc303HP9KIeUppWC8iRD4ldQcZGVZgraPzWGDXTIN+XhHU4HaovLKcwp
urrAD1+LKE6OBLzDF4GmqegolkX7g4ygGWfJdqDxpUrSeOf8gZmlLOrmrK2ltWBYWAIJ/4Bo/WqA
zaSeIY2oS5EUf/h21f7gnILRAmEMPlEFy/y7R9vNFJ8ALcN/VFExYYRaqWwa9yeupZtXQ9gpTFBP
NTGuaRTzcDlQEZCizPYQL/4AWsdg5/6rjVNp0ytbr2YdP455b/h8A+umVZTscYgLLhwXBw8BgBKT
KvahBPSX3DvwPuiWEIaYr6dY/wL6zr+qLx7JOaHF277c9XP7eTbYT8z8Yd5oNDYuf5IQ8akLdmQ4
M4AbnG1q5HHb+2b65qxE/pf2Mhh9M1g1bVjKyl5xfo6fSAsP/WLOU4rBuz9pbjzRLb7Y9ENCfqW1
Qwvjq+ATUIsWuFVPXzjjaraKW2TGMaS7+Scc9K+vxGFjLNJr2rwnggy2NkjiwIRUcCsuqFV+Galb
LtTzyAv1VP4NYKDhlWuFizIDNveql5QEGJhhWhXOVLswhc/hmcRpCfvsmYC9DzmCS2qo3OF1VCEF
hJtBtQFFieLX8gjlHxkC0sp6Yl9uVxCfL7ES5d0CgRbKugQvkTxXCe2rSYjw15wPGq7itsuDUZrr
i6ApXh0PG0JiFbMDZQhfd17OLsCrkl5CId0M1SvPaH10wgoildXTSTKgjQQqk/K59uouh772V0am
/Hrsh9AAGXcmdTsINya0TnQSzABNnnFk6C4RDIZjVm5nLBWRSZOB8IuAQGI44qFfmmNFhik47306
k9BCr+T+V4pH6w0NTBszDnNtK09QE+YLPxnrhi/y8vSz9awH8oGzKvt13YlNxXVBCAo2sTEyDKl6
euHj2GKp32aINgVnbZoj4b4iLo3EVrKt481cyiAR4fwkaj29A+coMvD33KbmqRgjAvMGGvBj5fAt
mOjMNyCu7m8INNsUccEeD6+pU08C63morV0IXvAkv92erF2aEPbhSLPPyvUOfFGkvTMZU/LlcAQj
LHIKTnSL818B1LGlVk5pxkuUATOwlp0uAvad1VqdoVYLa84kk/vHarbk+C6sOpYkhTpVFAyq9MIB
B18kwFz1W4OTfcxdUirJstXjbJTjCjlQPBsSsaW20jdA/2TM/VRNd7YhRVR6VwruOzNH3UTr7si3
7rogPjQZzrxVxVxRQXrgJ0Shavox8eFf1B1iAArexmE2WqEP0NeYwfeN8mVuiW0mTRlh23HtDQzH
/vhrq9aMtertX8tbyWRnohbGG5dwVKuWaUUDAUhS3NLIK/Ic9mVfEFQMnWxItdgc0voDJZ+nFusc
5jYdghxxCmmbYT73Yg+IaW7W5Vc50d/ZrVuZG8zVUp8cHkVy7y5MunFzfH9KMI8mEeekA32d8k6/
cZ0OciPpNRj8Uv4wHeeF6trPPNWSL+WNKcqT3zNZ7qpqXIDrSzJGDMVOJCKlC1hOhtE9QHJTJP4Y
lOFhUYkgqm/lAqXPqPAiKQRXecpN3UAUUXjcfln879Qem5MKgJjQaAZm4rVXrjLPDcqCeA12FMpn
PV0xklsKeZ/L6ZdRkhM7A3orEyjHGq/zfDJD92TZCTYLdPP+5cV7DQ7aAXrjDl7GdQzkiY/nGZ2O
kp9EscUGEHpsjv/E0qaQd9kOmpoKBJ43d1MJGJlzqv5uEsNBWftSNPrRnR/qZGBupzzBxmbAHM5+
XyEIon/+CFsGQrXiBcPbENV1GBykZD8/sbEnfuhdLtSeTcKfLFppVoUW5DbSm0epXcnn1BDGgo+X
X1jvQSHiZpKvQPy8wlAutxRkOZG9UNqltOy5q4RMD2CfM7AUZGGRiKXFLKrKwvAcHQSFx5CmDu44
DAT1nMc+6ykANtjVy+vy6VoR1g5TQwSrUpFniorifxCGKzH3orMilCOxsaPSGezKuyT+d7Llb3pL
WPw7a3fpxhN2kZa2wBEq2EAB15cJIGC3nkF/6oMggCgHxZOl6Jz2a3dtcAg7JsOxqLoTMeAqZM3a
Hk+S4Uvu959mByK85FoQ5PBxhj9VYMhE9QjespvQL/mSPVAX1ixbYbDuqfLz6fSs2OutMyEfIKtO
AHjcE/5A7J1oR6IQxWWRTq6yreL3IPJ3Ef0khYrBUz/00zJG8SG+Sbm+o4JgPra7KMlyQSemWpq4
72QCLkbFV2jDyNNEkNFfN56n1yJWfToL9vj8aAuU1HuNHJhnh8/iuxQ1ZXYFepB5478EFBMS+euY
alQVGAVbnHpRuBtK7T8HLI5/U+6G3gWWLa8+xi1U2AjWZ1XjCjaaPyrg2NQRWaXIoGl7MKjwipk/
4TM1gcZvkiEE3wqCFjXctmnYWXU1p8Y4fUMiqIXlOl0HNTcp6KU9tZBNJ1ZsasdUI4E4OC8TeDYt
WMALA+yRVBj/dNDFE6qmRGkSb6ZTpMLkCVCA4MITNlGWUTx3J4n4C1H8mgzdTF/7Qxt2tX6bhw+Q
FFJzdemvjwyTKSQ7nv/nROHVuk+Df9D5T4KaXu5TOEdSJJhc55GhezERn0X2UT6W7s+gU+Z5TeBA
q8AzEOSxd44Ir3jS5GjGYow+VW39D6Ngk//0+72Jrk7ShRYmt1lhep5rEdWteZEmuPC+G7mS771j
tRQb3mEtPDGQSBq9Y7fYQi+OxiulwGN0wPP57bvQfEo/d6lG9J671DGCmJONDHPusnqpnFrkAx0g
MnQ5LK+Z2d+WC+hfdye5/Xz0oHp8/x9x1wBwEAEOwyKVSNO7/T4N2PByQ210DFAsE590jKKKULEI
xa105QbGsdWngXPaOc2GGYfJZh5gyS5QxSKg6NtzYOZgjYnmdnMmaE6ksqcPG8kL6BCo0qRwSpgu
BPhXtI+f9GXJYd3uIYA5W9Sr1qyI34/MzQ1m2cuSBQOGfMvz4qgqzZGmbxuwKsTgWuO9ZzJhlepu
MBF7gUNrRw+R5lpytL++vV3M3EoSHIev/MeX5TeUxwWQdovrC2uNv1UaZah6rycmtKuzqE3VulPY
F1U8f5GsOtXl64T5UEu24OPonb7Tl1/Q6VlcO8/yvfmjJe/iIrbMnz0VH04DT/z0fiF2aRUJoit7
0VgKUNQRC/7XeowKrCSE+0srQUAzNnfqrzqpaF+q6R5JUJmWfW29Zmblpp+FjwEASUXzXzcUd1X4
Fn9ymU2qwlHjI1/Yma9wRGqXLnFedzJpHZL0NWoFbREDLXNUIQ0qOuRNG27hOtvg6jf2A/jVypon
ZYVcs4woDzu6qSzdpykzllqwc62zYOSIUTdIGpqXfOH5n6WW8ejqdhSrjYxrT7g+3l002nevPjiy
B9KfT5qd4ulNXOWMr6XipES1+yU1S+XxKV3+kuGqJ0jB7PAvluDpp1Y6okkL6JAUo0vDYIgLd/Em
qv8exGG+SXc5xmS88L3BXyJuvZVRpiap0kX7j2tJD2cYnIeysj5V+RoQZVnr1fjU2T6+hXJcdiCC
mIpXcAzmlS08JzaWw6TO/9YSCjrOPfluwAty9DZu+h0BSkBY/RmYOYPN2L+rDKFUzFLJIZHDuC/V
E4rtaBKflF/R+6vI/qn0wDKPLCXGufqfdkqEvH7I8X7ZjvrhFnJD0tWX8WimXTAoBJdKXvU88tUH
NUZA9MJMt7zmJY+GaRtiT3NYYYVQuWT1c5N5f8w4KqtGB/IZzfx4D2Bu1JOtF/yODssq2sKbXnJm
yEuxq1XNFg0T3NVhHDAQl/ue9T7SmSWyVvCaOkXTo/3tStJWKCc881/XBfqwn2OXz/9rKhm4vsz6
KHEdiEarkYlNHKqnv6dlCg3T43l2FKCkiNd75c2J9UTfhia3A1CIqbW+IatiKplyTMcOkRJ/zpr1
GhTwUQjkZwemnJcoBxqx2dM1c6OFITWV8xwsLZ8ALjmC1EQjiTqHaXs99IDkrL7F/tQPR/G8qkSM
/5aMu+WSQevmcTGqiqkBO5jJDb39hYp/B0mHWR3LelrDh1nmdhTRZcro6VhoPPB0MFuHzadXmYks
OGXP+F63NplY0bahgIqYicIo9xId5OGBtN88VbGk0Sq/rQMVGpqA+nNQj5E42GmJMyBIRlzuKUPE
3wOtehFQEe0Ya8sZkwGIcC3uQ+nzBZvwLV3aJekmG8YtWRBxCurcXw+H+tvgCW0tQK2fPK84nyFh
XRo1gHyriqOQmXA7tYVzkilC5gujqLal41XrT1gCKXq2jC2rSmfWHXO9/qRmOSbDLQgVQ9/VXgZf
U1zmzMHyHiPbsvv4889+zpfhxDSbqDh4xqDbWEU8R9xIOdWZAsDgdMeOGGmWQ8VxG6cL8bMso0EE
kuMgLFMGn3IegsqVzkEwJ5TpoaaE8Ug080eHS4kzvuEnLxGnq6tvU3S/1EFEm0p2eeE11D1wYXiz
I23+NsaIhAU0f8nInWi3NwIB+LaDywx0Sl+qsNjsqSDeYi9JHJogkBkC/xC9t75lXkdKNeDqReBa
6G9JCWPyjpbcY+YE/Mrkege2Wf8PLt8J+mP2aRp/6m3SoKzExESuiDULzRgfbNya8iY1gA9aJCUx
RsKxc8Efs8op31e/d8729NaQ5xaXo9q4B8Kw06O5XfBxorud7oumNAodx3KOL7eGeMvJZAaov06o
BHtD/ql0ZRGk4vDeWrS1b1AcnnCA4BUWt7ErYdFP6R/rEURs+ViQNexM/w1ZAmZ7Tc/ZUYaBeS2F
5b3395EnE+aJXt+tPBp/8XQ3Gom0yhYtzCXMG1TL9AjbUFASMWwAcAYqh3GRcL7BdFpzCVUDRoIw
SAxjAHftTFdD2WzOar6rfDI16egI6C/7jvlyhfASnQKK+hf+XeatbqQQxymxVyqpTMAhEi8aBDU8
ozBKG2Dnz9rqRtybNPejIFEqmKvqzoBU0oLfZPKGr8NWjj/EKhjvr6MI+P1v6qFzHH9dU4fEFAzp
Wh8JGGMo0NlKx94yiBjSsKUsFEq80rDbv0OgocxzlI4LglXunWXKNCYrhy90Fath4LOMBs7Z+a87
6krn1bLZ1qL7jRHJHkS9lSaLp5h8D4Z/G+LfV2tuoVBHZsHOQzeYYniWIc4BJ8aKZ8EJzNT6TZT8
Sjt1FGYjW+jZ6HdUTsianb6KcIJMNkBv7qYbtFSguJ22+JNO9q6kFer8TJ0rRiGg506sU6bjeYik
X4pIWplGFl+I+igi8np6z/Olx+eBTyssnfGwx+Kd5L/piolKElhTPpjFgGZSkQuRLFYb2xQax1Pi
5n8jvxQWycBpFnktjj1HKj0nWr3cZ+r6/nUeO4QeMY5+oDOz3MewndOiwiQ6B5mcjoGD6RMV+HRf
mkSTklZWpIYtO+1brFxBeH0F+AlBtMYCnvCvGneStk2JNkrSHQ6R2fZ4M/6mnebWOVjsFpGHIi6B
+eVPkSkvlOQ0VH6oyQsl59/SyYxtl+ntOs7rkZzQZFiv76CP1y0EtByYZRbADBLyBcstmteKBPrC
fvDaytI74hLRmF/KNVgDI8/phhtCelQRWj8Ks2gzoFNIYviC6fM55PZazqBpQZ0qcgg43vTvFRYT
x5/ZAebb78TXthol7M730Ol78nCy1bp38FkG3eDZeNqpCyw8B/zRt9lLZzsAp8D35DsVLGn4Oq3E
Uir1EPNIW9nJqDy+gpp6gO0ElEPgTRGUA0tShkvFqOEWDYFfsyH7NItf6ZAJaRqiXOdoU3zRNlWl
TSoZZe0r3O48UGcSdfyTf4sUZYs+f1b/zQTccSpX7dt9g/jPT2UPhcefRGfEX62x+R/qp493pyjc
9HNttV5r4K/zzebkLeY4SRrJyBpA2VjuhkBJ1WbvCDIlJslWyH+btf9J+Z9MZXHCKBjr/t+BdYo+
j6viaSRL0XH3vx14TcXEcCt8Ij/7n0RqBHBb5rneXl23K+/V54lbZDAPeDoTNjFJCXLVJm7eYa3K
4sJA0Hh1A0YMyvQS2spGYz+mUHiLIdNi07CLrtbnesf/xzWho6kTOKp0wJweMY5pCoQbKUBPEFGN
TfQ8hJNCPIpblSFHGIOhks02F+77vU8ZrTSlLgePI8bGWF2+HMJkhgCj9+VzNUywMR1AnwmTZ6Dq
YXsyFTjK9ZmuYFuUjnvB3rsALr5FiVD1IHSGhVzY/0aLh7DGPZomlur/psu3cDGAAtg6IALu65JU
Rz2KtF3gGEFgLbEKMjLxZVKwcdid2wHTjqyUh20dSoZYXoHAUoqjjqCcI7/ydwxV8zHtXrImnGyd
88ra4B0+5X2VSWXQNCperRZpBwfp+vbttXrJatO7sVVd6pAaoYu7aTcdJ81PvuTs0k+UTiQ9eRJ7
kmcrw4m4cgG6v4vWRiiUtEoGhiAm3bfMvofYwUiLS31Lft1oqh+DdHHoq6Zn5ER8hV+UpBNrSrDG
1F+XAVh8/KnIPcbEWMR8oBWcJu+45pGNSNtluqiz4O7sJ5dkVh1xW2kKRKJ5oCjEVGI6o0RocqDX
dQAUGwCJcfLkp6A32Cu0Um5OjhbtytW/oZkALCnewUGJtOyWEo1AhE5qjzu1DH3iRxgrxAutb/PQ
G+AANpG5M0Il+c0Cmv9k2QOe4n9oJbeQDdEb+7H66jk8VcRTNGlJ5zQn4SvpOlxmqc8Um3tpwPO+
V/1hoAiErx8MQ7X74oFAMjj/y5rs7WIQ/dSRQu77dPHVMtl7DgdadM5hrOS2l4gGQKyvFyuC4Emj
9dyHeTG2Z846kAvS2EZmrwykc/47BQoljkRcODcI1dI/oe1iRr062BTbUzXDF0wTP3sFLM2IEI48
moQpIFciY6dYNBr4igICrH8ozC7NuVdfxWkxyEAn43Cq2WTawa0/OZ5jJdDAQZrTLF4vKBGfnJdN
oMtyT9IWWdfuIPLB+/JAj1g5e7JLQG07vSJfyDiwlcvKL9+bgpeSZMHtT5vTw4YzOq6yBw3g8KQH
/mtuZ8WgQ4t0rHZgaYotYlZ40k4vkuC7NyFXWzOW9RRckhDWEQXAOIJwpX5nMth3EH4JH+QgPDhH
6Xi0uSmo11AcYmqI/2H33Y5UniPtAzMjMdGYUGeKyc+Tt10NxsyXWe6p+7LDUsk4iAjCkGJKMHF8
0+vVUJmT++mHA2WKn1WtRTkk2GD0YZdw3OA2DB5onh2Hgyx/vB/vstU5n5eWR659wbCEdGtdC8Pa
9CPdxn5BBWuA2+1F5qjZjbYMocuiRUv+7NWmcFQzwfE1V1bnJQDyLm5mH+0o6FLU2RGJwdl4ZRHG
21AF7ZZIbiC8cXRap9tDUJJA+hNqJdWZdjN85eB065Il5UXdpbEvFCpjeIH+V76FdKoQP7k00phu
HYUSwh3iC+cKyTHrDg58Lk7JeRTsiQOU3fA297nccy4g+APAQ0I2frXw2jt9KYsZEl1nhy313dFt
Z4FYFQsIM6byLSBuK6QtlKQ4vrsiNv8hD2GFyTSCvpD1qO+kswPuRy+/+SiAIs86Obdlwwn+VF1k
fLkaLlPySVkrNF0j9cF4Hjb17O2QVNi4Itvg4HRymJ+RFXX2AzZazvP+aPRjzog8O2r79ixoyH7n
cGuLv5IgOpxYSzB3VucZK/iyilS8OyPgK7b3V1KIQaf2285uQc4QzfhAkvc9eh/ZYplN56xssdiw
1Nj5VSvJ8box6coOKEl5Jr83PJn7N+2istPm/0rP+DaQ0s2SipF3GXOPTlp4Lu7t29CABMnbAGxH
TCWYTnfT1ESif5IHrIRQYFsHlmmpTj07k0bHD3qmYw8zh8FNhyC1029SZNdOr4iu6R5Q8ObSPoN7
WqNc+CGIWeWE4KotTmzohEvKoeV3G7+7wtStKt/cfcEB7Dz0JgVUOa8lGmZ5utHW72dJZbbDlg9W
DEe9zjKOZXO2BKUd8mQJPrVSJA0x2Dlmub8F77DQXnlUHgRrKye+QuBTMM8+XJ2rLFVtSAETqDeV
2yRLY/aA7SVYhfvpmKTgz0mMeoKvEr3tuFMXzZpwC4uDtSKnLVmaFgBUsYCdFx3a6cyuFCVGVEUK
qjGpNN/2l1YBaMRkXpx2jWfuF79r5PIJ761QNcDn0JO1cHH7zVw4v2ADV3JTBQzDABldpYLnwqCr
Ng/OP0Be6AE45l51807mL5HBXQ/gNQuavd1ibUDEXl/VXZv//t6dNewKfk5TSBTwgjUxHkdos78Z
7Ya7+srfmHwSEfOeW0H0u8CYlZejnrbwB7zbZxlCPW0IpiC2sIfC9pnyH7T6/Y9DjycXxPEE9Nm3
D+SKiDRJFKUBGUf8ddFP5qcr2PuvnSXf7L8j8n+wRj9xvnZB4+cAkGxTAYwQj9TFO+Kxd6mvuGhd
Nnyzr16IQfaCr8EHVTi1S5Nku1pflRWm/YuLQypFSW6yXKpiB4Mt0zbNsdWccJUgp9UbTUL5UlXg
abt5k/2u7DAVGzVsFSp4wJqIfXPORK74FNkNBDXXlQ2cWfUn/SjY/A294lsg31vwR6n6Lij/SL7G
GoNZCcs4BqfeAkD/7OFEjoAAFdmYuucDuZvnHRwO9NM3e7rOXpBPnRvqu+ks5mZGWRK30EqYtJvC
QphZdwg0i0QV2EUq+DaMt2AkPG97383/kbVKOeTGV99ZWHtj3XSAfHsPHDeHhn8RIru3D8UXe5wP
P9cmHWlz9wDm+K39bYWVG63m82x4wfeiDu86mK455J4PkVi0YcR06RdQ1y/q0Oh6x/eGaTd6G1qR
o+7UbfZWHZu3Fza6FtCw6kX/s2WLTzpjtLTkyv7km6enXa0LEo47W2TcuM6UwlH274X6KQpHXSbP
xv9lMQ6pw/BE8RI6T98gszJ0qxGgj7JgV0JMMAds5p/YdVyvpKjVdPl0mw71ftmM2lo86iDSOhix
iTqRFJS2YYiQLljh+VA4DW2J2TjwtdURTGgwel5YQ65R26Km8ifSi4A5sJ1gf0L/Gcv2TeK9gJ2d
VG1F8vpjL266lD+LVnPaGNu85QjHtDf9NeWTI+ddROz7vKuQfiCywoM0zZKALRvC4bgkyN9/JUe5
nXs5717hQ5cJG2VDmvFZ4Q2ANeiQM6jxp6YAv6M2VM9V1Wxy+d2d3rE7o5TwxRQmLaklbyhs67bD
uAN88Qs8uwqvQOVkoIyRcTIbaASung+IhCRHt83CR0rjvGgoywWwtrd5kcI6t0vArsgrDr8iV44e
bYHNNlKV9wZowc2alU8B0kOg6DDh8aNhqI4Nt/RHkz/oKphFl52qrQAqsTa0MA2wn4/rbxnfLysC
rtH8fUp/GwnHgiJ7HeZ26JtXWgOdypY2Z32Y3hzuopr2gTKhHloyVxztCwZ1Rbh31ejQ6iTY1kg1
rvd2/jnqW5LDDF0tMelg7f0HfngdOmjxtHS/54FY0n9zl8QSszG+PnHe8Tkf0lIG09IJbjWEhmRV
xusqDeQBgj7soF3NlMRZG8CgCA4AKnrr9QEz5DYAbubQQPPiawbvVibsie9EEwTSvhwBGr/WsovN
gfpK/WCY2sX/TIqbmiyEsDlstWgIyH2egpmXD2xsQx6hpbnTvPXEgLmB66cIM9fV3thZ1AGOqNzq
iheXDsH7ie1zQf7DYrUcUdgmwAVvshWbMOx2BjM75eaa9TQhUZ33C78afZuGDuqfSrP9128S6WjS
VwGRG+rlzaLaWEMlmXDMqXneUygxcdyl0zHisF+oy8x1qdA54CewZLzAxWrMEesFAz+EtDP54qvA
pyACUh2UDaEUMQ/K5w0URKXOub/8I7ZoQCdXlbDURMqnYKHivouUIUrkFBALgsr2YnYa/VmA8/sg
FKGO9uxdyf4l44nDt41dMiNIlSNr8c77UN9/QfiMqP0jy35UQOBVgayakgKK216td6LLBHa7HXry
9tK4XnMGeElPu8tT8HCHN1s6udmDb4NjEz4MIx4UaD69NU4Yw8BnpGjaOUbMm+kNLXtFlo3B6nva
p8uPBemmVL2AYTmDRwbiJqQjj1ZZ02UJcm07wEcl4fdBv8mk+u5sb5XRuhkrjGmvCLIe+MsI3u1x
J7e1M5Bg3AOovDyFnzy3GJ16TqjpvCg4TegwClOKm39czwrD8cffd63lKF+Be/b2CC8Vkd6aaS89
Ahs/HPWcPlbvS11T9e7+RBsuuLrFQeWNzSfIe45CvXnOCvi8w/oX9M3LrvfPxY7zoq8ERrAhEN3n
Aa+mZ55Ig94A8nzjslmW78jsutnjjKJ6dTpINqVi1K8txeO3JqCcEtqjZLt+xUjaUry+Tg/8Hdtj
WmOROsdxfHs7JjiXXAwbLHgF0optBuSpRJ/FeoWPKi1KEWHwQTRaN3vCTdTme4uRy5vv1FVqx0PP
Ojzfq3QkkRHFQIDEfnxLVJAaAtesDoISdo2rBRHU1LeTjRCw10Wpr+Slof0w2QmP/6wLP47swKbQ
sAqhBmUl80OHolRi4sLYRjMXfgsus+q29jedPEJLRh31Z9ITbVLj3r0mNm0AgLF3XUZ3ZFY5jW5a
ZOzjdHv3FcCLy4GKiV1X0NJe5imsYRdWko7oQktYTxd2zwGrEBqyMm/7epBmhW7T+9er9zqzCSgm
k3mkHGALePjAhgras+Kvg15RMGbHuALQ0AIumNd2KZjUAQXDzqn135ULfzB/zxXRlGradwFm8Ao1
K3f72K2FD5G2WksnSjPQfM3t+5n+524bjaMHWQ6IiXGH5VgxdQ6ilU8jO83/R6MOKq2a4M1c3uuR
olY8CMw3nZWN/c23g5A5V3lOSN3mGrPfE+trmKu8LgKlznmBbIYiuFeZRKakV9VZ/qGSjn2QqULR
7VHmpV7a2Pjz2Qytsq0iHfuezx7BSOuF72iZqKs+F1AnDbTD8OrzCkJ27WIiIR1zq7bv8H17POw7
aMYBWdR2xUOH6ICulh4lh9X3z6Zv9aAdQQutPbxJPc0omnmdYGJXl0/IOCXSK+DJsPMY0YawCsip
rgwYMhbmU2qZ2gQqPEQBPTAeZnPDJYteBAzVgeYigqyVJY2JCr8JQ856DprM4pu4y8k5/yLB4VJu
/Wo7C4J3LaqbtFNSCtAZY3902BBZC0XSaf3XAN5DuMcHSisVW82AoP8igju9l743Ht8G3qCfA9yR
kM9gy2sf/wMpA6IRVPV6X13RpdlBbMHMWKATgrloQv+rFlaKS7WLoGIQAzU1Sw6+tentPx1jlXhg
TAxeIqldQrNDlZH0p6PkkgltE/tiuL5OTdaK6erNq2M3RS11Ha/oQbnE5fCWgsMUwAyt34y16ZqF
dIQlhR4c0e4B0FdbTLFkwiM/J8z2a8DqHbC4XqAft8APblikGdwY0b5PU+eCBC5YFykPEpWi4uhZ
UZHWrjni1qUjB6nkZjznOAv40aRw2C6pN543jNWJn4L0BXzJYpwT5z71KpCMVzgAL7SbWIY/A7xb
gbzSCtLPCbAfSumD1nbqD901HdMZFDjNg6fBBHMUDWGugux0Qzg/CXDmfofbUfotZyN9fvKjRWZk
Xt9Suj7c2ICmGicWbqfuy0KI8DmUmXZntMda/8XNdiVrtSZ40d6FzlI9kXO8Pv+X+bkdNVBjYu31
k/mqi/j5rCKua7VVpKTvYrWIIYN/JCG54OcNdzb2+pJcDoouk6U3ciWkbYHIZbDxHvFDUCLTXnoX
IM32n4w71gIZRm+6UVeFhP/1RdA+SpNgb4QfL4mBIm5RrGmzNXZQEcM2xPMM/lrnJzvmUvjeFK23
fTyBUrk1+TOZFom5URAEoYPbArG2feCqFLnk8SKVG/nxQxRJnEopLgTvWjvI+t9DYlier3dyYTCc
Bs0hCXJLJEi+cUCzn11e+BWPMNL+4FMut4L8fXEohZw2o/1cUwo1ZDQWf1govYz9XTkOFT6NvsF8
ztuz0J2srg431BMRa0+ycAfjghUlVXyaZYxzMMNJ/GFfULvir57fOxinuXNIwjbivx0IafbHaRg7
ZymHPRReHG8oKLtAhurtef1PXg1Fy7WHMyQC/nE/z0VcvGdi6CRQp+xIP5c0U4ldBP1FypP9mMIu
dwdWprq4/APMb6Ki8ilHib4cLVpPxKg0JsB4+7fvBUpgxLfzD7yxDaoJIdv1WJ3inXDOzInf3YR+
F2nB0uBtmvOrxRfgbQmVRRm+wz08VdKZpei8OdkuB/pQ+6qhebRKZDwu78eEDylBii88w1cqdYa2
pB+Wup4I8Y8xzz3W3gTd7VXVtxEayddQdnc3lN/KbOho7JMmfB2Sym7cp8Ybm8GudfqHrwea6z3q
ufBaK4iwbMuPa12Fyusck/n9zUsAuesB/te6ETKqr6o27cZlFXyzUX6W8YYEgJxwPn9J3rDsKJnf
2pW+bGjbUfvlXDrQvbNcN23oG7v8NxGFM4cRUS+HQDCQBkOcwE5y7vfBTQhIoF4v7rmoZ2KcTPQH
Xh3mEbJF3CNiBYuszNmMITvSoFT0fZxnvnvQRW7hH0BQVjjD7tg3OfhMx5DmLgVW6Ysqx4zQEnPT
d78JoxQPsfPu/halu1ReRiERzyDTX/Gb/vzj3LZ/Qhn8Gtw0HNBJmAX6otO3cgtoOHo9qHlzg6Pa
7VAKnDgbsl9UiR9RNS9UTRW+HyOgJ3eEDkuJVYghmGOxhGsfB0gHl3aABkbeuQh74szjo8DVVudg
2SQ1KpXXEMJBhaTgp+UtTtuzeU411jzyJf2RRnSaB1dj1zUsEOceSFflBRJrx9+Fc1f4wDNEjbtv
lNMQWjyBTdFxprpT1Tl2nag/zhMnrF/CI8yQjzxZAb5HwOvnnf9IREveYNZPkTDW4zofSZ4r3nIB
Z/7c3IcPqM3St07/MaFiKAQrXRZR5DWXsQzNNSDqyT0iNs1RzUYF5zBMTaTyj0YmHJJ4BAAH1kd0
n4IV+PGgD9bjdhiUqC8MplZh68OKShTpNGjlnRuKAhtuFoKauJmgKZ472GIfouDPwNEp8jmAVS1w
dvOjHwhb2565/OIeapykON3DsS0ASHwDz/UhiqXGa0vUbYkzBIae1FgZjYRGEm0UPuKPDJE22O9P
x+7S5D8wMa3hprvYGCz3tABRAlAVv67axpi89zeoUWuoVPbYnV6LeOqE0Vau/sn7tRQryLzRVcjC
K9C3oEd2jSpLnHwfDqYY1mr736DR9W6Ot69UyYJ2AC4vLomnzOJpRHOA23LkU6D0Mphf1CqknuBN
qI+sLo2y+3kBjGjlQ+utKOGIQsp5dlKQdgjRNepIbdcUS2q4/dGokPRajxQyHTzYnbaiuD7BCGgx
8MSpWHCPgtpfxmEvPdeLd1HMx0biXXqQ/+xxN/GXRPaRvg5t/+gX7Fc7wPM5SzGAuL8IcC6Y0Q6t
A5htNsnGz9KWuXl/VBDyN4v3p+Y3O+fZhVCqNuMOhDgPkU8M9Bq7HBc3Oe9k/6t3zwZgoQbSMtMZ
MpxWJ43Ox0klEF+Lv+zr7nGshaL/5fXc0aMhoUkVn9hSoU3HjmPuzFvCtu/5lMXA6qZXrWxs3FDs
y9bO7i+4uHEWxwWGMA/BjRo9kQDGGCQds+RtqH1f4gdbx6GnxPUel6/pE7yfMX/0acamHSxmkzcK
VoDDmdOnNg9Cj6kB973kjHLt5Cf7sIokwJmDrURu+vgzDEToBmaERKDsIviLVxOtsv2UGmYOOOmR
4j4CTLBKyJqvgaRVM8RVwA5n8iJpuNHexpH8zHltujB0I+JR3hFjnxoZe+Ywnnxh1gRw5pWevR/p
Wz95c9meL0QwOAq9eDkHf63pbPURo+NOs0Jqx1350rQkzZ+cCSG+1NZyK498nFpcOP5fYQ8Hxb+5
WFNKnZlybu6nlLX/ZDU+ukpvRourcmgZ7BfB7N2dFIQGjptwGrFSDf9QIAFV8NZFtyTa5cWN9Q/e
vwBZDLqts9tNHpuPLG9yy58mpfdi1NYJMrHHcByYd5ekwxrUz5GahvkYzj2dITabsk71wnAptQvt
afwB1VZQDdfpOtuESYsbMX1ZcBvQxU0qY0uAklXZMl8eIYEE1OeaOpPnoFYiaR9T15E8jKy9DLlM
JMoHpA/JJd/wf7Mh1LSaBfnXw4ffD6H1imomMSbyuEiC0FClatm8FoAaja6aEWZBn1o8keDTVD+9
ZiZewLYVSm3YQooPdF56df9lP0waySIEjoVLPQDnXBEi2eCy8gDgQb5U5ov8U2vgAGS1sY7x0Z3f
elgj7pgVNYD4Cq0qwjyBMzYhw4aEIuwy0+z+lHjM9Gg6wBTZUJjOZSHpkPT2Vr5ed4rJj5zWfhTN
7H3noyILsk11B58qgdJWrJD1XG7MACVnCZk8o5IUNj87ChPNLjAbiiqprUfr4yjc7NRuKMB+s721
vIyaBUC8Bb1C+H2hSHb9mx5Fwa0rnUmD6smcKrixH+dpURsOVgTtwCD98LyVUnFO7eONxRLZP0Zv
X+80G/fLkNw6haQHZLppjhuvQvpI6tw6Wkr+G5RLj2uhLGWVqNzvDCEgsoiXw9yci6qBwwabUyJL
I92MRoRzsuTUlx6BsdsJ+NcU9AawzNazshGhPYGzb4aqJ+pAQqaxkWA1UHw59VNWqaxQeRwzj295
UK8uOUQFNMeYliKp8nAbsBjGVq3vQrzdtpZrdkAxGlsP7lB7S6/hzTffQCabufEYc+VTk2+w+s0k
ek0E339bhgdDSCQxioHMXA+BNmDKxYnGkMIUHo+CzVgDP/P3RwMhhzgAPnnPmc3Y6iXyWrhOMxzi
/a/giIUCkrHcNR5MoKs/NOI74/ux7k8Fo3c2hXEYlQMb/X5fDpmrKKp/i8YYSp/SJUteK9oX0laj
7YCc4TVhOBa1ZMMqqOIWN4+JxCTZjJwm66UywWbpGJRZbIFS8pVBqXF0ZlojBBd2gsaZ+JtwzUai
NfAwsalPqIzdGmL2Lo8vPRFnCWYOyhE91uh2wKDjtqxBsQY3Cb5wjLPNkYjkswDntPQnKPWJ5npW
B8aGNO5U9byKRoa+pEfJFzDt23BZNYxHZ3M3ehk+DXyRqiqsRDU8QWmESqkgzLvs5TaUINibmnv/
S/fgeYkwYfwmbBLv+OAfxFmLVdsIJyqzCxIYsYUxieBHgNDaMARGi6YFZEhLCC0XQK5q2Dt/Yn9x
ybnlpkVED7GtesBq/6I2AeAhz9rR+Skkq4l4zj9jkl0YmYDveqTcmOK4Saoet72pzXEh9bvsq7ki
cHI/wFebS/ZeITn078vj1tsOaLa8fmYkvZdI8pRJ+KearMd7V1d48Np4P77iP2N9NIurMtI0R6/P
PSc3/kImn59m1yz07U14qkGtHNxPPF9jvNpKDebSZtoyy0L4h/k8JNZrLnHZw5Wehh7Ltq9Jw0OB
yf62OumRFcas2U08uVTpPMPtbd5g0vXjCpiAnLLEIkkTvs3k9EfhpDoaL6T1TYfQ9hDUZ6YbsSpd
7U5i4Gz1UGymBK620eqo4furzsdn0pYfeb7UanforUi+YKOHLVRu26CMvH+FvfrBZamga0C0G7VY
XLNZYZ/5gU8+e1wJHRlQTv25v3ZTUv+zevEGmcey4w9Jl1Zhfv+V6mYG4OxSgU0yDINrXsVt4J3e
OdVqoNmcH58lt7hU5Z9GIMCh+cGwRYWxQpaIosE8MJ7LlPAoA7lVPZ0KKT1sGuJpqBvZJPhb0vnj
hrvRzl2xzjVhmV9Z6/d23z63cio+0OlY5ydCO0SRfL3IbgyTopztTRsAAAdRlqBza5edC4rvn/DU
8YZBd8RQJFyuIlDGl3W6wDoL7mqYFnucnheqmZcMA55bl7xuDiIQKVmTbMMTD5QffsweaOy9f4RS
x0LhUtpTouA2ToVY9IDh7qX5egxZPQQIPBVxZ1Xs2KdFkaRegxDe29aqjnieJ6aRucYaMPkKzPPT
FDSpszWcM6oymvnVuPLkG+fUmKdFYCH7X1b7KVXGbzkWLfWS+qMT5oS+m9ElrmR0yHwN+y6NZ4fB
J8EROZR8ddLEognyuWe2Ly7gu44HAs23t2KnXYC6ryOgiv1wThBpp7vNKpce/ef1UbvgccG7Y3FS
s83Suxai73jRLAdn1HE8R8aK9iKknkCyjHtrsW+oPzG2edkhu/c1U5NFSCnyfVaFHsxgv9WRGnRu
ytD/DqU5qWl5dxRqYp4KAD6pjfXlGk4Y5LDGMovxQzIN9IwK4yXWzWVLDivqFpefIsRvXc8tc+iY
O3BBDsjdIDB3+frepVAPxjXVzyuVAYuOq2in9rYtwaOcjEMY9IRsXtmpgyhzGZ2aBRegTm31gVnG
Bp3O7I4pa1yOro39IfA0xpsBF7buc3uREXxekYl/EBfE3ldYIO2JCYhCPaem8hvak8Q0ALnHlgsr
wpw6WLrjmZhC4mgHNARgHf6J8Mj8LCqae5y5wS7JUwovUQ6JSH2SZk2808CTWb8HGRVj5zZbSPQx
bwD1anedDLFvrzpIBXzZkX5dxtUxFAMRcy6yLOWFba8/QLP9th92/LOZ255zZnRgJT33fGPb3vAt
5IDXXltCIiHv9vbK94+I1IVWAJ/CCUMpupZWKtYHneixN35mP37Y6GMxBC+OblWySIPvalF67C1L
2AdMfpu1E/Tspw3cz3ulHeWVT2QeWtZ9+0P9m7ZYHfKklPDj/Pz4miTXiUZ0SuPtSfg0Ck+7FyNm
y6O0vWviNwGFuT+z3p3DXI3nyfRsNYCfgdIgD4Ae3bREBwnBAiKucTuKI0H8VMEEvjB94yB0VJt5
ivWS1uIkirGZ5U3YBlieLRZZHfphrGFfE8Azf6KSnNJuLgT4BGNm77vZA2GsyFLxH6wYkkBdTGRk
ctpYVtJ9fPhfseHTJgKDVHr/KU3NluJ/mRgN5cYq4HKcz0WAuTKG1zXJsOhSzZRQacVgIiFaDfFM
RWkumcaELC0ZXynyG2Gnng2Lkxt52fatLzy8wDxh4rGA9SpIgDJAeF/11rqBV2uC4u0YJbcRALNC
FqrojC2bsTAZdd5Osp9uTFAT0aMKrL1cyNhhxfgNdOMt/tH3xJuqyJd6zJitwfIYin0QzDM8e899
hjhK7wwMVWBJGd92XRjnzUhTsPeklRhZDa3drSBABVpMPUSEdma3gAKT2rjg6uGNdb3CfvnvY23Q
m76GQZIrsVu02oSqKK/JDdfrvZz2MWnjL4wMjoSL43VlOo/NGOCpj/jRxHePV1yYJtnrxnyCOvMv
1k0rUGW7hWT/cBq4A9CksiCjZJn59GPLnqqyctFm9YKOxqk5FBE4fEK+Vw6W+XHRh94nPihc8eXY
mSH/XUzldFZIL8f5KeFWXedVhoRvSXWWmsVus3BJ7rWf+ddukFuluA2rWlCrdZ+fJNCa6Ev/kqZg
9AAuv80BNO7UB52YgEemzSqyZCv44tmNn9ieiQH+eYBo1tPCsnFcO+ra0parpYN8CbWQRdSas1/a
4ReCQVLvlgAcFAKcj3UTltOgtB72lZBfMa1A96AYHWTkE9V62JYNX6koLOHMTnb2iHoNmxcg7UIQ
GecmuFPjYNxmGfLcxMTanzmvYZiu2QATTkKktKJxC7UFpjJKpabya1+Jp2OR+ZUua4atkatQFntp
Wl1KX7Xqvk4O71dglY9OKanjOalZCmoHugnJetd2WeRgw54BQNQfm7yUXSTHJZ66byOaREB3sWkL
LU1/np1YCUNIz6FJME9vxNR5tRZsDfncFdwta4aGkOJ7QBcydHLWv3frfxXu/h9i4326Zjx7x0WB
oAViyjdyb0TozfS/yyz/DpCqxGwDStLBOH5s3BvLaKy4PoA6Qj+dEUlAt+lxBqBqQCjUA1oMmTDC
ZCEhoZqvVqoHnMz49I3vtj98+SUzNcf2mF62GEWKShX7lF+3TDtU94+Xph5EFMzbnByzHACZXdfa
aHxnFQ4tshiM0OjjGLQER59+zqcAKvfjH2MqTz8Ho3sAX7qK4ShxjeIJKFSb6DPITP3k1TEoj968
h1i+DiL6XPEb1VWceVrcsZv1gFlWpO3FgAfpf5jMq1OPiLGSEryVT5PoX79TNB1mIhYk0+6p/5ZE
uBlEufsWMBasI22gEAhKyBTwMp/v6QLJQEQY2L7GkYZgc66Re2hvJoySR/PJRmh2SpJelBpO+U7L
8REEDNMJVLnl4UA2+p6plf6/n+jCLjAWcFxZ6xpTGeCpBfJJQi3s1gV18WISIB2Zikq16GStqrV7
04FpsYVOnUoE32B7ssc+65gq12qeVDQ8xGRF0udgY8juATJjeZ0rerwuBNxBiELZud3i4ItqcHIp
NTelKNLMytErzfKaDgHNnKBslrtCgjcfoPSjVThOVaxyips8hEVpPD3cZDx/JcbQDlQ/rpUZi+ok
lvIQyTzVsoPdhZumrFcThLT7eDP4RlNWXJChfFg2ErJWy9wDa51EYJn/q//hcVqa6S2VE4S7naLQ
lIZ+oU78PoizD2TS6ii7YB53ZXwL60xx+OJf4d/4hBwXwuj/VfattNjUIIf22bqb/WB5y44+jBn7
vd9LoyLcZHcHoEDXg+jnqMwf2+3+AWgkkOR16JrPfgyr7TmD3MJw8XuVqBRFFJUoEKt/NLJk+/Sc
be115R0QEkE42SFetqtNkBdrnqE+m/7U5R2PJbIRWDtOAOrwJa1xL6B4BtnRnZEKFzhEDM5jxGuz
fww3EavDQFGW1XdaJ1m1AP3Jk+RQnvyLyMMrrfRRo6D44FwqydPuTF6ht7dmlT4nCO5dG9Etfs60
aQm3w9nSXHOy4sRstlRObqIcAhOXqk+zWRij7MJh88qstYNfESsBAXNPwTfhPiACml2Dh3YMqw1T
KsL+W9CuCtmwEH6jQiYjdZ0Wkj7QBp5PBKiPNrA2ynGKmbY1pDsoRSRK1+uobipGtoK6VY93CD5q
2GVX4m2CGYrsBwwmdBXjGTGy3vo+M/j4dmZsC8aqoP/U+OeFwtCgPR0oCciiickckGxMn1Oen9yR
UUDOXU7l4QrzSeP4B4qmeMBIiJLR9UE08F6JvsUUoA5UUPrMbXYG1/o0HlNk0QN/re4YZldiZRYc
abDtG+yFQHTsRuirWaOsQfEzB+Y/ON7hXQYBYiTdKpCdDbzJgJRAtkjGvV8D1exPmamiU2nRtovo
YOgUx5o3xqpXCPdE1qmskz2aOJyKzf05WkcqmyPbF6sg0mFAwx40MaU1dAl88SwV3wgnbGbgWaQT
DPlMDybI7qdN6bbVhPW7SoSKuO0wp+pieAdoCb74pOIeze1ZjSUEMpn+QTJJZTPoTkSx7gRbZ6Tx
+OgpFm2nCFA7WcPiH3MAF5TMb98HOTpXY9Hqqm+xUQ7CP1qzbuXQCg5GGlC/oTML8dA2wS+NjFYI
hHHL+PRwSdH8MJs1DrA7UAxFjU1UwqL6u4gdF8LSegkWINOaEyhh2q+AXCAZEcvsU7iZPudxDCyR
XSVZ73Qj4Tu/ACroO6HYT1yuGhdFFSg6a2iNkwABDLRL+bJpibLUbt/GlFUSdx54d/3+tr50W6UU
e5TJHCi/nqOTg5JJtHwDD4QRRgGwJpDZblq1NtiaZ6lANGI5K07R3dj4tfvzlFmgNJEGUMGegcxL
YIBTeQEf9asRQNNgH8XJSL7HwBglMpDpoUzeUOWBdUHmmHKEUmq/9JSGEQSjLlXAvftzPplPiWLa
MPdMfF8fZkgIohspM8PmIAP0RCSsYS4SrPQlfJ72WB3r1SRzZkDZiKOmriY0aPeblzSQ/CweXVXz
80yDX4IWunrMgAN7LRJF6WtFa8sx1ger3acyT6PU9ddfGX2WTcDXqSzZcnUOGJh4KFQsXbBgz1Rs
FMxdiZFI3RF3Ndtv2x0kvzo44r5wnWoKFuealif53HPR99s+scP+4marH2nan2IIVxEASeNmt1FU
VEFzzaAsDfv1RF3VyFEf68B9ZLe2tCU1lKMvjh46ZsXz7pKvftGTa15kyPfLqnSsV+2kOUN5AoL4
j3c4AeKzyjZJYLObFWSSzBD5H5pTPBZHZnDc9QUF+hKQ3HZ45414W0OZO34GkJaFXdCofv6Ly46n
i9o0+o2IxYsOZ1lwDNhSAHGzYFxCmAZVkhwpkGSwwn2c3Jn7RzJw4j+D2peF86f7GgmcZVnil0Aw
CsLQRGCydyh1BtPjY/THAZ7H7Z5zDpRjgKc0oX9vsp7gvzroLQ9SRRMcsWhNIoBiQ2tuk1x9xTv6
jc1AyPhFqIhZoVVnoJd6tvmVgbf7i18GNdSwuL0RyqZiqM6zk5w4A2yb3cf3589THaMygoeFSYZv
KtA3Sy1aOEcu2J7txHIR2q0SLScRinsY+7GVoCiBIlWWKvRqLZfz0k+uN5m9lgjD0YQLXn1+z1XR
dg1vbkagyei9DHhoYl93K5iERPFjiQgnxrcpmGqbXj9kynM8cVlQE0ozVnEg0x4xAXGRpKCSzaTy
poK8Dc5zj2EYKmwoWJIlDm04pFZD8C/dkzI2qj/orfblcX2QqyIPEboVEcAN3VtnYagTFJfVxA3w
gwdg9CURVvyaEy1p024lRzwP/kIXFZu3vFOKn6ReRDJIB156tv/jaTTUHeiu+juTeJYWzACWZlGv
IncrC1oxjZv56kbOF75KWn5hr93+THeKfn6pFKOBxmxLXq9yEsBPC8lqpFm9YrZOAduBr0dmDtlz
XEm2cildQT5tNw68dWxA8vjIBo0f83C9pEQUlZSGoivPKgOX7ASpgx6oYh34XRG/rqo8jFAHOzVx
x7SedyMnjZ/rqcLWDiScnYGgOjq9r5gtGF5x3g3xKAe3v0EEj2P8DCEb/XylTRBsRJdysXDw1y69
NzzM8pLmoHPWGiKT+6dX4B7ik7aNfTzFu2kVk2dvhANZlu8+ZjhDXAsW0RsvQEM+7hTvu6P+/rFG
MH5vMsXe7282zlqSIcfShajGAWLdtLVpmrIoXQWZolUnar11VYvjdYm11B/qcPlZP0e0NNj3kp6M
RCIDtB2yBM+r/k2JvDMAfHPFfIm7sC2Ww90cs6wpZaBqOgpNRGqy+/gFgukOHzgsKqtVJxGUNQL3
kP2l5XZIN+O3BaUFOjjJMUGfiziLkKewWkGnQRkYTk/9WyjDD1ddOUd+sxqndprtL3eIplwu4+wu
Dh9fhRPChvIaT26VS6LuCurXqyfWDq/4PK39ZmkqofPo++oqw1KcFF8whvcXmejaCFeag8QFTwi1
nFwMLj1U4Eiazyfal4U2N1+wY7tlfDS6Rea2zBOaBlxPGeLRu8Ff5z+I7IIU4M+WPNxJaVBUsaPF
LYP1mO0G1lN2VvDdZKvqIm588PLG5pYGoBKp9O0CyuWUvv/G4JLdgOy6v9D59luuCrf932Lz20jm
dEFjer3m/33s2T5rmqmIBJZvFFMTK7eHs4r1qk2u21i+ecuP3kZLRR7bQDHvbilPB7qZVS6kEZOX
O4MsCerv0wtw89ivcrkwLB24p59xBUbDohiAsM+6E1X6skcujsIYY7+flej/CynlvSEsyalXdV4c
LGLfGPxLaJuFInbLydY5jEO/s+X1fekY5FTewIrhkdhjH5n5GT80aDT5GjhQ97dcus5B2XS0ix1N
tAyvGTaVWljjgcBXnQsjfF4OSzxEqVFjYcLmhav057juv0nY62uyOaylqZDHotCH7inGr6o/hQvb
mElX3vhOI+7WU/Mwelf8ZC1e3Y1veant7TAChGn4r7gr1Tb1g3EnWjTeAsyFvIb1ajrcYV4l2Gri
POZkykn2cwmQ7poXvo7M5XuxlkRXCIS6G8YldD6CD7CXno+pT2D1IlTT45GRac14gXROHxrIn6cR
HKEZ3ekycabYXTxUCQbP3ipGriYt4KbNLsHBSzvFpM+k8r1d10G2g2eEhhn5gQ1DeIpDrAyk1zBU
3y70/Hcdu2YjrDZSnQvy0NoFK3ywMoMMCbC54Q4t3Q+7Vx5CE3pFyf89KibAIkvpo7WYNuj4I3I7
D8SL08ivbXh76FaGKrHMVa/qdJLA0wl8VW1n82bxbGBwMjhIyaJNBMtZggGEaYi6rx9tXUvRZOCz
o/Rywn4QUK64CXh5waiRm6X96M+Qa7K0V+FYeWXexIEaUxAq0opiIiildN80gpkOBS7oiDZ4BSYh
Ijd6Ss1lLJl+Xyx0CGQhhaDgnEeQvgYoDfiyRUxRQ26CLWvwg9w1gfQgmhoZmZ1pwRrM62BT1MFu
Dv2CeXAU5xmQ6R4tdGAW8dCh8jrmBitu8C7GTTu7GqeH857YBxLvl3URbL7I9Hd6P7M15kyaHNUI
wTBJwi0v339EQjJH5mXN+NuSKKDKC6o2Zn3BZ/moNkJfSzXsh230PnLwCbQ3WXdxPt8FU4jIwxzG
FXKJDXLNdcdtl7kon9fZx/ZK6Oy2KyAfYg0d6D73t22lCvKyFTT6qrnDDHt9W5xow9nwf3Tda3DN
Nrm75OoyboLAUuXGtpfCtykk65DFPC0iyyvDktbJHUujUOW16Ns5wsNHk+P3SnKVRUve70M++wFD
oSfytvrUWvaQ+F7fHKLqFS/kQr3eCHPNaK2JjJRXapzG4DTPubAfq4eLBGXJc1X4xsPVaFPsqpRG
OkfwzXSPJpvsnB13jLK9H7lCPY3V0IQ/qF+bVuULHE43MitP7hZf0ZbShEsaAKWXS6vdbGtGe25/
foot8yETuGh4f9OcY06upxTksHnNpv5A6dXyPXS/ZfZM2O1+0i6VNmYpZMxSMu8WIogdmFw8sDKa
avOvbflspIYzUb5nAp3ch/ofPPEby/FNBxA9bbJTX0V/G8CL1BTf1qIl9zS98FCO90CoB5EpDbrE
c0ixviOCWXMxDH9L3LKA+GvzO14e0wc8FaiGwMTAxqI1puhK3DwQ9v3oua5ZF7un/1nkDLkoOfgP
FK0rMTHtX/Ce9NnB9hOAOE915DIas4YLi671E3Q6YM4kmgolXYdlE52tdbIjHL5ONsrZZfQT6EZA
hGv4tCNrKYRsSUWRsiwMkjARt0VJ/a0ozJlYw67URvXnyJPFxK1Q2hQ80KPjW1zYV2PTUlO/q3OX
vynBoO/3VTUhnVlKccBkFgA/tIUcXKfgcDb8sw7uv4CxudEl9X5aWxz6d9cqWvXw3cVeZHpG/7c2
0lKGpu0O+aGKUahWSTorNjyfUnrQuJQshKrMFDThvyAFP47PzKRD0zuU7X25HI5gPMJWxnrKsHxK
e9aiHAVxVRKjk1/4W6FQmJJb+Tm34wnLS/4sP/WnCY+CtJojDSWdHPIhHOcNldeptTNq7fIp3iC6
8ltzgMheF0VTZGvP8Vykajd3TVKKMXshh80Sgmu0Ej6T0M/BTuOr6i6vVqt0dnwTJK7JIBIPLDkz
ElCcltxFBfwD9zH280LJ2nL5XEI+KaDMz09B2foI2qtDqb61EKUYFsmn4EPEbIUyRjDAMVnan7o5
83O3VJtgndej69BWTvRJ3lbvGbPdGy8y1wsVyfcF9hPEa9/+ORFEAF8yT+ENsQ8KcBMliYwDMcr1
Hfbenr51pVpnlQVXNCmfejp2W76urATBId3lNZvHZ8tZ7KjXvklC54IQpIdAED4oRmD7gfR+LHiu
yF9mykJ5rPSY5tezlKC96fSf1GgrywHBC3z4/zlegkikP24bAMXwvuif4XEbNt0+HhQH6tQbS9zx
AzUzRsYGAPNgaYfM5sQ+Fu/D4haZPEqSufrsnzIfrmKSwjXF2vi9c0dVvXgFN+1tiFFxGr/uoz0l
NB879tGLvoyUjMW1mtoLLyzoATi62o+psMto7at142XXT1qtn0Rf+OnSESb2jXadH9MmCTNKlkfl
RQjucGDQ9s1k6t1uppACDs4qUsSm3qINKrXwbhIyEGgMfkektitES8i8qt6eGniWoW+iixxsD9T0
+oYO2Du3Qg7FSE+eJKPYfsjQpDonDH1ZHREcUCbfZcsUp8ZaKIEuJG5mgUMYJZmpZFM1iJcdCpnD
DPf+zqxW/N13davfSRJXSugiTQvopj43B+JFwJotuXpFUlKDkiOUNwYK4E6JpZt2hV4zfRB89J0z
nzgpk9StL+0JsNoZ2bU1mQZN0hGvSQ/BD1le9yyWzb70uv69iPU8/27aXH+W9jJRng70k2oDWF4Q
960Hllc75Xma4qC83iGYb9yIk4YHSVV05mtItBAUuOZChTzETUg/SA9ypeupw0OYPd/FOnTFrfag
7tTI6Dw7ZfLpAvKFYX4xMkroYerhPOcoq80Qh3mdHtR+tuee3vTfhmNzmyToAZZmMaBkTm6DXSv8
QzmJYwX78ANKmiH3MQ9GAVbM6qFa7bJpMxZfwkNkzi7lQhy48mNqXe2I8FKbjGcAwVqCu0npvM4F
6Dou4MW63W77pIxwJ3wcj6gwcnyz1kbazaikXrkV27qVCJ7E4FAPc/G6XlHCiZM8dMshDfj04YPv
Y66GkuGxJJuaQPJLzvOwaWxq7sxYX4zGA3PsDrjeQVWLHz9JUdAz7QaIdOINuhd3GNoAnyUHGzM6
kE4jsKdLamJyNth+xvEzhY0Noo5BM9Npkk28h/F22fjhlxyX6+0RKHMtMVRPQnSLUgMsrXeEjdQU
zRkfpgcmgdo+P7DNwFQ9Uqnneldo7yoNxSuPYcHnV+2k+JcHp0D8bhIC35sbUOr6Oeu49fcwyS1n
ZQ88UGAhDEnazXEKqcGRtJOmDC/1rbruN/i1DtRa/Kxs4fQbhLLEmO4LNVRr5FQP3Wu+MTN4l+zE
dpr/cGXX0ukvZRGZLlEF8xNMpp5V45xOfTXga33HKKuntDf1yYS7oRU4kZg5FmC6dqG2sDEqGUM6
Nomg+YaxBkmqdPf4pPp0UqiKqI1+qZl4GnnFk40yNS9tpwDa43BF9FZBXXTvO9gZ6NATHyVWrHlk
GUZMJ5MxOxmuWILHibFn2CnezDmWICz3Ji2D/LiU2+C5yce7b+SWgg6lwyVcWH/1+ie0fvxcaKsG
0b4Afktq/uWqan/0H4hR4ZjbrZfW+ixnjz75LeJL7u/GRA3AbnFs52cGlaNNJu0bjfvHdmf7308p
JKXic2NZtbExMXVIlKaAAAIyTU97Hr3kyybbWKlY4Uks4/qMuXZC4tvVL0f6cxQ8t2uKdEdkbkTR
6MWXESemhf3L/vJbtYeK7RWtDoK3DdjsiSEnQXgVqPOufpzyOuO9EbIa9OhhxJVlU8ZKB+LLKe63
u+8+/fEmbQmftNu5elixZM83mE5LUe7/41tbduESV0KBMMso6ZKtzmznEyLfoO0JYsSE/XOF8gcN
S/SUYK8RpCjCT0b3FprVfGAKfJqVA/fGTn1/kJi3a7j3jQC7DTRoTCSmgfVm1r9rW1G4alqxPwD6
a39Jhj0MZe6LcT6ZKwdRIYhtbtTGQsfvO5LlaWpfpRAwUhwocYDuWjA8K6aoXTmaytVL+K9PmMgg
lUzA3Jz5G+HagQ1VXcGeTpaqhbmpZbem3Hyam4y5eZ7BwSh40tWtCwJ7IOVgrCCQ1rmYGf1VhTsc
1jc2Yj+BgwLVOThtbsWsc0oDfB0D9X9eCSsKNE/Tx3+d0GW6C2cJ9pE41Bs28vkTb47Pxk4S0aHd
KFkx83WmOGaBxixmlybnD+JWR6H8p4Eq3li+qZYOIZJK8bmHPZ1PYBs6I5W8Q0l7VFmflfDqGRP1
rCmP5Q2EfgDZCSOfGXuvr6Y0vtBrpGPSwcoOYGtv0N3zMZMVILu7UBQBjC0bHJ90jEknOD3S52ck
UQEAp+9aFkCgfUOveHb0JDucguqUXU9hcfWSqibVJaW0824mdVnLPRJyvA/UwstJpuhzScpmmXDA
rSHyUeCBe0cWezuJuH8+DI/BF2gCIwR9Y89inM9aKIs4zvMhqzoq+gYvcGTjN0L3XFh4N95oF+Jn
1e7Etxmx+8LeTevg/UVqNoGY7Zuu+lik+wK9wfDXoUMVaVqVhs+yYRfkvfi4mYDZPA58PxPwT85R
rSXNTMWVRAC0YqZwoD/kmANRumlPw360Qj4A2Tbup/1ohfWsKxtfYXSpypcI7JNlAO5IyakoZqpl
8LPUHNKcgQCo7KGotoI0dIWnT2/4Q1yGgl92H2nIDfpX5GprhWm5b/2L7YbEe5KojC8u1NeNk2Jc
3K0ckisNuBp+hfA92sjuiNnOfqQgML4fwNrYKSs6W1QjorZyKm0MkQTDdTfPuPCcgpazRM6yJkjt
5QmFUJqe71gbsfcDlyE8xoxMLsitUjQCmGSeX4Ko5omJyS5X7ERFhTNy3U9gFMMJSbDwDAlRober
ewjpfJoM4UTV8vf4WS2JswQErzIn+G/XYEBqX/9gzKm6g97rVWFlW0aaO2rmB7xrq9iMZ1+43juk
r0/u0HpgWBs7fD5bu8M2pi/bz0DL8VXVRDxrLt2trBJPEgGA9gdz1WRYCOeSLOWoY9bp4XjrOvD9
yajseOUPNVjSo0UWUQZ+0oVeq7OOQjx7/EwSZYODBa+3qONNyoAMyfgjlbu/IHQZEfQknZQlOkOG
0xPmPO9UOUCG8CakUFvMpZg8lR+SmRNCm9c1/WJwB9oU49qfj51ytn0hRWENobTzLzzv9rtcTvkm
zrEaVjSJ1piPK5U5UuDfzvx88sLqheMpGetmBdI26keoUS9DkJSC/8d/o/yP8qeBqpBdxt2AVkbI
O6LmZj5R+fXiBSEeKuRYTGn2A4+dAirdGVt4X9io7hzQ5Z0IjHdVizzcm6xfSADTH6zgeKcMPoej
77wgyER0A+WA8FB/C9Lzoflb+L8H0f6jsJWSNjQ77maWZkRo1hS3GHDS9nw59S5mJmAMuD0jboNQ
ZPuUXRfhsZQr4iV+VFcPgz05n7/zg0SYVy6ud4S97DYBo2achDGE2vuOyzlq0+MXUCeavJgGQpkB
PIayHVRW3tc+dsFFf7SF4Ew/k8ZojjLjFL2X5kpw6nxIx6GQlG29gQ+4VyuijhbTl4hzUTT1nVqE
2dF89szt156Vl88xgujGFzRmqkqjMegjEQq515uHbINHEW+3N0jF1UaGcgXKII1gfPXVrJfp1fMF
q4DScfhb4oVmOjaD0U/32egSBptudt/qM520qZUU3OmIaHFMziAoAcUrR+DfVcsiL/iQ9y1aHLkE
G3Yn46I27+OxX3F+zTnHjoj9Bwrr0nzwPGY8LFb61+YLPv6i2deNXqDG4Ag+/WZG6DGcODXmn80E
uh22jIZmDWZNgbxEtfnqyId+JnZfM1BA/mbCrV5vd6ZkBm//C68DAOD3cm4sjoEprihprWoOAg01
keifPeoQS15Dbc6kiW2LdyUDjC3I4eZxzSQsXSa8Uzp6ke2UBbSMGBANnUF+F+A4j+qACuklPt6d
9vJ9IIYYmVoJM8faO9oxTD7bJvkEl6bSojUilzjEOXvV4aDqm8Gs0qpQJ/tsmo+auK6+iQMHSeQE
Sz/qie6iquyVvsPNDmXlgX5DZSBuJhVIoXk1OL7DvVw3mko34sPnqqg3/aVTM+57tagbi8Qij/A5
Q+foC5UZfBhahiuBYRstrD6QIjPcyUoysgI+Nqf1Z+qTZoGmCKF7f5a+fds1FK1ffv6fzWUPZlLb
GTAdBsqYOmazfGaXoqTW31gu3Ws4IAjoJokVSSfkeu52I9QIrM+mrrRahk+b6bhtWiQ4Cig1uSyz
YZXRpT9pgHpR++Ui98XloZl5JGfjAZc10l/gPlJVlPk9pgfTxx8sBUGr81P4oSlGl1EZUWbxJtXD
w084O/iLnKXR8VhQVWbh37SxOfZwrwlBOZEyP/+0MUsfDBQbskGLjjWLhJqPHV/049rKyHEUS3Hh
0/o+IYnb7AsuaEDrQtaIuGAZ46v8YIbtBmPqjGindabD2kVZEb/TUdMRQCghMemhk/z/tffA0zRc
W2mFLraLJVrr42DMoBwZbILY6ih+SqjPebD03lJZlT91zbudV3cuO74oggfsKbQyTr7qSfcF7Ygp
IJxZSWm8AK5hUyU7823o+2gDGlD6uFUKVRLrvJMYUjiB/uHELCNvm2dyuemospIVn7eaKvSElEZs
ENGAs7qkEKkqY1WCCCmjy5mYhnw1p+Q5ZcGXATLQbcekA3Z3dCJsU//nXh/N96fPg0HAT8pAVUvC
VP1dG3Rz47uGq3UvR0ot2ixPXiWiiJwj5Ix/O9tXLYAM8sShNLsztOwXCU+ehWROWf4v6xbCNFfN
Cax4BqnrOmySMRvSzFnxR56hKB3sCV/4ufXza9euIxMA7OX0KHr3JsQdbfFGqSWQ52x2VmUhKAuP
nJfxxxaQeE4seM6o2ZxQY0Izv1SMwJFySCrCPD3J998VSYdC1DfPRMg4X1igRxOm26dfmeCNk1O7
prFgEGXSkWcTarpK8HSAx3HKPyqY6QptZkmWd8FC045NEyq+KCLWFxg0uO9XbhKLR5uo49AwZi+z
m32oSht5wFixaRl6vZL0ppLHqLEWUvmUeWWm3iKjPKZfVruq6EsY1tX0T8O4kRflSMHIWQfsgI2S
htF9F6VyNpAwz1G8lsviQ4oUUWpsnjRb20pUykcj3hsg3IMPxIXht0elM4IHivTFuOJjA3A5HmHi
ZudwK1Hq3HCNYao5jYO4xhVIFLVHsk4/iIA2xROPTn1WDdbyDccoKkklFwJQUhd4qaMf7CUigjgp
fGcyk/pQiUgwfCxrb/NCKqSK72qn/kfuOFwglgIVHdSewIzu7HThH643+bt1ASEpMqqdkxb/aRwe
qKdV/6RAG+IZO5r4GczIK7oMss1dWEyVw9LDs+teh+KttIt3ZMekB1zEi7p0OH+rwpUMalUtyjSX
p0eIBaawQ7Le6LXvmhqyoYRtutdHApUbzZ8vNVmFhFaWd0z2xj0vKH0qw0e6ky+3WkwlDria0xtP
LrD/5D0Jz0P5Pqz3Q3O6MLz+jyVvBy54igOuGDZ2dA2bMDZEsglxJ7jufEl+m2V28QjkrCALtxjO
xf7n+72x+grgB2gMrBBvBs7dsryY40l+asGyiVRoXo6EDepiRaxU8tJjIsS93i6SYKfXi/kTvvoj
Ld3oe27uqONoLtP7uUB2qXcpUDXcwn6jTiMuCgoakXI2eHhIbgW8IdqA0MUtjg502cxZVdgk/wFJ
3Z3aygFdtM7PfFBTdO0iQ+KVpRbyb9Y37OiU4xnhGhPIXrGSEJV4aNkM8uy0YLZr0BQls+fmzovI
b9XJ2PyAGpAqsPbPrA+wJGYhZ8PmVoOtKz/nl4ZJfexVOmmPKnoT8Mc/QO7KxalLVWFSWQ2cVl5M
Ho8eDDYQ9gW13m6hR/slZDrb0F2mRcrvA8NZ7I4lejW/cQ0mdfWgdm+sRQx2+SS7lqn/9NbtXx95
QpMFMIfctR1JnoHFe53Kb60o8I6OKPhYaCGfCF3jXMBEpvo4OizMSa99SP7+lqvVbMDmCSKQv9KH
umI0cHDzzvRLUWRniAM7q1QphpmmhpjI1d0givTB3VTFxvw2omfSxYHW02WELHKuWZpt5i6kZFG2
rwyWDPDQEe056EicI6w4TSc1bPkVt+jTaON5OrCpKIVawQyqcTuYaFMirkE4AEMreWhYGaWKJNjp
7/i8OH0nHYigOJ6Z7Jl7BxkVSZor+xiVnVrfbIQprkUtbobzbZB4wK7jfZfA0wNQQPN/6+564R5I
HjdJmwpTNXl1qm/DryMpfKdi0018z7Avq1SX8cVR+fIpzFuzrjc7vUN4t6i2JRVo2/b0hxN1yWqR
5IcgMIW8fFDVoe75fmwazY2uPbiw9EmYhc53qS9NalS1dWpIL9PnCaTRv1uJay6IYAWfjmskW5vS
kGTSZolzsoo+HKKlOV5OpDBEHiltVLbkLo0xJDPq27+DJM78dY5UK4cRc26P5V2xZWCAbYrLOhmm
DNFOVf6LVkK6mIa4QZ7yZ/+D53azk8rfrgUuu6GyFMT/02TxCla4mFx6Bc7F4GkOdVW0n1rXc8sg
ee0EKBj8MAmUpqZ/2ZtHdcl/jXlF8kAazuxPT9odVpg/JMOD29bmrJm0K30fvzUpSkzlSi4fKWZD
fZQoTPewPBZ/rq4sS007JD+jbgmf57boha2cCtwC31aYxdUfpj4MxCEvaP8hqxc8bnDmnOQbOlNT
DN07FXrc9T+yBS06VSil1fFDJobcevXFuArLyuM/e8R8TxZ5vhXtVGkveYTug5S/e5RPCyheiSJZ
bt/Et8F3y+97WdUzO1xq9iBcerSJqHbiOWIke38E4wEILAdxod34xKJ+0Hx6ExhjjFsiZW0e+0Cx
priWhMkHN4u6jyFgfbRbLgE4wef8vHkg/qUO9VrFUEoRVrUunKr4r8KzSEpeRFtDUIZZXTfDTkQ0
05WT5nUK8wzVX8zmri8JhWs1yB4bDcpv9JBnEQlUYHrqzTa7Xj4X6dkiYp+dOOe4ub+Z5MDKXJEx
YrXi1Tr/QLKgkRKVH3s7S89MTnH2TS5vPM5LzeZuWQwXq9cFG9/JDsqFS9KIJgYRBPgV0kqDaaZJ
ZPHeckDTVl29zI+TYSyLS7tuXX5+GQZGltJBLzBDNkaKLeHLFxdJXicepDzG6FasJ1vjVltaMiYz
NKdyRt1pcWyRbmz/n2cmz79OK3mpNXegxrcjDcCzOp1c05a/gU0cJp4u2N/j1nWpGHa51wd5BxXL
p9fSxxgj+ytH3BQQvYO92dEEns0rf7NUpAYi3/qiLEIrn7L+luEKYzRByqxJe0JednXYMFsVyBpZ
xIhfeqW865F/B3sP2gJVn9Wfo2XYJ7a+rd5gjWZjQNLc77NjztB3cZL3pW/1zhMFcKVcdhtfZjuU
/a4O2JqZlLvk+5Ka9MCiyBFM37RTaT5cId5lbS30Uo8P7iW01RXyFcqC94oVzZF+af4NT7CG92b0
4wJgjMPztduRE0WEsJ59Ud7dzPrRTgHFsG0O14P0G4XKJPeTN+4NcHNE9HaCdlR8RHF/nWdPfmpF
Yio4453pEyF14lOuBlRfTQy+Wi4/MeJPOYtXGaeUIGKJ7TJ2h+PhNIjWjZK6Nd2LraSSQfTBDeA4
PK2j6MuS2tSxKpOmNfK6A5nDPYGooGa4IGcp/Vky3ZiPgpFcdQxvt1YFNm6u6E7oy0AxFgDOQyzc
K07j4s8HYVqLIJET8d256QRZu+owRSFDA2IkFr7S5xYxHzn1UUo4UEY7Ex6kiB3AD8d7dknBF5kZ
rdJ19PUVccghFcErRIWfJ3cnI9XYDMXuLw8fUqvQNmv9yfaslpZ4CUx/Pi2F1iYDcba+Po7ENx8E
IDnNPxJjZU2qhqoWeIhV09rRyobzLXx4RrVKF1+02MV2fWp/Hc/ZMNlCBQlSk4AtnGkdRGfxnM0j
9+x9fvKygMLSPjEvVfmzi26uyQK6HKYQdBMO0KhSbPSuRjG+UzgE2eBmap8qzX8IaA+n5jZsvLJe
8HIkiB81S5negvPwKY82T3+90IU4U3QVo0tP1Q8u6YmwisNinqgosX4jAuWo8VY11pMQQFzPKfxP
mExgGzsUC86XME3DhAvxEM7Z1Mar/Bu0QH9JsZqoIkzXYrJ+lqMUOBivN/EfV1k/lw0zXI2QIprz
UZ/xKSNG4Mekz/MO/VNHuVHmMcwt9QoTQL7S2z98D+y8eR3utaeT2zbVvjJ+A7P5VkFquf6scG6r
80nM86If0YezqsK+WRCv7wZ/mJpVSHcNAqhGjogxS7pIOGJPYl+qakF/9TAIH4MeW3gzPqQ5RBsO
X8Nancmn7Jc/WjCt+izKKSTbj5BXJ+jwt39umDqEH/qRwPqvRO57p131ckhm6Voia2LW9K+m/GBR
nbgLvjV2rWyTQ7OleBV7eXbUig/9rn4I58+3LBeynZeBIOVPqyNfZF7foOsEBsVQYr6sctQYk5ta
I1hLhUW0lHYkCf4D/Ub2fXh1oma9GdhM6K3IOQ2CdHBTd08tqAtnRW+e/xAIbo5HkSjCX9O+JJ5p
EBE3gnVZ97NIEQD+CcbIj+kt+UfUGpwLU+i88rgMvBrMIMRn/pAeJ3spP0JCwHPdxZ0nESBQy+gm
fu7TN+Ma3hn8TwnbrDnC9ygWqCb9kmh07hkbPqRZ0V5AJM22D+dmPbGzg87KqHrBphgzO48EcWCe
rB8B6Fc9pn3ZJHHGoBCJAOFr/aouFjigG1zf76fwqwVo2mPJJ3DhP/HLSQT0m0InK/Vzyuovr4yF
gz3B2g011EjKPrTVLmmLHOtGbaMPB6nOuO+jprCCgvl5YnKfzelu2isDSWr1ir+cdEeOJCSTfQYP
3HaCaZcqWE6GNC1zpjTrrwoIPjZc6jybvwVqSsV7zJWJ7mQ7RgomEpXlL2fUGQVMSXaCeTQlI3wo
7FdLLc3gIGw+xp2bHlTlRAV7N0Xj/qS6+sBCxtIDrDLnypyy2rUnmTfaBpFiadLLtzSYmP2sXbGF
ncIcmxDHcnOov1HTN7nyu3rXGKG/dhsCcj3USaQFxU67CNkrobF7EtOAr82oAY4Wr4vPTDOg4YfT
T9Cp/KOdZ140EL8hpgpa+GjpGI51eBuWbOy5m13Z4RLQoNOqsOC3uEPWht2E7Zqs7v6/F3dSjcQu
Y5fJMUNUCE+Ug2nH9gs9w6QryJeEq2MhuXkrMq8TtMFm3k8TJ83rWd9ddfhPgcXofd4Iu/ev5L4s
hVJ+xXuP0S6X20B3odg7fY4Ebo85QfqiolKECiOTp7B/75Wk2ACcFfVPVOwIV7R54PQeiFM1ciAQ
bPR/X4T9GwjJ4d100OBpRVJS3uMY4LYaY+xpzhkF/mqHzimi0VQrlKNzU0cMewDC0WlFj1NIC2/h
le0aIdRPN5fBxtOBy2rtw9CieKrjDt3s2IU/Bhqzp5GQl0x8MRwrj6Pg1Sfe4t54JnX8PUbqkjbY
enz2EU7/O3/tkJDVYuS2r4poDe5dIpGNOPgkEj0o7nVoATFruVE0ihzvCFiaPJsZgv5t9uYrsixG
AKtx+xqmlsYbiIFe8/Iwa9bf8XeS5MvmZaCuUq/z2FnrasjyJyGlKkYqIjyNvTTnvRytcerPY6Hk
ixF8Ia61cCXnPpjDDMFXjuzEEMRu2R7LBC2I7qLALp++Zui74BCcENJGcvNt3vmW924LOtlRT6RN
+W2nHYSt+MaUpE9hJ6rbKOQgfXLjqu38m7F3fkVGGyZJAXH4u28C+UdXBFSTi7CDK5tPW+GSW2DC
b+oLargoAoxPeqdprnSqPcH7A4ZANC6/0UEOULUXiASAYQIN1e3ZJ310W1ptW8CdvRjVyzsK/hIz
VY6v0N7f9UtNtPL87itSrcHrpNmt3mJovg/ZJdxMeXT7piFlzECXJxLrlS2cZ7AF/Qx0QwzS5OTy
O6e5474tVVE6S1aEXaMa7vbCn3ltkbBibZEb0s1WCPI4kW68DKKAjGc1ex5Qe5tq8hH4w3nWpldW
/1xMz5tFXhUTdtVWZDzdmENam6wNs/FeI1qqDmFiOqxkr+CcLDsLihIBHT7WhR8pRxT6oW4BBt7I
/6lnJCLjXTFPwGmgZvHFLOznTy/szynpjUzQ8BpNsx8Wv46eEVWB0Yhmv/jfrxK3RTRVDMhMLorV
DnWuOyVP6n3r+Ae6hVKH5siKkU8fbY3dWq90lGOsmsnWt5jWyE2CAisfBwOEoJPJxbRZfP1i+F6+
gqS+itXKtVF2GsGnKBDe1j6JMLIq9PKLuwHgEFyl5R53t6i6hVSuUyAIm+sZaQ81/BMb0GqeJjmx
JjQfhsC77NUNgxDnjewbhW3qsffWjyhq2zREtLW3x7TYe3Ambbk+uvusgfIPCrWvhFM2i1ZncdhD
01RYIxYRsW41yvaEoiDnOasg/5MF3W3bQPNs40B0P0yWs73J30IO6P/knFZj7g0BwV5ZrFucqO7Y
7MEej93PAwq+8QDqhoxCllov3dcMTbLdt9/KTgki4Re1tNDcjGSDWjMqQqxhu+1k/WwqUCKGHfu5
0CDr4nxzlHkD0Rc0BbVc2k72DH5oLSVvgHRxn4XZqSliwmlvwtHnRCGg9OfJ6ikGYkYuh4Iptdvt
3Rbim+ADT00r4E9TAKODPwVS3YyZlZOGsZdlyBmMkzWyhxruVTqsOnKbxDj3j2ogdGQu6QsSyGvN
agVl5qC3IPPq2LbuznnukjdpM2RbfY54lulEoQ+n2ruXHJ4Ya8OxQotO2tokPDoKs3VFxbEhsa75
ohZQR2g4Pew+iwXfLnGaBAaxv1CWtirdY3Tum+UR2x/eWL5LFa9T/PuCdeVw/cCVHgAKns0O09kI
mMnICEgHhndPYPww6leSPFEIlsuPJLBra7//zpOOnSR1wWmcsyPnctMpiluZmK/NYhJWOATx3M3a
gojkZRwz7yvpnJCoLYCjB6JMmSkqIz/z4NX9w6NahQ+0wiogR/M8dpC7SS81Vz90hOnY32QknlJ4
b7L+e6tA+K3WAVWQjux8eHKqpkD+S+UzE+POaRK18x+Iv88bIwFNSVhHD7e9LRuamONlSYA5oXKZ
2IxezX/qRg3MJLh2m6IkiG8ZKd0Q3xgcyEnHlcwv+4QZHBsmCJIo5I1bZrq9Vi5RZaohPQTr3IFI
eVahntkthWMk61tWBM6LUx4t+7KdwaKQq6Ghkk02MzVHvqxHL1bKLVbZhHq03WuyX/SThmKAacwF
9QSgB3UzuSYtZTINidX/02vpk5AVMqYwqUEPte/hR/WraihSi6kgRgrOFqs6jgalgef0POEflXmJ
rWVhbuwwpGiFBQ4SdRkmfV26AECjsFH5eddHI7okDpGvxqUvwrJ+4fm68OoJQUBTDUCnLba0YWhn
somp2VYSB60FY9cfl+kuqeH1SrvxqEhE7th7BTa/uEQWxON0fLztjeAUAlvGBX7IxrLWklv2VkE9
WCy3v/rxajiuynIDSMLnvgUZ5SQe6qmjDwBY+JTFPKuPJLV9n5JbKHiSa6dFuOTABVXOP1FOGG14
CfhJV3n/7zmzY454Z/veuz2IGYJaeAf169aQEohFYUDjcypEBCszaJbvtcqWyGf/C9XlrCEvY7b/
NLXTEgICPveCRuXwD3u7eFLjGjFxUraglV8/Vy7sn5jl+TLU0RZt0BgSduT/jrP5L5CdTg1fBtM+
q88+G+3a4ti5BLyJQHCk2hNnNE6o0a+HTmVVVwiR1nBsB3YUH3OLtXpT3RJi4c3ZVNgc/2QL3YJl
5g+tjw+XXF6VZNKMNavDnZHuBwxFa+RpUbpgAbcQ4risdbjoVn3TdDYkccCE12MhAwxOx8eXRiOm
7ouUFpIzsPHrx8WBtPFX/ehTqH4jxCExulyDv5qAizWVdcUSUPnFYY1K8y7ZcBKAhOuLSSy8aEmx
l4aJIfU5noSTT01wcqYRsyiYsIJzZwnAHqKFhewElJ3ngDLmLAAqMfHYC4a+Wu+W0RZ1qQEeLNTI
QqNqh2n6wruB5fvsCENnLupOozKxG8Jc/RKErfXV/0a1W7RkAlVWRRHGKQG8EHRf23aH2cvp0Tcr
FbEH1w1esQ4osLq7xEnDdBRRJomv7LcD9RZggEkB+W28dj9wwLVchSm5vN+RGW7VJrloQs2A1oc2
ZK+jnjep5IJQQAJwWgwuhz+aJnu2pUrYM0DUru30DO8N3Pvj0Zx0twEYJicsMrvXYFI4yVKrlTTP
z6OLhLiRhnSAORYr3LG/HfAj095ZN3ijXT9jvXezfyA3mbxH9chxz7VWtyUXsDS3Xm/1a/knq0kD
ZTVNEQqhHPp4IaYrIHGe9jrQA8p+11nJM/mHulYMmmQT4pt09XbrnMplw7TSpIWhw5XaUrSepkIM
e4s+1W3+/F7qBkt/ycti7DT/5SfA8LYXY3GIDxXgvAj7WhLFouwFqOtNhchmSSFf4zopANURreo0
omNa13xYiSChxU610WZW0yDoUHNO/vZLWI6K98ee/Hf/BqqdVCRHJBEwHOXlAf7vVj3yi4YZryns
lsIp0oRivog+qd5Cd0iHAQ30jJx32jViU+2oyaVB5aaKWXMIWW05fCszvm1bkUb6JrV821Meu4fm
c9YEQ2DrSl2fTwRj11g7rKFMFRSy0vCvWHWmXoq2dJF4MJwVKqSPfBotltwHOB8QuabnZUtX/jhT
qB+MvUgtajNJDJxGjzCY0aeEsTYwPyAUQxOt7U6yOiK86pryDxWr+5Qopv5hIiJre+Im0MM2kTaA
1L7u+Nn5kS3vWW8K4XOPZOlgS/XjKq5sQRrEqXiAqv5JiQauUs8GFHbbOr8nzNG6bS9m/DahYz8C
6KJanKEY4qS0tYXPra/a+q8e+bYEBILp+bJ6hGi4imUTKFz70eiWtoDxON/l3b137wlnfya6uVdF
h8e7+Ks8k4M6lw188yaeokukft/bK8Tx4s2pcywF0H2A48GTTZgeK0/Zd1Aee2ToQDf56Q5dV+sx
bWx5SsrdMOfF64Ifk42fbmXCjohSaL4dHYrhXXKXmEVVwGjDE5c9TIyOKC4wXkg6QFayKgW9r+6Y
GBcF5pUoxZ2koDz4BIN9cLikvK481ZfoQNs84zgNVIyohnVk6pc6NPsoEcTmRav6d8zK3AmCCoAx
/NgdsznygoXYyGCL9fRwtlZWRw74znBPHQhlWeSAwtr4F3en79aQ27W3b1R4T3+iAwl6MZunBwhM
Le1BIu1XN6S0eXKyuSQmZf8MNt3aumE9SAD1+dTdpC0eF0OqIuX0Ecr7NXnH+KLjK1rUQ/aC2R9P
5BoxNiOx/8maT/7IoYs+09kh4FehZr5YlHL90nzo1CHJorok1TkxgBwL9aguwJnl/i0XxfeTkTff
NcsMgUiZPmuNkuowwA+ChMl67a0Kh66EBqP0xVI5/5RPFp/RQ84K3I/E3qSroQJrrmrA1c0TJFi6
CNs7YSDGA+PRK++alGcrwGVJ6hsttKw8HogjtluWe4E+15ycR7Md9A/AXUaIYv06uGP0BwZKQH52
Bh58hGX6d4p3rY8+5KJMcEYmKJ/bBA/51DeQKuMtcQB3zAoU5QJ/W0hTJ8Yy0WidZXIG4n32IRXx
yaMeNWvfdwiAH4ljg6PAH9qL19bkyQPGjuprrzA5Sp56xkWS0I5b3ez4upgMTk07ixFXdwjkFfV5
U8TS0cdqC+S3iY8FmYZw/Ye4G582E2SPwt2XM8ANs/+V1KGV607phgffQCIJim9TFexjW7r0zqqF
1qDoGiDOIZXC/S63PvbIkcYGs03PdZfU2bEEOKU/B+2GD7zpAPbeDRrQ3SN5FtUBBY9LUap5VFa4
JGWu16pGkapM2M/L3qfsjBnoZcWp1K5Ji3xddhK79aR1Ho/5SLFjsIaM3s6HxxNCmk+8doxshbLf
fsvDoalz9ygD2yOATg4sqTIT3Q/CMowFuB8sWtZhhk/ctlnxkqJwmAV/w4qbSVe9bX9j04PWrhrd
GPJFlcOvCEa8pjpzuQKQYrVnoEgXgfkzgx1Gfk+CMXHQmL0lVeSrVRrwgoYbK8jtGVmdnsq6IbH0
6AbVCbiLqiozqblwE8RX18GobdOW3XrAFnmBgoi+TNHPgJvivRiUncpysb3sm+YrsfM3D3dKqPpX
il98vqFXMpx8ov9u9caTy9dr9rdOi13YPo/DrP2IRRna0AqTdE3sqrt4pSXAlPICPRd3oAWLBGTW
kTeiqe28fhO+aT786M7hPiiVxEtyGqaLEFWmS7ooRTQGzpk6cCYIeHybVYyCmDNLaXtvJdE1/adk
Hz6bG+J/CUrb3QrZAnRDG+n9pFjwRRMRwR9Z5P7EOLls4cj6dacETooqluSLdpxLiPi+9XJOdz3w
HAs7Yk2/VLXFI8ULGJ8sToLDp+F/QDd1HnoX9hRihlv6rNHJqe3yulG+7bnjda/ytLoIHJm/kzGK
gATNZJUmqX8/nkY7pWTw5UpEthcXTCI3auyz9h+PCgsPD+XgHpV0PEuCqrPEXlZtVb24ZnSbi6Mw
arcevMhuqIv6SS80XBoMDjd9eyhqlTC9RYrKKmz4PJ2YxuOoAq47CIyacCvzDO1hbr8y2nP3P4W5
RaiZkMe5PNxc33La7KZNIXaBPWnA4pr2icazPbFFzz5u3/kP32NypnnMI3bPkrPCm/2bP8cxh6pq
PMbM+Q/C++QUH6QxD9hUeKgFQa3K2RBifq+zouxpKgN5R/Hoy4VR9hKW1O/Z0+c2v08dHV+VeQXq
bkY+Urcie3E7uiyUQB2eoDKYuGu14TOwq3a4G06UabsNv47N/fN13Pb+IWJ6wOJlUjpNBaQGGtdk
Su7l8eo5XT6WTIE6K5InzZ4Wak1+wlhKhYBFdwu9UFl6R/auQY/P5AaEebuimIYgLPHpCgrtnMHe
ilAfdQBlZ1JYeKJN8RoGpEv9yIlCCBJZ82+4R5DRxwzfr0pmF0mmr5AldRqf4ZVUOCKOeKP3C3zj
iiOYlLTFyh4Ibj67t6mTBEWA6dNm58Og4nQjkYHku5xR5CF6Ta4ysXkyqFWbT6iOTzqWh6KOAZas
Iyg7hhuIowhYuMVdj63NzV1YBi5bXmp0pRI8ZJ3zTohk+tsWjIe6yW+WNo//pTJr/MBotOP0xHGW
bz7TvgHERa/BC036C2i3qBn76qkQeLqYEn5hFYGncG+Pylx78yRfQy9guj3f9kASyzhAwu0Bt+IS
VosZc+GBs5f8mEN/XlZ5VhY6dF2JH0OGiNvTNFHV9Gy9ET+agNIz/sJ36KgMSuVwYEPOObT9Z6GA
P7sw9FwTG0OI23ZgiCoIEVTPNEKHAP2qTiyhUNG69BXuRu6ceNR6abTZJPKZvzlsEoWZGVm5Soqw
gJLNx5IDxW+Zvr/qmg74cXKgHpIqo2y4Xhn73fLMuaagFcyOOZdUt2a0izylqHcodHs0B3uFmpPE
71qJHBk4evaqrLa05crqHmfoH4ReKV+KYcmNMsbPXe+neBc4l15gN8DsW9DYajvOVDsihT0swEyW
cBJBJwoXTy8eweLhenPGvDQV6qU0qoPSwSLlkL246MTcW7gCT1y9G3f2wL10rQ2AA4vsPQsQ+T5w
w/nVwQzxjdPBhBi2ZMGyfUSEf+Vqynyrj+YrqqntkC2SfbDGieUKp1wHkN8ZgbU4XGqtfkGKbOds
HB+O/fIWKVn3pn/wl6F4KgIhbJJbCvlwzCxKeri1kwR7C25BrKPn2k1peZrWoG78o2gSEXkvj8nw
Ue3+2WeVAwmliLLioXXI6x17xcTLfGw9ubYMfBb7QN9qq0fhTYZ3YeUcooh0GpydnIZ09bFXHvEC
DDf2wSpLaUGKlWvWyA3NSH/9pwl8dUWGC1vpTXYAxz0V7fJgWT12H6SB6PAgXJv5LZ9j6VvrIiIO
OL/ZpTLInv3y7Fhl40Ua9sqkXuU6k3iScr9nUpTKInWkGvbxRHHQqHamcZuOBETA8FeRBnU6z4WN
7eTUdNaNHpMsjg6cZzSDHXVV2Mb6C61M/zEMa2V25tUoFecvckSQ4gHVMz9C7ZsR20pruCEEBnW8
1rpidiqT1DF2Ga/k6CtVwxfVS2IkSMk+Gi7utugXP1roOFfwr5J1RvcwN6aEq1bA38qEvYnbkjhh
PzqjZ9nPodZDDQfBbor3qow3fSIu3cmKGUGKoN/OQvnx0yecfOmmwhjaYLMjju1yfwb0bkaHxs9F
226pP13xXRVnpHZ/WzJrarqBBbetXj2CS/OA1HicbU33ngywoJUmIJ3wKO3Z1qzHv1q6NxZfUP5P
0SmQK3xwvmpjX/EqlO9sc+kq5GVELjsc+jUwlVgzw0mjGz2ZWiqmDY3gVPCcVRHj8T5hEbmmjurg
KAtLGkYIW+PCTOcEKc9mCWp7yxmTrYF+9Fm3IqVgUjL4Zm10/ZehC2jhx7pzIhh6YqxbhtYhn/Wv
TpGygybgsRp+5i3+C7RA+C3q6RgCF2mhSDxeQYoNF+2rUO+dYNjuNJSyIjjEuEusgvONAgEXCuDV
pjpWL8sFfsExKqyrafG2RexOU57pO7q8oCPi6tVSq3dTnpAy7ftWJRUzN8CH7Nz1J/zdKGojvNLV
s3xrGYJ8PdfxOxHmc0ZcVCf+iLbjzuJ23k0SRxpWOxp0zk5l6TP5WIc7nOB6PugUO9E36oMKDNU+
PdvF0u/Crd0HPWaXHoUuhcQx2Hwq08mAvmuX7ZqARSSuSixJcUDAtJCLF9iMzRjkwnFph8QmE+Oe
Zr/rM9Qup4paaoAr4quNavG30DjsQoXo8aCXPCuslkx60iHz5IjVG5R2/95qhGZQLwOdB77z5ziR
OGMa/8UFJAmKoAJ97wV4s0ibJUvl5yM2faFGtJSjq3qQcR9ofK4LL/+cMb4fPjHPxKDwPwoy5hZQ
sQpGO5d/plps271w7AuDa9fGE3F9JCpHsoQ2gAX0XaGm9ZeciB0sFLGtvDl4OYKUjlJJYaNurBad
vSyadW5Qus3VZwDfZsYHtFUGlkX4opn21IdYWHIhKrqx+H61p8B00+3QmXmxt1xD8KGF7dx6RAVk
fALopYnrhzZ1rPPQQlRO7af8SC/x6D6UFhvTchPCtrw7TG1M2c0Juw4H1Og+foH42/+1ISDaQ4xg
aiSOpn0gwVAj6sil5g12+GnN/B2u5/+rYUm3/+DUkjEgfqJsIY5JwefMIrv3HtRwJiNp7xubsOiY
Hfc6BcrCpaOB2y/wbpVkgfTB77nss33kpsoThdLojkrhaYi67pZaffFoElPWkXuEbuaBs38uy/Ki
r75ym0PyQvtA/fNnc2L5+mkqrocX55v7X+PigglJFjCLUsSifqc5Adgv2/xEGSm5ppkeEe9Kom+M
kdEbrr1PHbdiLXv1bAHhw0odKKci0JW99SQEbd+r6rHGbGKpuW9oNDQ9vlyCBGw12HwL+rcTrbxn
Hf07p/fpL9zpEyilH8znyfjBWaimwUoDx8QME1Mh0mmV/0e+XEyTYLZPeSZk2GMYRuMvhRJt/Duq
es3UOmORFDj6J8xFRd2J+5O1U1m6RGjKFHYHhcOP7iJcxpn4IaMQPjNsodXfEctGZqXxI7tnKy/M
h6ZMa8uEfoFXLngjSnRnslfrNcXE6Ps2ga9ghcrtr+yS0k5kU1+K01zFeqfONARlEuwx7/azLYrJ
g9lQnYqbf9Yi+4rbcM0p8ZgL7doBjK8RFOVhsS8SdAFQmslhtf5J/xA24I5BDYDIYCxwlccd1R3+
ExnkyAPkToq3UIVsQw9MiHtgrXCbGkeavfZSYm5kLF4oBJV6eUwKMYWBWkdoDo9TxV4qI6fhldUk
K5xsJKQYx+v028m6nktOudEN7TlumjMECJv7yr7tf2w+1oOXfxMVo1txiGvCe8xu9rqaunuTMAaT
6AVvJOmyojd1n43NIX5UxWiQdVxG+vSykJIsYgnB4VUcGxZYMHAeKI7Uy9rFt1v2YqIksiBQj+iK
dBZt7VkVn6Hnf3ZW2AAcIA6TN/tFh2vkouRO5bs4vjqTaT2zhslXwAW9HX9H22GhlFNvV6kEI/Wv
8gg4qHDChT4X/gusV1j89Fjsf0Evzx/h2z1+AcBwYBrtt3LRD9dUKz+c6WJJQj6wk5JGHzEiVAIh
NNlfX8o3jSPfhBJOKaaxSK2vM/Rmibj46yPQnnJl01/Gfu5gPx03C1q9iQ8HW0rKrJgs1UsSLF7A
dCPsY3wzfVzO5Z6rqzuIhKg77LjQldIaso1X3G+r5gpr8PnELFhWh1K+RnSA/xIRDA9FGKwBg1X0
H33NxqxXjFVNUNMkMl7mnetzz+8DonzWllsQHg+rtGLvZLFD92uxuCLdzX3ikGvdUFmr+fTM7v1Q
ULiM7EmYdx1qpssSaVvR4R1fRePBvN6yWUQrZTcyQ6F0FJEEpklexIW7y2P2FeUyVsgmcTadyt5x
TfDsGZY34a/4PdrB1K1lzgJJ+RKUV3jyg6BtYUYv3Yryv0OhHTWClBCk40CX8l4/wwqxozvBye2P
BSfcxvdKWCsvKQ5IWZR8R91sApb+ZpWcqiSRr8JIcV3bo/9jC2y+88MbtNaMTM8ihdz01A7Eyzjw
2a/5V4GCudtoMzgcTJVv8owkuf7LT/YGAxv6whxKUZ3CwKM2vRNB62qx42e3RkXEfXqnZdNbJD0z
HdCDKT0sKPV+i1gXXlA94WoYiT8bayVuwVLNG5+pTRNOeLCMc9Q5OfA5KFeoretM14L2kq+i2GL3
Bpr1MCrIpBP42916LBHqJeqCyQMUbERH8nrKC3yPakaOc8cpxygSdm3d8gHZXY8Dganuo9x8IRRB
r3c4VcWiNvejESLEe1OGVheXrnRAyjuBcH+0N5Q5Iyh3dYhaqD1EZrf/zJsYNhIMm/ZAGu7D7hlX
zIr4qUrXdjxLt6IEIkvCjKuA3kFJe3TESTQjrsYlPb5d76CTJWo3U2qZ2J6zbDPNM5PRyiuQt5mW
J53lbDFxlr97vgyIsQL8J38RDQE+SaS6aZ7gMYnNYjNsDzIRCtGZG4S9ueyimh2lMN4VZOT8og10
7I/oLhxH+682VV/BX8TrXXcGYIgLQtvVsof5t3cQGstgTm45b6FlFoElMNlTNUB/h+rsLe99Vu2B
DCxfYiNe1abfC5gQQ80h6jZapnUgGe2JF/0ib3k+VaY6DrVr1VP78Xg0fTYVu93xs6j6v4Q9KyLs
JytPQEHpSY2jWggiitBnPpiJUGhfQMyKJOUEZpsuihANjN6Hx9WtymF1pZ4KAQbg1VCm8Apz7DHm
nPb5wWPlmymDidLYfQi5txVEMa/uTRo3i6MSmC5UinJff7ICiGh0vv4MbUsaVY4NmLJuBzIbCt4C
5J91K8Px8PtkHZolHpYryQ0uh+5/Ut7r/wMZ6PpFFrlDxGqn5QxDvRLVrFa9vrC78KpfzPPKtGet
8xkQ4h21VyjaSea2EYuNCFzLtCf7ZdsL36tlTsOJcx6l8nzFkbfQphC6iPndbHLekBBLhtBPm1vE
MgseOS+ffAzKVpOig7HjWef+PVRGy04xrV5qtsNrfuUzFdm5Ewz6OAy2j3OxtmArlKAyVx0V4s0e
N7+uD5+lue2PQtZkAUbAwlAtU+rFQ1wiifUhNF+XPKrno+iBirnEYlRzYwJ0HFLZMb3xHItolMvs
c/kKAMT7dhmchwnN/WyzUVArfQ5XZ6Eezowg2gvXnyay65RkSaEohe82P5RQ+meHw3ow4k1TR3Lj
5Gj4BZLjblg8woomTDf0UUWhW6XC8UH6NM2mKsmoLXRO7hfczUEqz6ux+Q21em8EpiKtfdCEpkJv
2WA7qlmh0rCfWucnHzTiBs0wUr4MK7qOnr87Cz9HDo0gNdLtgjgOvTVwkyDFznFbshKkZzWQet81
5cTHatTHrgQxM0xmev9WNaVuHv6/ynJFYNhRMX4bitbyx65F6O5ks3giNpO5ycugGNQYCUnB7Ji0
1a0EPi8eCJiOw1v8pcXcQrn9F21PAHjrQwnsh5jo69/FV63IsdfMS0sgR9dn0ZBPmnOo0O/fEUWY
jiI96qDEKtQNnZyMp494siNBv5ak1M2b9UqQlWoggwHYFNJpqsAomLxGGp54gcbQ6kJ8nkaYrsFM
8J1PGlBx9vbjJvTJtPp/66yPHofIdqQgsVi2SOi4pql6FFuOgGZcJdEryXI5f/HoCDVD+Uqhq+E9
+4CtmyFv8vUK+D5gVK2umAari4WYIiblPfvummgUmFENzvTCCp6qOxeAyPMPR9uIMzFpEgizxAue
b4B5p4wuLJj0UzHdXAMn1rJQi7mJmYRaX+rex+DSQ9PtLCrGL1Qeomq/IWQn9vzDFyxh7pQ95F1Z
SmCKI7lIOdveO+0MXQKFz3KCgKwFXfgLoHCy923n1QaVex60ByrLXk4/s9ZG0P53SBfVylKM3eAJ
Ih9gJopmtspm5EUzCfLrk/WyxHvtEsuPh/VcoKvD7AjpmSKcLQHIoUPeQj9iZafyK97TDIvALLRF
8XbdAunHx17VRAZla9RJ+UUWOD7X/aTX6dYuNcrBgRzuvCfFZNvfbYhNFPsSHMNUAg0D6FZFxMkK
3Ojxi+epkGc8WEMD6FmpWeNvfP4CKnghWpLCvZvhhNgCj65n+ghrOrgBaQl51mSDd+q/F0z1S+np
V08/OxI/f9GouTR1d2uKtsC3B10UOfey+SGxV87FXyp6alijky/lCw6KQbRqB/viUZfEKA+/7xXj
tGL20zLnudpJ2f8XVOkyc6CMueHM+GScm9W9ImnmbIGNntrCRgSchY0YKlRCATseF2IY5P5gktDZ
tN7k1AHCLNgVZlkPX0a4tEet4m4FxYaGi55B5n2n2tTKzT5nmnF2gYM0ve5JL4C8evvxRpsfKZc6
gUD9aELiuUhjV+tm4HNJjHijDPCAzGDO/YKCNYh3MzZFOfDUsWviiniBLmGjuCYD7cLdOYLyz9NE
2fHw6VRyK7JMJ6sdV1b9KM7Vlg0y/UMuUnHCfxSvYojSn/BA/9Hl71jijjbTxub5pB4dvsnS+KM3
uSxEHugp60LG7Wt6aaB/gL9KAiLgJ7OYNaagzm5XH3rb2Y+YH2JgE/F0bzAkny3Uh5ZETjTSiip6
+oNNVMU+/hg9NrFPyW40ti+vgl62nq78Ee6b5f2vjcch/aFBwbovv5uSiKvDW/o2VotKtk281+64
VKigAweR8y7gHiaGSL6iA4CsswVd8ulOAI7oTfIBGBYZBLC3dflx4Dofv7ZCu8u9VYOC4ZCXZZnC
fL8gCR5Bgmq+yTH32H6wkdbusYDzs3x9R4GHczj/3k2DCZ9eqhIxMkOe7PUuXOShCbz5ipt6WgMn
fQYAemvfd3rRlXaWGFneL8vz2SaW/4hTsmBB865gseS9yIeVvBLcvhLdk8BFeuFAV9QNaxy6Y7zF
pcOeDmtCTYhoRywu45PXKKlX512eSTb2kJdI1PeLOLQfhAA/JavWqgv3mRfwqPDGSE6R6KRYPckT
+ieI1NJqZ8APHl8Zd/egGYP/DWUGHgnVTXIF/JEu5TTD/yOfLERehrwFfCCzpPx1ZWduaPM0hIGC
M4Bxezc9oMRD7DKKElpJ96GTu++zHIzmf6x5yaf0UQZGlO5cTwXbcec05ZHXGX8igfpTJPWicfNw
KNmJw8RwabskjEcb4u1EVWuGN6J9eNqQ1OtXCeC/nFcAT8n26x4KGMGz6ex0JgPExzvqrpcxyJld
kkP5tcmcFFvFUzlzE9gTFYohBFczwMxDFjdL4RVzl7WUCbHU1VQKcqUGxKLoIegAlcyv4K+0KgiU
En790Dqbxyn4OCaoIZuIgQRuN3Jgq9nJ5e9kQF7HiSceofGgRhk1peUpl1Bg9ggic6MjhRyKWr6E
AvCVL5LNFtTJFrhrzR8c5aXuC/BNrkfQCJCjq12CLT9HfIja+5jdUDmqFdsnk1ZWjVOVyV/sHNPJ
iNATbHMa8zaXV4Y0aM6ALsybyluKhGSBFdKwOSUi6jqNqQFzKsvQmwTXSdurguFll2YyfEcwWGf9
loEghuJEXw/ocW7icdXEHpZeBIKU5YxSG+XqMRLF7afq0JJddRXF+rbqAy1M+oZjsuayiGRb6H6q
tlxn2GbXMQlJOh5O3DRj3T41PATEZ02MenPXrnUB2PxZrXX2fiFNeqLEep1xDaxrCt79repZEa+4
zvvmPdI5B09beJZ3/Js/2i1bxKevaHuq1wJHXrO1dskBBrcGiu6ZniXf0VV1PRQBZxNUz7OdXXRV
u8qE1aqarL3q218bvoqFEmoA7v1J+xRm32TqE7TTFr40MHez2Me1mCVlA20iveZ078X+KPk5u3G0
ndfAA46yuQmx55KAPCxJNbmY0fOAHw9EKl3PHYeUAm9/XarR+D0VioMtLwyEAGaOCIS/V1ZTiM5T
+7LWpe0YGriPg8Ssr5yJneKdUK1Jcq0/udASMrrKHhrIwaw8MH9Y6D6Q8G/8qIqLFrlWmSJCtYsm
15GO9LTUqqnpox0r/QT59DIKC+K8fr6M6KXm9VjmnYlDiLwU/J31bzQut4cAlH4btmmSx1IolkOn
i7fGWY0FtRNrY6DPzf9pBhY42SgjYeQtklTKcWNxgnejv6cAfqUPHUpP96NIEf/dQQKu8ra6gngs
nBcoRZhmQoZAyn3afPrldznkrPZ6u+r86AzQ+YwQPwSfEmAfpEuWTugLDzDHKlCygBYfOsCExFKf
ofVA8UiIudjHQc2qXHnzmUqng7ENyBtxp7QgLoQuu2JtXspFGDyEyYCgOO26BOarRb7SbnVv99hZ
May8/QsAcynZ9eNcwGdt3vQ7Yjns1WPyKs9QO+usRaLTMSu1vinw87Sb/OxrhnB+18qBKfkVKmyy
dBuc3nGfnJlsGyzCIjEX1OA7se0winchWbU06mJo2U01dcUg+TWBvD2GDji6he/OyOakxR6ZyGgK
FgLj9Rq1BB3DNPAyk/sXb8TMV1z9uQcYpayfR+OVhw95/VCF9syVlEtm98kZ7mEl2gpqi00HujMG
cGxxDs6Px/9Do1IrEqrl+iMXxdR0uJKyUe+w2xB/tfWv/FssPGrrDHvcS8p6r/UM66nJpOcJTUvc
OS8GDThTurCo4EBsqgz5fUj9ul/D8xuGqDh6gXyGDIew521lD2VBstCjUP5SqfiDNbYJcC7KZFWK
+ffKW1x2Nm6QWGHPa1cm3BmuDnqS8u1jph3YfBW3ZKECOuO0dn5NX2mdLi6rINYsxlFOD4q3v6Ri
kk4oKXpcZW62GsNDuRoAQf+/dQVYvhmbQzts/yFeYY9feufhOZ9/J//hwrL2Z8Sv0hy5+EriiKsB
nBeY9BOzR0g8sRaqSNlws9rnv8RD9N8KnKr8aN3GkW+jUslyEyQXFuA6SooeafjkpxX4yWL1caKe
ADxxYCyBZod9vxYrEl0pOovgj4Eq8tugvAIyZ4nLQ0gDH023EAUORLlInZP9yxYMSomI39Vz0Pcf
Wz8qk6qF6V24mg9+ugF5TuJktBOz2xPMabb8VYia0NmHb5fGSFm9DsuWXxZ69VrXXLjjwoNMGexu
7HpOh1Y+XAqbRBOoVrU2Cvh+MampDuGkhOnPXw1+S4hFlNTSYMLND1iBppp58tnmCDXXUcPg3XMj
vwUA50sfWc9uWLfKx5JTHKPVHT6Gj2ZcwCgB2Dn7Pb/Iyv25mb7qlMiSCYJR6DN5r2wamkOUrd2O
+MLzhBuMLMOaoW+KRXXzby15kOJHc/+/O6M+/VxGiUSMd2dofcX+QmgA3M6mDrjEtslW8CVbmdH8
a+W9AsKV5V12cabQzd3p5xn/0w7Rj7Cx8pJdMkKMlu4Iq0VXbwCQhF4DfFI5ssdUpRt1s3KVfoyc
FIg7gUW870zva8MaCNwP1xHYnm5QMkW88iw/zaf/l/jZ34VoXBTt9baNbbScrVF+Hjv2nV2G7xp1
MSb4aMj654Mi8cnDCCmSxaHQ/qqDr3U/GplxJIcde8iKAwrkMxW7P7ZkO+OyeF0H4SK/gnBNqygu
pgTE8rAQnb+OeM0KZf696eG9pbRSE3RaiYiLlsKd25WpxF1/f3MWo4HMJmEtJWKN+ObU7LrQnhml
ig76A4wCPEO3nmhh8plPkjsD5vXx96UArrcb0TVLujYZy4yBVsxqeUYQYXFQHEpsVAuRa+I47drW
ujxmBrxH0l/RM+05OlT1Wd7okYaT4PNRpIoYl3rj6Wf0urmxFStwdgW+tCUEo7L2EfwqmtZs70Qq
c9R0PaaDBJ8suyDsJ/zVW2OntFjxaEt3sSBTHqy74PnOQz+MP017/4wR2aQisXbVNZ4zNLOeVsB7
lOWi1fJRRFAfgB0bz51O65DTViTRSJDqicZBadrBGY+VemmJrZUcoEO6JfVZQwx0diCflsEcUDik
kvwZvN19TJyecx/dpfsu8HxK4WRvvdCAmNOOXStv+nUue4lkTJ8jdA8eM2Jgv8U4jhcMG9ENi9n/
YJ/Gzaz1URmQxZqEFl0qjhL1238wTmllqoXgK3+vruuglJjHTcWNNfwVxXPjriLq/bcM+9y+tzXH
bJiZeUyup2TWqeGxMIQKfpU92n7V4pLKNTqwA9NR5U4rmvrv+ehYHCtl7msiuginH1OLrD8NSW1G
kwZwVlkUxGbcwcC2kHVqDwhiyftIjzBmSuCcEugv0PAzIAHVKvqKJqY9QCKMMBTwzJqpnh7CTY/o
IxJ0T2wNrNDWF2U7bQoE1J/C3KOlQsmVWt5RSgTTtb9uRLyrXsfb+rY0qykUNDjO15vkZNDJWJo2
vSWgukNXR6+HDWYV8JGL3O9JpDDFXQQAypdDmxGhyZzDy9wj3DZZhSVA2qvrtbpc041pIXpw6PPb
aYIofWStAAFlp89Tq1bmwQnpEnEy+PYMXY/1ViWZuz+vMNV6GFX+sbGE5ePr/45wILEao9dow1ke
/Ae9Dsk47WgmF721h+QjSyCe6UhuBA3v5DscaTnU4OII13RIO1H6VdN8zS3FQBtlSgRdQ/rDen87
J3ORMKj0YzQaCvqfVWZyPsxc7xZasOM8KxAVmmM15ak9OqNn8XR8/KfOhmqay2kz2EAH+E7VUBLg
VFGoZWP+Bey4cVyIXOVhLcPT8ck4e6UBteYqG7GY7f+Uz03NdgJH+nZxBAJ9tEFtO7hyqbIXM7yJ
PNKPkbP6nHr/ktj8KMo4FM11WwT6f5CdL8MA9MYSpmr8+CioR6tdhRN7LEPozPePEmvnck4Gst7r
J/Qu4s9BRDZY7U21UUbv1OCLTZ/Ra4JS8japdMUWhh7JvVs9M78A0qFOw2iEE32M8mrwjtdhhE0K
KQm47VnFpDuZoalIyIt0mpAQDs36pxWkKLDINTNLmYf9YIk8YBc+1XEiog1dMqIwRobtXLZy2cQP
2/onrS5vRPtM2Tj8kMnQl3s41CE0JkfoRk8BBmGUie2gV23HfvDG3snENZJOWEfxHwFKx2Fd7Jcm
zn5LfVvEew6xuxVLL3mAlViHRp3oy6G7SY0YDLhlGUyuzOQm0hdAKh3o25Y2yTGB9asxbdmaBUq2
3bUEh+buxNH5nQUV7dbfBseD+SMrTJFxFq06SEIo5M6gHCMuUpZ6ssTysTykNWAiCl5Q33C6QRms
UjzY8ooPJEmAi8Dfai0JkTGMepXQDvCWb7e426yEUYsOAU+24MG5bCZdygV4uq2xOS9lZmvnFeKn
+ubV8f+ZBGZFsMUWkezw97sUqOdlJ5uB19VMrzHCXlnls4NNm458Vt0CgnOnPvbHj7v82DPYlDzl
CATNuUEO+o/iTmmNu6jwt0RYA+gxPMdrDtmZ44EMBAJq5l9/8j+GSFH6cM9xwIqNNPuU1qGq3X6T
ZGx16sbprhZtmdqs9g6QD5JWx3Amyj+Am+zkUim2E9LVjTyKqXsxD6/VAfliDxI/d5zmIqH+p0HZ
33OaXEGy38ZBTlUXc6x6lpc1iSCMZeNYzomdh9nwVJQ59ArFmRSVMJxSTwAn6Zay83SLeDRvnMCP
iUT+GDxjr1dRps8lV4AGxfq+NxT3xNHXjDwmZPFezybt+z2TFSYtrEJT2AO7DyX5adf7lcAGXpvm
AujVaU+pOJdo6YZmKYNxZIKIRPqHoiL3e+/smjAuMzCI7eXFqlGtMVI/nA3XTGh0GTvoEgqULmT8
cCumO1JgvECWjhdI1Tw6ttjHEdMgigoEu/5d/dsDje8Gj/nSFLqIMtBtxtro8iXBllJk1Pg1df5B
cocp3nVif+4IxUpUTKGoUWBybfwRz+iOFjZVngwoHdxg9Jrizb45OgB0eKRTxOKiSywHtP1lTIEe
Pgd/kxIdAq/O+fBxUcILeWFVzvBR4lFmEdwgjAelRi5AIZGoG2JkTq/PKHd7sEkfNRtL3YtE6wnX
YHVCg+x5L509kDxtr2KlTJiCghQNpzcD37utw3neQ+PcleHoQt8Mm3LCJozkW0uKsoLzr5QgIy55
dIoiudROJnCmPPBe+PvhakjniItneagtkkcyqCPpFR/eOZksy4yZk2YxRjjANaYYu/OHy0htqL0Q
qGhm+VwADFuFG88TYOE4CFaplR/LNR1WK/WAnu8Qe7J4HOIxlJZ0fBFNI2z8pe44H6yWE4/cCPE0
GG/7AVyVAAwGefoqAhs4xo+HrYnx2XPvOyYo3hHGpTgE/823vBQSkw5kbTqdNJDPvi3m7F5IlCGq
ctu9wILFutAG4CFTWFKw4b85QL167twxVsJYS7tToseizy/asY4tGir1YeTkruFa+hzDF6WVIoiT
/GWgZ2piHt7M+OLryvWp1bepAt1/93Cs7LSS61/CBGHrdWixrAQsoFUKp0RaTYA1uciekWLF1ZZh
cRUpCRlmjuKFd1IfzUwhXEebFOM2PYeX7S81ia5UQXrj81jPHJ4WVNc8u1LdvAs00UaLQhQRmjh5
YYDPcUqAyBFeIubKZgKcIetr/IX/AqXiWS1MxUoTUQ2m1wmAF+vdgTeNXPnrexFLjrRzJVkwXQ7Z
XWBBznl3QNLEwYITyWdEPksYqwgFAGCtZOv1gUU7CZ8dKnE+pgiyMQSrAdKZuuyD+M6esaBQZKna
B6vS2Xh/Xzuyxt7PaHOjPNHKgM6DVyBtMQPKIm0JflOcsXmgsIiJiGFxFPd7442AFZdjj+pHOKTG
jBp1VHw2HvZL4w6ffbufgWOq7n5jI56V4SrrchuSQbmu53+Srm1dcJ0m65vYn2LLqxL+HBQf/CFz
fiQhXqUFR8sULLLClfkb9l+GIBHys7FkRezk6PPIDSK/5KUxXsGhN2ZTNLnp3d+LwjOiCOVQ3+pS
J0lPIr7nFdNM7XIOyl7j67G7Vs0X/q0V9uFjNMZh8IZ35L6s4Ece2DBXSLP2IPMH3tQPFjEe3y/a
lRu/A3v0XNgM7KTt2zmoOFzGwCt1XhZMY4oEFV/vRon2TSfrb2r4opVtwntp+wRVbmSsdCXDKODs
Vf1i0HOqfhm9FOqpW+XQ2x/NffOYEzP40RvuAZhT//ofLf2zX8xnQZwWMoNeYEs6rknxIzViowX/
ExnBkmPLzzjcOTfHLsadT8hMzOiCFblvU6Ex+kZCQWEHGiyCjhRmkXNuu2mNZ1Ljgjqkjq3fa4ha
U3MSxfMJhZmzLDk7gaZVM4FJ6clYEyy6AxZNyr9Rofahy6Oa4IPnsniARyJcYleCE0hWohFoVcW5
2bP7i2d3Wq3DwJX31IJdJllLEdm9WqsiuV4uRmq0i9nYEJpZE/k8d+BSUOssRU9VR4OYZDMuXt9p
GX/U8YlZBjZVmuXGwp+zcnK68MoWb0fhtKc3WU7HMn6HDsPfvuO2HI0Vx9DcuYv/AOK6NwTPcVfF
/y79V5ZDyLKw99o32/OdVlBl4LZrUtBCPbtZLoJzrvMRNFEtnatqsKrIKHgI5nyYGyW3OeNs7ES+
SnE6vO7jeBIuXkMeG40D9RzfEo9mchRsL50Mump3rbr07XpVHWN9f1CPlZzl38PNY1A0Wr1fj/FS
SSSJp69Ix4RGnHzDFSitAyC1pqMrqDWFO4UfStY20XxMpEIbGTWNUM1BOEiJlvaPUfbzKSrFah6p
KxLni409cvNPmnSiQKuw2YIq7s6sRjApJJ+DpFUqg/vAG+T9K3YcpWg0ogdPY0hAq4Tmzh4nR03i
UuDinumqCwL8ybzTEbTYGza4DYpFgnWXZvF/UmJmjWHB6IqkPcIPdBoUrm0TmOlll2IIjDYOr7wi
E62rjTg08gakvVShpEUs6hwPq43PXY8t+/M5RC09ovyN8QKRUSLCVwZXFS4Mnc3kDAqeQzvwvPBY
lkoOW40PGfPkmB/X0yihvhRLppOwonHJrXevhXATjai6D/ZBE7YLdo4ELdKx4+LRpCiWlKvhTPFP
QmjfZcSKek0SNwDxwreATwNxd6yvf62KWqk7TXrESAp8xsK9SP0b1iZU7FIXouUx7pTxjRs8LfM9
p2l9kF8r15eH3ulN0AHcM5ayM/uLpFEiT4wpRW1+zozfCI8qtSi3tZ44jJRhZgrLEeR7Y5O5NgIl
4VVZ3BGr5lejOr21jjnlc2+CxSB0rrYidFwJfUcUljCrrYqdiEDkX4Pgso+f9POIAvFVUZZ6N5+q
f/0TW+TBT7vE0j+HCziZC3LUGYEKzZrKMRJTjdx18s7kB5+mok3mKU44wzWaR3fNYsmocvASPLXo
+JibGfdFp2mQ/eaP3DO1mO1IPcOWFuR1ROO33gU0pbReNk6rZIZ8sazd+uhcUfKuVCsvpK7MS9R4
k7siDGS2vTTkhItwyIf3OGSUdoeDT3YX6xf/XGb/V2uu+53hz3XIFnILWS4puh2X+41i1wg2XTFo
5xgKmzUebEnz3m3bKeyvJnFGWgTJMbvkGZIBjuFNvarRO/bn8JseUBatwWZIOZWPNzNO94dj5C7p
YQ9QpjRr4DtDjuMUe020TDXaG/UEbBu6v8jFw04PQLWkyq7FJdxSFPG7ntXnru2tOPS1d9ianeGf
qI+3t3UeJhMaqiC+2oQgDTV57bi9JTgMZRIPhp8VlnFSep8vHNKBEXaKaHYSbw+l/tnmnUnd2dfY
FvdicStxOPpGM5+TFwPOr6VKKw4n19G4UpYnJWfECMpydf85Ds2OSEtSmu+QOoZypztiIx/39FFU
Ey4Qd4luioBSXQtSFsNwuZMAI2L41s1+Fvw5a+9y9rpwX6ckMmgeOd5DC3yoUjLiKcIY/QhJJGa4
R3l568WJjx74YP64e8RABroeXK+CBpbxS1PwLiIlWArV/rBOzdoqoUwidwaOR8IOW/gsHojackav
WfDXJw4y6PGQ1bAL5lcUMovYrNqf8TpfuNc4lMB19l+tEUMPFJk6IZWVOrN9vkxHyN45yZhlb+Wd
emD4M++QwZhqDDKNBoau4guBVsV8m+xYSaxqdJsY0lqhd9sySFmmDbQYFmZFgPVoH6k+YBjP2kVF
qzPwbXzKdoAp9TzzYkkDgmtn4q4dz01njpNSWCoj4sH2dxa/im3tBryyyUqRwXsA/UBwOyK0d0H1
4Qm/w2c2p6y2qjorRYFG+ARcb7LtaddjwwBc4uGvvVks+x4OJXTdnnFfglxXgX+NgLzr6YqC0Lvr
lDRvqbSkhZK1IKM9eFFMrDnZ8bUHek+c2nNTAXWeKSPPJ4n7nabuuqRyk98MXjWcIgxeJGkE0uWt
qACqQbLcz0By4L9dV7c1V/hq+NdzXZPpfh9hwg7SVy2lUSLRS2dHIJIOro5QncXqtPqyNSW05iRG
midQQ9za8GY8R479qckV7yn3B/5q2n/PXtNC4jU8hka31U1stv/4/8ucRUvPwxVyjjaKzxKIdtAM
c1h8HwbxyoJzjrZceZ8rkQwl9DLeejxIyeK/K2HwW007Jxp8dfLubh597EuOGRgUNhtqF4B9TKMX
Y50QCLwANTZV4rS+X26gFgEpkvoH6Ih68+46nQgwmVlMNz3m/yskKMNnD9ZLv/XoUM712hH8vlYK
3whlveaBYGC5lYHeD3a+Sz1HsnAT6C/o9WObJY1kSGWJOJy/lMoWEYs0KTloN4lpCqgId2qjeyXQ
zTCrt93JUPw0BRykC+RrnhaaXvxyOkKgqTkFt9bkUai855xVHMst8iHTLOONFdCcOa08DIDRlL0Q
WiOUanhM1VaeNQD2ZgKkpu2CFbc7bx5owBvo+VjhYwLUt1UouDqbu43H8xAwemSaKJ6/25fr2UF6
PKdM8Hjd128vRidxWROQe1Pw2IqE/gIjWTWEATuIhoGtfGsILRg2sb3WWnmQ1oEpE0kq7eq/GDSg
GS50hbgRRBPp2iSk+5q3+tSCr3sMNMUiZAc6EOgpJ4u8aX0jQZw5YZ0GpnDv6YzC8lKtP57nLzLf
t9W96CQznIE9nVV1Pnwj7aV/YIYuXSCHO+xhAC0y3wtHL+TLIK9HHRMc4xA0OLTnKAEUVv3ReGkq
lqy+L0oadugVJOu5kPNbdb+gl3GEt+s7urWSoVCbaGkVXyU+udbPlulKU29opVdW4MlN7Sn9F/0b
S+LE676WYwy3FXtSYwH2UV5L1GNjoEUVbYTWCHWX5ZRI9/ao+F24GJIkzex+Nzkp9HgQlviSiMhZ
EFdU8bUEmnf1xWva2+l0AbQDkoP2fbgwZuSB3WnN0cNrnGhd2hetNE2CG+lUwd4z5OqZqSuPyikD
jjzkxe/WqX+YC5Zm02duZdjDPezvR9deDEt5ZLWXQiVz/S/BS3sm/C0uGlunbh4IXxQcuwlhqbGJ
I1YtaJzZKE8GR/wEb1gDw0PbHrOQJeDPyGuNJaEJnohry0oFXB2c8kFsFOj880dJPoT+dUsQI623
vdyQVidLc4Wnex+A58B9/VU6zPV/TDdwidyjjZm1kVWCqnfYVLIQm+WzA4Vpu9trCexXFu0yLMlP
I9BC/qrxjBKp6MuQoxUpSiaAq76b7KvARf64zotfRZFTQlf5z6JKDg9ePI7C1xs2YBUdJb3Q3hIX
GNrVEnD1B41W87sJp7rZbGwHDZ04LhVKES/wrLLdEbvhWVtuIyGWohEdJPOV+doWp+w4o/z1vnxx
10aqW2e5pPltA82+PcZPCmzgNUy9LssAeMnnfUtNVGWVUgm8gw1i/qS+n2wmaRjSoepyV4rOjG40
gwMrhtuD9591F8qO0FZo2ExJTPvxCiP4wAmkOi7C03SprYjU9bu8SvA4u1t6eoZIVgSGUP8rOJdm
jNxaNIRJgjgzj/EmSnc1//5nZACjfwNVvQtQLZoeQapsK2ZaBHAoNCqNrZTTcFKVYsZAMD9lPXEL
XDkGJEzXCENu7/fPvw6sK8XqFmyqLohB2UL7bvDbdVwCd+8rlOh8OrtVXPC+KA3eIuMUB9lahzYb
lnaIHiatUutUSj5IdkZ6C1WtyRnSpOodrowbhOuDFKhoTIvVkw7GcOjZQtfWBYzmRpvslPROOh3R
Qs1/mZJISr4xu/vigcHVuJHXUByTi+GZ5f8e4+sXqizK1QmYXMzIx+oB//xV0luFfnU/a3/l56Dk
rUXqEULcvHJlEfNQUGGw5MQfkg7eKD+bXzRbfz5bq7WUUlM70c5DHDHEssx8A2gB3EAPdmg86RN0
TKPDIuL9zq3Ns50w8v5QbYOaNmZDrLrBDh3KPhdZib4vzan3n4fjtJlfV9y/x6YdIyQRs72I6ub/
4Ox0vAMMo6BNlyj5HKbY1i6zNzo+m1HPTVwJqpN0YjePMMHYqP4Gfn8ORjSqnBn78LYMpgZd9LZG
0gqEie8DdeyLG2vjrLerliAcJP+FVuKBTVuZJ1TN7NF9GOhS+vQg56UkES5I8qNDmmI1Sh/yZU74
LM++k9K6smcodr/caichbZTXp6LkmY69IXvaIEZGhJEUZvrxM+HU3umzwXUxAQmA1kxpFmdOV+5+
n0wyrYIYFe4EhzMgTYe9S7lLove4+MVEYL7YcTSPmIwl89/zsCEyPL2qvhwWRCgWqIInsC8GKLfz
G5jphTXTAJuEPpIZJ+pJpKmt85G5XLVfq8Zr3Zr+mHP7Epx5U//YhJAhreuvJqsB2VWB3tGojDpj
m6jxi9MQ13bob8g1CP95zhpKJkR4cHlnKXuNah//xrpF5bYhmhRzV0ZSRjwy+rJA81onx5L/nNHz
d9IFwWEd2gNtj7IaIwYbxofEarky3cTjBeRPdSOwN8MUD0Bs2oI9EG7fIxMrqXUoPCNpDx0SYMGl
kgW9bcZR+5fVXpn134KM/sKMvNYe+DVQAozLhFbyJWT+FAOnkl9pGI1YVkljP7gZJxahF67o+aJm
5g9FwgLgFWNojapTY0DzScWeh1g/HzB0p9g7J50p1C9WxLSAGZorhOdYWEdMArngVW7W216u0yB8
au65Vi/1yom+5q427pp17Rg+9lI75nivkXMXykFGUn9n37RG3K0/bQFiY+HvAL+1zyTIOJ+IsW7C
UCTrYuny/YIS8a4YmZabNHg3Y8atX4pEz++5J/HPAZc1LVkwzeIhXQeXjnWD/zmEGQJvKX3Go6dF
JIW0wcK8F1O3unOttLJqfciv4/Gz/hhGabKWVqw4vX55/GElkTkAOoAwJdmkHtvw+JRjDY7bncPL
m6nbAXETYFB0ozHhihzKa1NogAvL2ex9pVDvVSqKwVPSVexkTtSLu5WlyxqV7GosLTgNvCgPJuA4
yxCVSdUET0iK/i4lEB1RMdCEG95L8x/3ujBproM6f4QF1xWjq3zPePBAzxBHqKvF//VWuijUHXNN
YcH36wHNMhdA3Obxi3hICs+7EjVrln6ffAteXL4Go+bywuTgvNcdIllHQk9JR+unynn0X7e09Q0W
z6eCkjYhff3jrpyjIbX4sxNPfLuPJtZ+XAndrZGTE++fFesDMa5f/nJYTxrCcMR4k41Xo19wSJ95
bEMoC2Owe2jx0WvBmfx+21cgBY6PnJXXIeC3t2NFcG0/cCPANFZHAOfDVS6tb98X+6He8MuSPvyl
6Uw4LOZMa1aLbdNuf6Gj68GOYgFNOIlh1KoYvIBoeEBebVMc9EjMbuJGS6P6Q/0xlXp7TEjZ5yTn
QY/D4F38QbcIrbksNFsYNmsh2xrZxuUhwzxEveIaoXNgBP1XSK5sQlqTR17KC4/6NmI4TjtUerkD
JcMnk4gFv5ANj+KnK0bFNbCtp8DIecMBzhZr3IMSlOe0e7/gOJRZwNnHnxkwaJEP/DxDEGACP9qo
igVhvnZXXoQxlaupjjgf1Kh/GjE8W2u5atBsa8aX3E5VadL6xGCQ5i2JhU0+fyv8yKHQuoGkMm8z
XyVNIiUIMVr0y0YGfKgJ6mbeJ6flw8Hzd1iUZUI3J4XkJXfarmrNC7QVxyQrV4rV3juF/cXYgjMN
EBwF0EjkxG68QkJYxleAkUhmZB6MQqTfY13nxi1Oq4iw3wwN2071Npg2dAMxWTUrBn9U7Y2oNf9m
qqn/j/ELoQug7NZ5Z5b5d52fZlU3mQhgS4PsSFDyq88AU66g1YtdxCxzBf/Vz1CvlLEHA4itp4T4
7WC0jUAF3l0j+pFB9NpkcsdbnV4LnWZvXfiH+rVETnhu4YRK8VoSMoF65bZuEjHUJrvA/xn+U7q7
Lvsp3aKw9ubAYqvVlQFqoT8z464cYNrDTCHDmV3j44J/40UI+yM8OYwZFC3oMvfN0L/EsanPyrkw
wfM/1qCWlc6iMm1a9JLXM917G1zZIYO8KIY+jII37RYaKqU5ELdYfyOO4AWKy6wbIMTKBIUad2XS
nPwLirvVBx0A1InnuUQi8H26nBidrxFTsNIEv3D/I/3OLakTXBXU8XBzNb93kr2ZC5wVfd0Xb4c5
eq7oQDWqR5c5TNPM7qGKMPM2JOy/EcngIe8R5HSU3nWZ8V/QDsAKmaUJ4VrOtFutFclMk3VfmHwT
9cjJLq+xfUrFsBXa2mbw0jMoZq2VxKcwgIgkdzqU4nN9omgj13nud7pv8r7cvdoapb+jLTiZXhBk
IBXTBMZykeaHu3HrV+NwzPKPdj08pAQJ6yzG77S+CXl2XcQfze9wDjPOUENbORe8XPWvH5ZEZ1Cs
DbmCXYXO5ZAZWPcEx8dky9Ne+1/1zsJ+RZLr0KmZey4rcra7xxjgiF7yE4Oh4aP7tc6pBas1Bn86
W63wav0Nyr+DADk4iXVRA2mWqhTA8N2c9ByaJXz7M6i4e+kIO+vkrsMoNSzaPwSmqxZ33+8xhSP8
n+pUVfNjRAjreP0/Np9Yn7HSG+ixeB3o1LvDfEXhn+1oPE6rH9QCcE+ft3iYc64ZFirv+1GfLev4
oas8WZXXQ+Ta/Szbx017bbtYz0Y13hsur97XpWZ5sv6StJAw1n0vjcxAna2AF9FFCWQVqNaT2FRn
8vKzRaxVyPHPm7yiLpH9qNz6je2EDba7Dab1ivWRFZCIbiStomxC/6/+vVgYPehFy5aO/gsJsbR0
31oFJOz298H/MMDN4jyw0dg9gZtvJaN/FDk6EOX5ShkFnUZ1AsBbGDplgLbpPQqJiyQpQCBVDO4A
bGljCXfFmR6gEXKRojGoNzuuN9B1Nj32RbmLjkIfqvhpej6vEnWyeDr+GPWWrcoMKeHghWlu0XIZ
jmM/LAdqon5zGe9xJD8K3X9VELlkiY9+1f2x3kxm+Ip/wnNKAFs9qfngaOXIBYTZ98dsaff3AFXj
+QgwEdW3VjXOYiEZOv4RyWlHP8YwrjdBTziYLWKQw/56Tu1NxcjgJep7Qc+fFY9rSVX7R/l+9ga5
PvDUL/cjI6OLhxJkY67jlWcBS/kPY5JY8oSUGacs8k90meZJyStEuQZEIKvkc7c7Mq2tP0S53gLY
z9GsohGHsrJTWwgaAv3e4WOmmfVtlTDL/2+CfjyT7ObOU/JicBpQrvNJ5E7rQOxeTwQwW94egapj
V3fcCZDYfAzER1Sz3+iI0QBbdH8P9EoHlw6aTjn9Afcr99I4Dom621nXNEvAAmxq3zOANDb/K8lw
p8OnJRnSzi56gCpNoQ/TVj8RsjZNCQJJLv7Uka2PnTKU53F5O+hoFTmSd1iM2jm+SiqwgYl5sL49
uIvuFnQ5Xj/N6Gz0nRp25oKUETiT6pwBat7FycdgiU4VVtPxQq6/D7IFUcuixPkOADRKJXmqDpL4
0hvWNw2M9h0gGuCCevr7zdXfvBNVUzb7NyyfeOtizTEzLndWwkP5OAp3NPQVDT9dAqzHd3cNmQ3x
chMa89f/BkgEY36C2ZhQjdmJ7w155rmSYTAydD+tadpsjheX8eS8oKjekthxTvDwuTJF2bJpUuXr
gvDAVAr+7NvQmz4bJJD2PXwB1wCOr1pmAM+StxDR0L1krEj7UOF4HJai6icGGAIDoaPI5/mrqs+j
970kOOdmy7IJKo01cCujOrSwClV4SiroFzEv7YBIgS9f5WjbeG3nIDlZjQpoZGb47X8Dd3Cy4HEe
i0j60Zk+TmbXydl/3lriM9a2SoKLcr1qTHx5+L3n8v5AKmjY3uPva/yQlckjV/GItRoGar5+i/F/
lDFpXK6x1da+ZU5zR4pVVb5I+6yx349Iu8qsJagM3aiRrgBwDxprMipJDPJxPajOey85xjSL/hLA
pCExp/Cpypevnot385chtH6M/eg1CltuB1iNTnnymhvqvTNG5a0+tK6K0fsNfqPqziTpE3kecmF3
1xIFnZxLB0EaUt2wjL3N4VvCJuQZRxuaEhAkTTVhLHLGPeEUb4SdZ2v5PDkSDz3yFC3JYGHXKx84
RQw7cxcdpYPMs3frv/rydsFEQsxpSw1G7ccEfvfdPfUgwiwuCf6sYPZxjxKa3qtOzaMkDTk/HM9g
9+Q3m1lITt0PsNR7FfsVhso/Pr9lSHOVV4CT7ijXm+ndGoMskIez9wWrdC9/vM4ChF6VMsIxgx4l
D+m9B3DkgSnPLZWtnC+NhOx02hhQek2fTMAK+5hayUipsSOU3Ex/jFbyEaDU8LVZMzhaa+1xWEwk
Eix5dD/8zBAYJGk+8eYyJScn81t4w94BrfnXx+2tgN66O2bPXPSf89LVGe17oDH1Cm/k2BweEQTk
8WmiOMsc5co1Fuz6VpuwwwPBUKkAWZbGFoX/sm7l32GMC7prxl4r72WKAsIUSva3Xth6WqQ5EGmY
SAwccPoFe30bvipnnu5Go+5rOa+8nuslHiBgW4xZRqnb7GV3aAeZMi9d4Bs8hpM7HhjxAGUfBqGL
sAzX78P+u5RXizTmLi69ce4HGhRJYJVjYUBl7BYAU3LvXY9aEQ8l8660TG4edndRGfL6KX9SsYYt
yVjfmMd9wd23K3wyTsDEUPNC8FNXkOYDeqBQDQVbO6WDtBjVTzzwqeKa5siRTR957UfGLwifZcg/
8g0YKmlOrru7CfD95Be905VlzW8HCDNTrdn5j/d5953e5ZYV9YhCX8VqeKzhcfKvy87wUFDAe0LH
kJTp2nCfeIDRPeB8k59ih3G8Qk2Eqvd6kzvYX65uRor5cwFZYi5RaNq6vWUf3BujQHggAgt/0rS8
drj9VRejOO2vW430sG3JK2nr6CL9QfffYErLmpmDPOi3wSWX3aZZ/ho2fQe+IVznbbKZNgsoXlSQ
tKMow/AhT9ol88dyhlMLsu7gEc3KG8TG1+XPOOo2XTn/YF4ugXIfBl4ALFU7A5/OQHLDqpy3oyTN
LLYvnBiksbDO/yuoJ65pft75B3ST1e0IJOxKZSDRTcc/meX7Kb5MAACS+/AVak5G0YjBAUqWO1M/
O6nsrAHJ9yl49LBt7ayEAbzoGc/mVny9KIUYqwgjnR1B6vCRxPHWXGmcFs7JLLMiwZDWaXnmIKJ+
jTFKzwzaCBWWxeNRAHghwOY/0dNpG0TTvOYxtPRK8YW3VlSYOvVZfmvKC11Fdc5qwTijzq/OhPYp
TtE8xR02uflmkQ9qX5lfGgdVl+T2lKjazmwDL8r17JTblOC93a0fnPmzQdOGVHTcKj7ZUpYw6L3y
l2UoU1Sf6Rs7IxE3o/M88a4+AxJ8bLUSGag4kRjbmfc5by0b9n3n6Sx3ak8zyC9E/HvpkP5l4Kwg
T2SOqIoJ4viC9725rLf00dT+j3yg18c7su7pv8B7uq4pYGslsLZAxioWE2jrIbhQ7Q5QhFXfpPiJ
1d9Fbdvks9oDqeN1QIiaZIlmhTu9on9tkIuVKy83tyK/6x75PHQVYiEqs8lZWfOYG3CCp1JXkfqB
n5hHD9oGEB4t4wmiLfaONVkdplIQl1J5Kk7EJUplK73i/gpgHZvseEuToE7wQLzwIBdsuObVM7An
Rtr48UVgjsLNoVg8Pm3vDYsXxoTJT1+pdHSSboaUbQvI3ck3k3nsRhuJ2gyWitRz40UuMYzF6oGz
iAAkwd9SlHjVW0CTwHoAYOF2Sg/yufzJirzr2KrMsOpXIWcaR3ecUFT04jaAuJ23EH5ARhmXp3pr
NeAOHyv2Xj2+E2+Vg1x7bd15Lez7QjlZVURzZV+BXNr6HTqJah5C17iscSd34xH07YRy9zbZdG8A
xEwP3cm5TC2K4SQutYf9JQ0yK5VQIQ96iSNL5I9RyQ0+MbTxTdZsLBYtyrYujO9x40OVoHv5Lc4E
7Y/0DzWNnj+rrEBs8mK/HOwUjlkz5kMemcZcGXLGSNnN+fmchljw63haQ/wJye2mQfaabIgXWvQd
tX6fqvEwJtB+Bog/EvgFXnjM05hoZakgCvijte77hARVBeZhvaGp2Zod8qp+JLrpJaxxmVSPFZKx
vV4mH/X5k7L4TyFqZqph2uK+dNDCTIlOMjW0hNWFuggCOm2NhTgAorbftyA7WVnG2qHLao5GignN
MDVJsEs4DHI5p3n5rspZDSfUhXrU2tNd8An7rlyPYBKIkU+5R0wZPOZxm/VkT5ssvnjl56C6TxOp
AQP3VzuO/vnCmh3jiMWCkfXmBObQs2m/tZf9RSIjYt5i0pRX1F2TvNSH4Ogkd+ntFE/ajFbdtSer
JHYMcXUzO4GhRHN6T3QQoa5NDNKwYBGVc0UCiv7ba1bfiWX6xQTc4MO5fQhpKnpjmvMhpDUEte4l
zgr++dSVr0uDAbwWzLStuR5OHWA71Ayq4bbbfHs7X1VMMJ0Anhl8j39IBF/3iii7kqjwztu/v7J6
RABaT5qFiaQmBQ5n1h8eG8V7O8taS9g5lCas6k23tivEeuRhHuyDqDctlX0GSW0jLDTrGYeVX801
JXzrx9ZobUGxbrV+0t531sUpTi3lIy0xkByRlzC2/+Pgo+whs3ubKhQgInIqr522VxWCWNaja/z2
JseR94igsJsSMT0o32SPEKRxE1KlNljLBpClPA3mXiDNlq0xmoPcm1zFvITkZfOaXiLGNmMy4o6W
V2CCyU924P7Y1807P4ouHiPNZk6Eae68Podnbh7kDDOwGYzGcnSKHQ7Q7Us9FrnLvMren7TIZgwf
sfqd8lOLS1wZbSNTYAVyaLOrpI5Pe4qptKU8i9gLPzgf6fxGn+9G7RPwhRCWDFGt5fWbIHOsKnZR
mJostat61tBq7xM2hodjaWuwvICR9ZMh1La9y5bi1rJn6Qu0t9eHPMqndqjIDLvpDSLLLBAwT3GL
GvzaUZKs4e88L6sdlMfL73C8MKWDQY9L2r4o0aGyamRiB1mYycf9+T1Z/Izx1TSnlzmRWAm1zw2V
VcBHMrS5fwo6MB1dZDQhIm/NVQE44cyB/Rq7H1YtngAGqzpUIRt+vRApyl/VzSvG66rq0Tgt3ZI9
l2YRCiLqCo0tB0WjJdZmTFDctnt/0AkNxGnOoxsfK5JTR4NAx9XnN0mBnScmxITgr5ilDJySdQpm
hPFWAx0Sa8nKuM0rcDuhPDNKqtUH5Qi4NJAz29/Nx6RqO8gMSiVqpH5IkrTg6IaSmqRyOXyK/81Z
QNXHYh58ysjllkY8B2N6d88LJT0xPa/VtiSrKF7lLkB+oLvXNJQsNuNMontLEYwWLIN7Q9aVfho7
ZpMO+iEKmdpmgUrt9+psUOKniBcM7dJE4G7CXQgyGz6bz2oUJ003s0/vBkiEWUohLhtZVndvTbiG
vPKHpcPFeicYYGPJRQ5tphdWA30llIZOy9Wwrlj3AAbdTM/Y7EqFtczDOeOg3xy/5zzWB2Uukqg1
PaAkSib5tgBsQTMr9DF7v6TdHGEUOyVc7P1VFPhxi+w1XpPWucTvf1qhC1cNyY6ClsNECgMmWOkG
O1z99DrStObAs676PtbFuxZnVFBCVzeLygXUOiE4rqaygrTPOVEB+vUMeA8Gjh/iDSCBm/BxSSrU
CxD1xuaCH0NgUtSYL2DPC2zO50rx3pU+OaOvk5S4HXwFcRsg5XSoVFNclz4xb/bSqte6avliq/Hh
Ec7tIKEPQATlEW1YUkxfaWP0Wo0NGnPxHNfdRfDphLIo3RMx959q6mJD+JObvTb+63aB4WYS5Uyf
HX71baVMhWFfTsv8hbrbf3tseI52P614QFu9qlD7Dx20I6aCwIStmatyhUtGo+muzGJZ/N9S/9nW
M8VD8yCaifEL4tHIt46zPiyN+ElXoY5RIx/yd1ko8NiixGCHlt+igVVVgiQ08Tlwnw0v+R25tHo7
kncd4dF+biGxk7I4cPHeR7iAnl5VbRN2KnoPMIl0eEQWDnqjy43nMJz37Sbi/vMK3kvCMdog0f3I
DKESXQzA3efKQ9zzJoJPlNK9UdwEKK8KAjmeLLoY6of3TLX12AG1vjOh55T7Enb239OURUaSMZpV
cSgwn0xaWGS5dFge2ukK7pt8wU7oQXoIh1ZNUyf4bpuUQ4wXA07hRPVXyfxsMUdd2PeHZEG6+xjV
2mD2p4YpbyWmSfB4jreGzMDMqonnkmMSqr4C3lVgYch7k3bZQB7ny/YNMILM4b/vSIghyNSM+A6N
C7TvCOLzVI9qZIGvaTj/yK0a+zwSjYnwOyjgYIOwztgL7/ePeQe/V4kw2JqFYpXB+2A0PV7OyYze
Hzgchwiv1SLlOX6WQHXIJdliUTrYrTp5JYzftb7eOyz72Xjak35MFkEYH729fPNUbYMxcj+9kVoG
edZ9d5kWuF2Y2qjo3hSc8ocWtI6+VIjdX8wf/Wi//aZ8bTE2mmZiqqss5FzqInHMbCHrfhe5pC3c
7vpshojsWgpvaZq3gW+cLSypm9Pn2nHugeBoPNLW8KPxamZTFjJafP/Kmq9K+6a/DabRNu+GbCtx
MdbllRDDyK8onlorOSMEj0c8OeU9F4Hs1uFJxh7CHc1VfQMlh1iFzO/YoyP9KctN4lun8tdwJOp4
cH2DxwTpBfMHSeBd6tcMJd/EX34u6vNAxCIhSUVjaIDRQWTEVZx3nQhVo/yt1WLfjXSnbXscpufb
P1SFmqeQdLGoHN3LQRIRRm+NPyOqEwf9pznMQFS06i1eNWmf1lXiv9LSiY/bCtR0cQ96QwVMVOPz
dyvBRXst8nHGApsBeLxhsVTtg1YtHrfBF6QSq/HCgMdx50dIafQPLfLD1t9xGqsNtbO4V7QibON/
jCldRySvQRtg3Ex6dlFwEGThFMsVRmeiYfKKxSHJwdT3jqbH+/u5Go0y1QdDXlpw6cbei8q8bCpG
8v6qPzwhcf7CroTgkeudrJWEo68RlupaSRYwB/Jw7S0jWq4Zqw3V0kuzSaUVQ3zmFrfqR8UnMlG6
Cnb+1qMC1Bg6RE3hd3sGmguX709mzcR/ajO96KajrBgWRg3AgPpr2RLQYFN9oMFMRd7IWwmjcg89
KyUInltTw0gRAGqqwEmy3WdhQFCPOzOYik5EHwYB9mW0Pq3Xe8IuthVyo9fPlSBa5K0L4ac/2cyc
J1aeq7yKyCx/8Ql8WhCvb1G+ZeZcN5SNmOC55xSey+GeT564KbZlxSm6TNERCOvaZAJ2TsVRBnwl
cx1JgyzzizUo/A7DcCtQjM7furuiDDah+ujCtT3KScb4f5eUiQ0Sg3MQa32KzeOYjxhPf70W8Rij
oInT5B2D/8oFQe+lhn5Gnvp7zYxPk3wPSTJygahCUoKlWhxv+YletWYqZRQmvhBwAxbp7ktMvmbE
/AkZcwEsb35rsU+dJ/89YV1Tqh1SQWiz/U4CnfNANKJW3XZ+rnWrHaCxTNdgbSQoQ2lB0JL+fKHL
NMHtzm8t5dBsC5ivp8pyCo8mF30tuh47Mey5CxyS6XDENFW1NUSvpVVsQBHZIcGpwA9eiHBMqE3z
RfzkzcCvaq4GWKQEjMAoOljE2RzUydPBc19f/KqCWC4FeStD3pXNffEUe1bHRgQP/sHbrDq5kN1C
dn9qeMwWnMMlQQ537MyKQ7kMfJigF7WXCaG5F2hE3gcRotjuwyZs2+ZY6qVCHRx2lrqw+jiHt0Xf
kvjh2R4mw3P5+AUtvhgAGJ+jifd0LqnyPdmMksXod2wxklbdeN/0dC/D5eUTzEc1v1w08w+ZpCDS
j38YI8B9gFGBMb6rWQZ8hM9n18Qhbya+oQvGeaxgfq/G017lr2Jj9mG46rwMbARIW1IJPwo7Jtbz
L7BHrJ7YOfb/fqLz5FhoP/QKVS4LvnXCYJXa82a0wp9ENrmaZwEhLo3xIZgZarJWD3X/sCfQzCQq
H2YfIEtIj1UDdocdzODoxqIjklTj2p4gUIOP5ePkbgC4zXSRAaPzhBFbebHQvjHWK19IMGWcQFdC
W15MJqm8NloU2uFBtkDtd8RJKdYNVtdxbl77r+Cnbcg6d4Q/xW7CJPxvny5s5x75UG+9hVlhCHi3
0jeyiAGSP/Unyjw/BKUPMwpIqmNU1qq9Y1ZyC9lmNzhreV9MquSv8FU8w7g2LvQ9vuIScsJqu7Tk
TmWUByvJqSxyu3KIKdj12XPshhZRIhmOXz3KpmQhhlC5mZ5JPmEhHMysKRQSXPLGS6TTjYdEiOXn
tz6on4CszTK7UHDhy1+FQwppPiypJHEyx6EwHYDUscldyCOS/6EcVmrl3NDsLuXDddOZ1PCJ6ult
xyhNKLh17OUt+arVJIfK9tykcfg6im91U0Fz54CrEX8H2EjaUU4ZSaIWLkRrUUr2+nGc3W1w6Bc1
3EX7O4IbgtOM+Z253lc+IcPqcFnC2TvcP+/Hf2w3ZDZLtInd+vg27Ns9lRCie+HH8qnET9MBJ08d
DbA4ocLU4x5jNBLJOIrARvT4CA1WEUcC2Rfjt7IjES3NjqaMpG7JdGpCgb2trgTISTvj2IqMZaRa
xbX+I7G1QuR7yIzMRqqJObp4ByYI8xGEXts5IJ7ajSVcuf0J2Eo+TtcWnv4Hn4LJHrRQFCbkEs9M
UU9NQlsBg7oTFnTKWA931ZqtCQ2Odeahgf4G0W7M5PtO1EYSmr8KgzdoN3+/W1q3jD6T3U4hDre6
zXoJBaUmVT9u2sA+nIFQ3g/sZtVUF7qTdNbfDrvfCfMmN5PDwoGObhsimkU7Rcue6Yf+Ka7X/yiw
q3aafhdgSodDY/WotTrP9x/upviTi5I5Ixyr5f5N0Bd+0vy0BbqtIHjv1bZ62WSIes79+sG+ZF7L
fUmum21BWSs66m25bMKA843zu/xUFHCXnoH2K2Ob8ysinV4LuEnffG0tOx6TxhreaM1H8FDGLlGs
q0FCwfJE56cSfpIqihXwHDKXRsvLocm/+ryTaqnE1csJhsa0LIX65oIo4GW164lozinyICZ8pcrQ
+LkRAYwWUBhQVi7rg7ooYDYuK7cUdOpVuKdUd67zER0lju+vdHCfrZlO8vQdsI/SV0K7SsShU3bs
DQRTSn0v/2BWWoJ8F0gDhlcg8aTo5nyqY3xu9+L4pQjAqAEPPt8SjARhSLFtYxYANI1eJDVZBU5f
e0jIFfHaAQ4AE4Tr/7GzUDTqA9GuXg3ayNSGWbIT7HFw9ni/M4efruDME7Aikf9OpGOdCmWoLvQy
qcNQojHmVAGT1RrGPgRYiR9dmTFj3Y7+PX+Mm+78tPxfg/n30Q0ztkXKLzaqTbHzyORNKDf316L7
MZYISYjR8rmBy2ABvSKfUPsEAmUKSqa100coEHG3KghLZKxC581NFyagylvyL5WK7auP3B2Ydx8X
QqpBC5H6AJwwPkfqqQAA6eF9VKuVZD4/XRx9kPNqxA+z3xxkIwUT/qpC6anOvScWY+TZ7M1ZffIz
iibcV7r5yP71DZS8evQ6ItDcHgba5Aqvz6uf1mtULiNtUCd28RKdx9mnakfEylA16WhmK+mc0X/2
Yzd9esRbWbyaOKETBkW5/tuP+TLHTacyhhNeorBVl80JFs4WUpFgNe7qKN7bFe/jwrVAyY34gS2+
Pq+OY8TF8SZ6XL/yAmxsmarurUR9wbkq1ceEfpSSN0IrxVkY+datUKzow+Rc318sRh9zEKZHqkRk
aT8/IHRZfosw7Rhca0+gYA84gyWz0vqpisbb5m0MXUJuVAqri+H5GAwf8KOJXh4BbvHTbQaOg0Ce
JREwSY9R+gzTHN72ODzPlRzwdNdPkXOcKU1NUSTY+44yIEFrr6MFdF1f4RTUSHDRroEv3CWFKrGN
jxMnSHPrr+CuV4LqeIHREMxk6FHmEJyfrjpo3bYiflcEdx8hJkASJbCLnVB0bsR2YbsXL//ycOUV
Et4jgPTZtdk/Z3uzXX6QaG5U3ZNCowZTYAlZ5FziyOIQkbs+vBTGa378eckJOZrrO4dwB1iY08Nu
GcEpiNFMirA18BPyR3+aHCT8cOCebZcHtLutP5ytKdNexOui1KkeY1MiYICXuBoMT7qPmGka2QI8
qf7xFR74NdJ+l9qJMLv8BEAhFotBEQLVd8kL/bJScNnwTVaIpYNfzrlob1PTFQq5IWIQsFRKi4d8
tG3ccD9+6/S4TAEpt/3pOEo4FJWD31ZJkGo0Iv6Hzlhi9AeXHzW4IKirAHYq25PP33N5W5ny4sHy
KWt1NWfCf98kLTNwknDR4vh6tfGuG105R6DZtFDpEDXmez3GK9XvtSwdY8zLICzaAPgxYBfvrAU4
Mdx8a/uH5HksP1yZzXuXPZOLvuuo7tayvER+065/Itq+fV8nCf/hyc6x/NQsQ0Ws9/3G/KU3I+PQ
2lTSuOc3Ut4g4QTvAIFINU3WRv/Dendgfq8MDWjFl7yLTPpIXYy76LXhHeDNC6F+DDSE1lbbDyUP
YqBHv15IaXSnPuEvclqOjYdELlQQuiF0UI7J1rncMLON5XB56Wi8xNyHQtC/dSib1PJFwGjAbgWh
/cLf7NOIOA0zg4ygf1c2j3kAa8jYEJ2KB9Hp/AwusjfUARSgOdvN+MpuD3TIPFtaFgsI4Soqn5hx
NH9BcRU757dZ3JNRmfgiaDdcCaH8LCf3VP+Ijo8O7VCXTogY1WdD2w2kJFgpeHlLk/cArX57D45J
tq7C1di4QzvA8pA99BikIJQ6NFzr6EwrP6Sh1gOalra3kolw/hh5D9HT9mErQUZP/Uee7CHtBmi5
X89H2YHd+bSw+VZqedcxpKCnRPvg3EDJoniGGEf5ZaiIKA3vFhIVdx/VIVNuJi/1RtfV0Oj3EX8B
/0ihE3wFebrC8MoGuoK25WT4B9Q4NXwKf/8MWXI41VcIWVf3M+l1UnyPwlOWIxA0Zn/AstF99uu/
R34CsaL+AQ7F6OU6melFjC4M0u+uUamZxZMTHbOThJ2TsRkUArfA7T26U5Uw0R+ecbRm6aSpsFSi
gUp2SNWeKyZDXnseM/YraYRAGrLqUr3peYPnBsz3XMboj103aVg+abm3WuTgtSKASI62UJLHs7Q2
gESPHL9bXWqGoHmb/CZeWKY0N6ZHcReJJX6c0SjeqB+y5wE/ojZZsXRsPTNVCKlQCOHXRM3YgwnK
CIimOibjNauwUOWjxmcLu0tfgO5YKFtEevUJAeEb5ml8A3Ki+M5QaHgKpMNrX38lfl85NcaT2aWg
8o1gSCtxauinwEKrP21CnzrNv0ydt9CwDMjIIaNXNiNVmFuBOds03VgO/smWabYnkmi8UEzltCng
o1uI9tZb7CqGN8PmP8G4jYLHIJAS8R9z2OCPjaOG1F9VJ4dIR/0GEKvqI8cA3vS9BgiC0GxKbcag
OCKQ93Woa2PWUHOFI81j04okMhdp4q+xJxzU60ng1MKHXlySGg8c4MIt5xfdlqgNgnrbIcUtsIPJ
M+NzQ0l+V+qELl6oMWP7jGNIuECuXS84JsiUgCgppa/gl1YqBPOs3x6g4eJ8PhAu5K0rWaEBhiyk
M8egN95HUMeWEpPSHTWlS+3OX1p1zOVFMALRQByp2szljoVgnyVYGasv5aloPkNOwv8h8xp4mpXJ
EsV/qe+73cf6BAeYzI7RTAOZsskvxkfuACi6Vg+bzMciD0JyMw3ryNP9SdeWT0BHqIf6CCCgZwi6
bVFQDPzqOLUiNu3Rk5s63tmbz/kseItn9CJ4trIoRLQ2T8/Pwy3cz0LP1AyQmkbZVaGe0q4j7oAG
yqwh73ZZN72o889g/bMNKqHZCBOG5dSL4a7MFEkUaquuY/MOfJ+rhIaciM1ahkKwaFdIv9wIDIQv
m5daGnO+ZO/NN5UWOBXP8eoQTB/VovkLGk2Fhv72R7XziTPoVCcjvFhOZwbAHjHSgNE5rNhw/2l/
CQXcOryaFniS6BSUZJAG/15+NwFcWPkm+e3LDNehZqwyMTq+xd6u8PO7j25e0ueo9Nr+2+SnkrLY
+S0y4kdanJOSoRPSgSus+e0BPcMCMlTg/VNcb8KmfcLa27juYWL4zQnT/rvLHNgwCZE4dkO7B73o
quD1QVO9EzAsdCpLxSY4B8T3wgwAKLcYk/urQwNOEXyW2S3+JhZ30pV+jjtzuMjZN8Q7j0daBRMM
IT/iMjyRoSlgacBLFrU2pAVDovJ9E2bmHhrobqS25r/vGgjGUQi1HU3tFc54b1GM+TAKIT9ru5yC
hA/LMvel/kKe3S98TLmZEF7iDYcGCc1E3dMh3kL1O7irKZyjv5lxk+pTj9f/wbolnU8nG7yGT4Lu
n3e4B6UK3dtLw744YQSAOyUumocGr4v0pxNvN6jrGi/L1b5ZOFyvefVwg2+Myx1d7pE1lEuwv78w
KVaBCfr2p99qXg5dJJKM57pQBdgD43XVFCPTTthDNxnZBoUg4K8gXvtLGhoAFPyflY+jG9ixQbmi
w37cqLLb6WjKsDgWCJrGDRHawkap2KpLVGebkc5TGF6CByVlbmMIzwZotqv7TpyuowsH0fyrixpW
KLuqwy/HVH6rLIczYO0nYlfJcmYLEK95lEJJ/I/2dSywcM/iPVDjo/+/3TW+KvlUUEjXdk/nELlm
d0gAvH+5LY5Uy0FId5W2cP28gvoLKQNC2+mSqK9vuw4+XBPg6oNvjpO2daTcoA6VutLY9k9/aPki
Gd/j74i/DYVtx64NbZzTFErf0jMjEeYj4SbfUHNvdJXvFyrk54Dp0WF8naFWPtNtv9nFuTK74KYH
YCZaeoulNXV51nzD17i6sFtS7DTnXu/5e1a53RnGnozGgTeYtud+fuMlzy/l6u36XHbtQTm6Xsf+
x8Nxun0El7YgIAUMo7UGxF1SHMHnbfohXaSRrHNpkVbJ2/5yeqjJwGNJsXZ6YorKb8/jBMytOdUn
Vw42GvomwVUgfGw6QHdDU71My6Zix70Mln2QRo3szsHqK+AllPsreGTqrz7PA26lIRG7Oo+O3Mfq
SDgZ48nt+YmB7N99IFSUkxPYiUaUXLLe2kYloQDPbzliMduRtPHuUe/hceAvL6wzawJ/W0EqSPu1
N64rfvcYgjMKQrwCwWcFySmHkGHNfxgQuvQcS8rs2lI+ygK39xSoe8KWQ4vKY0aEWvuZkoi0z+cB
zn1HUXX98Ut4PVcTcvsvMp/l0+EWoLMzl2W6YxOHeq5M53TB07Yk3nlERbMsLvZPcz9L/c8MsQ9T
IWrzDYaLjhTCY2VksoI7gnXVEexfu65cDvghwco3IiuHjTUdeaLxSEuokJkO/HZyWjNyqyLOTqdh
uzHXF4lY6DN17XNYZ35LNR8Hin6mTrMHSpZRZxYvZUrceHjQi/jUNlm/YwUxEJOP6VkFWPmHOv0/
5Lf9I4DCSh6lbBEt06dgJloGiqARWGshSLz/LON1yG8OkwGusfZu3FL5UNDRtN0lK2hx2NWPpmnf
J3OQJwj7L1RAOw0tQV8+UuBrBFKr94BRlpOPYccSAZjljiEUDLi2fGKMtXqvm1A0zHtpaErLyWzM
WWjDymxUNMtzSFwQNQpy3RLQgs+ew70HQ3xqF2SZvEMnfrEi2iWiIFcS80pNLgu7m51V0+LW637Q
RHcIqaWJDIz9CYrvqh/9mm1qF0/BgRyRZZsJgmC0cN5NYo3SHlyjowOSUsiRBXEEH/RHhwQOGCl3
FLaOowUEuWgJes8ReXjmI9Ju/nOfeTGBLktHFtj92EcKXgPXeSQcRJX5D4lkjQFd3WEM5xRModYs
0CNGkpHpKtl4TIU3kZifg2rAgT74nFj/NpSgK9BXFpxnonnBOLbcGPRsCvGufRVBPsHfnoROTI2a
yPZ4eqvWCzzAbuLWyiOosEdkcuqJ97nf8uWoGreCqkApp+OErqWxAao4RbUA9UVdr86aUCWv+vob
MDEzG1hVIJS2fL1BBDneP3J5yhUpjqZiMxce8LHWJyBQvxEnydInNcE9bcFEhgxsvQQmHa10u2Kp
cM9Pj/3TdfiraWmfl3CLqWH2INj/11ScOg5hBYwSf6O3Yotywg/Uzpou1ztcI0HRmKHL+DWE7HIe
+OXiv/06Szl6XSuQ+uUhcwv/dyPLs7e8ps+vVWvf+byx/LDTfruG/p3wWn1xV2gK0aYFtnf2oyZG
hgVbDxmHhpD1bjf6iKHmeeibtmzkhgd2Sdnw/bZrAyZFJHPPiM4SsHtqkLHQYbfOqme3HYWhwxG+
EgyFjJ9OLblCRsHt9D8N2sBKknKlsD+qR7Ei48qjD4oyggVm/+6Oiur6AohBR1hzibKJm4mHSyjn
jP4ovTseCiQQToINLN8Q8/t9Qhxgd8kKkx2uwp7VHmG6SanyTDAwjI/aao/lgFJZqSHUFbEY8y2H
9PEVp5yerULq6xe/20GZbQ2fh462M3zYO175RXdTb4G5xBChA7Mb3HF1XUheEDJw5GqhinPKjOfp
SOZLZtRavFryqn8bOpgRYDjqeRi8hUGAxJ/QonSa5INUE8N9v9NaONvomBuS+IadRM61KvgVQHpx
UX2lYBZv54kJEGGqAVfnb/89oc40HX0EGWxz1oRSJwqIdXVuYnl+1GB7tquYNF6GClf2thVA+Hvk
oDw9nc9g3bqIWRl44XQWnXKAVlncQH5Rw5glUU4s7yl4qblWV+/LsBGDaGfWirx1Upz02sU3gX8N
jxKeI1hz4/kq42bJU8763iz62KSA93+ZMrTdNciLSWbQm0vbx1uJUemu/JYmW3IB+JoZtN2tZor3
47NNyQ86kLOnRjIJKU01B3SCZxcmdLa4Kpbb7kaoePmQmVxDrujHi3xoZqHgVGwJc8rBVwz2Sj7U
cebtEPmuvMCfIMlLRXVSrosugN5oxmJ6aQ962M4LxzfY5bXv1zOsYs0VgQEhA8PJM9shIB7kHnpJ
yiV3iOp2aeKI336BfIkYgBijY4qnD45cAypALCjLGZGw1Vr5Ar/GDVWFm6xLTUVLRi2a/SRXzYrT
drJBza3eB3QOW2diLGrA3xjEMFL97coSqnUE5H6IjgBnmM2bvC/JL2FUB2aArVHz1Aeo2BXPTP5e
OszP+qyjo6Fq5qTuQMiUP6leXGjsqGYjAa5FJ+ss6KeeIu/rCG4x2hc9Sb9vIxAUVSybT3RGvVG3
EZNwAA4xK8d4fYKWUaL0eAl63ZAa+dzpCywVaDfo5mT9dI0+jQVOxiCOPZrXYZhSuIdwjE2ImrRe
ZIfVJ4Xb39Jr1PSxrENtzjLzBcc61UUrnvvkDPX/CqGeOBkOfDybXWcMfPg9GN34CHtcMMZ/xPoh
aVucUEDe9+cnIzNzFmKMc+a2dlqVQnAYtk+XqFc6P0UV3isHMTtlclmfAJqAysmAwy97gjphm2G2
MEGEgYaCwQ/i2N7UGjcVdXxU5ClAjVzujzqNjjoLyQgSX85rfyd2NO/ZthHODSavYVqQQzvVLcZn
BTpNKATp3Z7VQeRTMeYqG46mVof9+zdzDUvZEfcfZtTUoPxpTzAauZ6qxwo2SHcM4uHmEBroTVwQ
fpURcXp4lbcY4l6Hr9NdCW4KVMpAp7TmB2v+6JeMi6IziL1zWNEDzkkGChPQq7yluNNImaNMsnWG
D5bewjIoW8g1K1wTavzs43vAj575XE40dvLWf1AB7gbVNGbxArNKT/h/U2tJQ8x2xqiBXJCrT8o4
nCzCkODChYUSRPIrh0bKHGi3e6DhFODyx3fZSsblHFFMffybYwg/xTx+sox0cFpQKNa3Sld4HpXl
xeHKCYy1CrCscRK1MFdo/46syLUHdR+EQzFcSi0/fJqRxvJXTCKACTsOOiI/WGeYQsbRp9rC1dw3
n3SI6ROr7aKZq2hFC3T4qoa3l9ZP1ZElrturhgV1bIPChE9x+fjMgMDL3Ds8Rff1DCOx/uuwd+p9
Mxn6JznYOAVK3D1gP7FXqsUYwiAV5/u/zs0+dPeoDKg9kiiS9Tq1hy1z+YrsBNY02D0m2b7YIPbC
dRQVgWc56oKtlSAh+/ETvUlgfybJVQt7ZKktvcuNzll9V0XWloAk9rmtj43zQ21rJSWxLsJewQVd
wxd3LOaT/3a3/lPGwPa+z8ZudiNqpBIoayC9GtfiBTxHFNcNsmzPDp66JkOPnb9TJmSIj/CpR6iE
HHIDcw8vcs7g6hQmohcceQ82WoqgvvdgoUYoZbR/nCEbQAF6IIfdXrcGeruT8wjiAOnwEwjI7zmX
N16rj5ec91V5Ax3BaPO0RfGVzBzdaVdZKiNzNMrvXpe3ueXcBCaTvGjOGaNPRargzBH7GKB+wTkm
d6asUKqIfFIWwrcW3pKeWsK5Ry4KC25DvG+BUdhzVy5tOcWEv4A/J5IRDbgHVJI8T4FfOJzxhGNA
IwuweK++8PeCyBg/0gpNcI5tI+UZARbvKPgeCbnxfQf1X+3hHkpw0E11AJ13TpiMItSIpIqTtZ7y
qYTQtlqMKxvLBv/U+p95SzR+f9um+oON7/FUI2E9z1hCQSXZmWZKGB7SR+ZtbOYAepmn/iyRWDE+
POYEqLFWaCRQqFC8slu0PaKqbY8rVwdo7EEPtL3IAEeCSgWe7BA+Qa+SpmZrqV10rzbcfIViGewG
fxCxtA6u85qn2RX1K4ifrX+22VBuM6PkMCNiMdww0USptgYxlVu9rbHDdPh5nHG6lK/AbejZLaVy
SWMCOfipnjserKg0yEwS/BmczlH8wuJPMvnJ5rsRZTmbnA4n44f5OEPL9hJS4VrJP2XpHRwA2m6B
gnK1dDL59lQpMBO/ZvcrYWfIJrQ22r+a/fAYY9r/G/sQdZU0iPLEQFNURg9morbdNqr9cZG3frX+
WuvPgzZWUsP+zL8JOVwWsh6h2G/38RaJVqK5D5rgXSZtEB0H45wGRfS4tjmPVB0iNrnzhxIU1m5c
N/Hz8ohQnn9VT1jZ9GSvlMlwq7MBzWWmJOd4m19TIZ1mQaGSkYI87t/lEBjmzmLsYGkfsrLxS1/u
EXNggjEdmA3YXKGXRLwVGTrFoipcCTKra4oQlwD/I9+NiuwfLJ9ATOL9U+EOcMWOdcVuwl2OqSRG
WGp76gHaNRLqLVTz2uuWAwdxAujcaMrQWmnrb7+i5FumD5ZkLjoSUyPoXRUAmHugwCyph9OjklqI
66GUMot1HtfG24Xb7JEuGsYe4uFM9SUcSoTGYlxkFyKYZIcxA39RCC+n4DYP844jxXoNMn7YWu6S
7z1pxSR3HJ5MPW//xn6e5LQjZ1QAyPNJvSmqN/TvEzNyaACog7g4wMVcuxp+3I24lJO/T+tKEo4M
OgeSfqY2o65CifakABdSIsjoHJsLH2dQLJ8aHrDjV8vu7uwMFzb/N570orLPeuoUIGkJAD2xBqWb
GJo1gwlDQrp86454kMlt8QTLALGVtb+Ils6eNHtQ99LgO/gJJ6/p12lLd0WoImkk/oEbcQNcmvh5
8XDEjr5Nr7h4AIWoYtTWeh2FyaMwJoV/m76xiTjs0G7N8kDCAawiBB2p0bbKJdY28nRTJuLBIcG+
jdr4ja109hlA7jbIbC4cDkEmhENTkQOd6tf15sfFbvT4HLLYk0uA7bQ/bhXdrtQWQ6ojFsZhpbxq
/qF5cvRoBkiGeF/107RkpVy6W+s1ij1Tjmx1T/SPt4nSGzBStbgLX85fhWd+DSHU0dSTMwq3Oexf
/MhrQdn9keT/3N/apIMlt83KJWl6tSl5cY346+pZZKxr7cOfZYagMtyY/24dCky6rrpWYOdCwALi
GxtxfbxxmNqRB78Ppdlq5iq5pDsRq2G8U4ixgBnA3kGSw9UprpprsNYYdbDGPd78XBt422m3V4K7
B2sdBQPPknyRCckPB/UynVL5v3nMQCK1kdCiLdRB3gpWV5pfEw0nTSf3xWbAH7sYzQy8aqX8bWgl
N3R3pToSs8FYiWkonjOd9zBo1Io59BI0Ffc6Z6/mwWOmV2eVIsoJMh1DiOoSlZZYOAWg32cKQ/j7
4E/QN3yE1oI1rDVu56PS4vkLsPiAiWIcBIAWiLn31lh+7ExGQ2RaopGskfUbf7+epedlbbJyaHWA
GpV/TTc3JmwYokPF+OWVa7Ad27PKyHFyFp6qv+Y77GteECJs0yBJNCHWPs3FrKycX7zclL6UTU4r
NzwwirhvCV4bswkldagigcdXx+7HGonTqFlAmMrEXBtRnuV/RErN7A4kP6fjLPcvZdNINOpmImhh
oURhP8pO6KVgNjekgNc+KQMBeIadDiPfcGqSUNdGl2Cx5Nx95V5nOgr1TNx4CzY8k2KspEwAflnz
R9jRBDPu8HqbfASMe3aWgXnD0eUXWxZjl++lV5bwH18OB8by/ugBper0FcB9MtMwDiXPzIj8U17g
a6OnuQmo3A74MBxxevYjxk38km9y4bqoir+TUDW1bqpKDNCmsKylBScLj92KRt7OInwzKgAeVma6
9SIsmXlO+HV1hQJnPHH+xe+j4fFIZbaMLkvfKY/nBfvfFKhsYmqg3+peVVryjK6uvCa+kkiulgwA
yIC9kIK006k2DNuM1VHhKahhth594UOG7wFYEW2WFN0dqFeo7fYCY/6Ek2yAYzXBslgMfQMUHojR
taKsm8otkiNLd7xZH9W8FYYgswkJSNgrC5w4T8FEN6//47bKPAnxOeviCeCkLEQrcxtr+120C0ya
FJ/5z/h+np4HLfKgm/NzTh9qDS71tu/Baq+3ZnjtN3mcwU39LTA36ob3cuQJ4TUZYKpF/ARwVxXK
6T0xgg2IJGJolKfzKmMRvHSiRNLmnByC2YHslVykDLUr5Z7uHd/mUYeuVG7ebFWMzgQGPWLWp0Bi
4uJoSONE4K0MamTlwQwuFVVgX+d6RGpNXS80kRlFLH0VPqEAueF3CBVM1YsxIer3aXxN+Z893g1+
722915z1II36x6SxafhD67FuUa2cwdceBsJC71KdydbzdXaERIcIxAYbADXrgRfm9K5adY7qDCg2
Ymd21rSQT9AhFJ/xJ7gEXf9bT8p8xc1P0b76e6w4oKDvfDwMnM/Yy4+a3VJHHfsteQrKYImTgHwA
A2vIersMg9L+gTnOXDFAKCE4vZXdMfnmQnCWaCkWRlUaYsNMijMnOs08X2/H+YZWT8c5JwsxpmRE
DTQf5NxH6jmSKqEXKo3MN6g9G2lx6L0pa3LxiI51lre5NBL66y1dmTJY+7QHFczuijCz3FdqGVca
fC/Avm2w4q9KXOUjYyro9bTuQ6M8VZM1S9qDblPo3OYePRY/K8xGSgk9ZL+G/fxkPoATNVbjyQYf
T1Uzul/T/w3QB3CsOScG1zdJ70Hg3c66FgIfNEcEbHkGp/vgI9Q81lRNP1t2FWe2TyhicmZRlvhK
TMqRyP+U6I5P6/8qEXyyX5JSkvnESedxXl6Lrt34MUd5BFhWbdJAt/0S7WZ+ZkiLe5yeu1fdADdZ
j4QI5mVtJ656MN2Szd+spXDZ2He9InsE09MOwNYHkgV/UBMwjkjX77Z5xVI/0NzjAwskUhDTQKt+
xpoDDAYmf/sGGbkhPivaJSl13p97YXVDrMw7mYYCwptEIdPYJx1u4safDcE+AhViZGTYkgXycfzM
p8A7EIiYHjq3SdLBi1TtdCe/My0LE9YExJJgEjOFfYS39DWTtW3danGkHk6Y49mEpHCrazbHDTIq
A6mNn8uyB7KYxGXvZ1CEhnQGl25mwUohhjloMKoduypmiSIMt3FGrHhrcG0aZvsssVpopBRsWEm6
mLZBF0jx8pLmJAYHGbE5XUEqOHO+pl5pBUm50QV2+G3AZT0sNWJceFyNOmXAZSNbiWle00wgdFJW
XyDEvuxhDDd5UOCFF+TsFs2i1ect1X9LIVw3FBP980fj3AW7z4Jd/fZXZfe8QM4LEmNCcxkbmwKY
sFwdXM8ElMf+JLJolzoELZxi61Rlhhdvl0D6icvDlX5Xz5ih8ddZ8ipyUnykDrU4lYPzF3Fm+NYJ
zCq/gUvnpBSShoVRqD4yH2YvB5We52a0GE+sS8/D/FlU02Pxwb0pHV9oZgFyRHPjCcQFqipkeZQ5
02wEa8JYM08e7KriX5WlS8x+nBXKfCjm5/lW1FMo1bn4WaUcyLWncUcg8nqImf4VuZrK6ELbsv7v
OG3ssa3edNDWFD9cbo8U72ZCN17aQbD+5ojO2/kTxR88g8A8sxM9DnjEaaN3gOnr/eXXHabTqY4O
ag687jzVbf6W7pzTbvj+Dpw130AjlDRwYoy4OynAdLmOPUuoKoop7EcH88oeMA+gyMaufufLO/AC
zf/x6RneIbVFpE5wm4VmsQH9Y+VxCvLAyp/8dUOK3VlJU1lFng3jF8FlJd6nUAvpMCUzQIVYG1Gy
BffWXzQn3V2kweMaZG/LgNkJN/yZhxM4sBzH1GwWTQ1zQx+B12gHkh9WsZwsybNNkPH0C2savFQv
LWqu4BgmSaTtrsyU/csG/qggRE/kmOdrPKEciL1eo3EvS5JOL/OZM9uAAwBwYmhncc6XsxTZd5ko
qKuW7v6KURCgCfR0fLfinyw/hOBhHGG7KesZCCQ96ZWyPHPEczIsacN1x/nYJANIhE6Yn/bFfdOU
bqn+ifnbsUMqraAGyPXJG7VyxsKGtS+IgWZVlEQNKGdhaSalfALxVHT0RGufgoLZychO8qQlN2FX
+fYShyZ7uL9tjxIBV9ALYCjcI0tVqHCjNxd1nVv0QKnDiiPCQFeUVPzmdJfSxgOjrsciNfJ+sheC
eZPxCo2Fvh29FNEGt2goRi6zhJvczFCgUROvX28lEwCAzjuCwmBWdyeco/Zn3TPd20LlnRiGUBsm
D4r/m46oJfLg9hqvqv/CVRp78Ql/e4dySSAZBv0f5J9+T92z7NRZ7FopXQaX74d0TxqrbJj0Wkke
jNE7D7QQqFi+RU+yluXZhR52b+uoTw/5UgpPyLulQfPQpGFTfdJGIN5C9+Dnv8Jt7xkcd3bcrBcI
hkob1F7Bi3CiT4oFHF3CurL/gT0OvE1ueuyimjFdMtoASaGH1hXq7RkOQ/Bu43Vj3EX5Qz6nQYOF
2UAfZBzEz+Yjxmn6MyMp55KRPEQlYycYhlwmaa+anvzpMCH9fz1GAh+M8gi36cxC0JFqidN/w+Xw
r4K/KjvLHVJzGq67ytEtlzD3iQM00ykSA3JCPTpdEUB1HXbXCPRBiRahdAeef+GUIAItthmpbaKQ
odglFMH6BVb3RQ3690yCGyDN3lU24b14mDMmMFnzGTWpNUsNE1dIQn7/Zh2Afp72/Kb+n1248gn7
VtZ29z2g5kCgwvRevzCWEmnINZvV4RaSPDZR0bR2kWa0a1OYw1NDpD3hZ2IeW2LI4ANwZS/g4A/g
eXBHGuQRbtJiMUDDMQw3Z2ycLq/5+WRDdKqIsWzc3+kX0vFQ/NdiDknw/QQKVQNOKUy1t6xxDdL3
LUnb9PSlbNsomJcC+xwyKwpcVUv/hblu5w06JzLknPHd+bbh8ssFvs64DH9ebpYIyrh/ycu2FMM0
ZZqFbG9ls5rMxpTVLaobiRvHvOWuZMR67Kp1tVa1zONX82zMH9fd8m+kuxhM0tQQtQ6NdfIRzzqi
rgG/oj7GH3gJ5x+Wowbm/+k+R7TOJEn/ABvJj7sn97jVYLpgSOPEGOLSJT3M1Vm+mh8rAQfutSZ7
clp1ekhXi0OiJRdu3E/EokUm/AyvEXDkCKmLxegjSr2TIxwosLijzpwSyi+w6ldLkkUP6LbKMliW
CSn1r5p1dA4hoesvDkD+H2Q7OaN28ixDSME1/dfI4bzHvtAC4OLD4olh0U1fIxJjA6vwTD3Q2lRf
Cs2p8+5gQexArjPkwranX9LBRpaA/hWH/qviSzcgOT/m8AWOEslxXqnHWGoEQjsxs++QsgnV28ZA
iVFxQiNV2Obo8SL/nPnjVIGVFZ/yDM8GzwLoI8hJckzJnXuE3kMCFEywm1cW/1DE59vqFXP5WVNj
9UNcMtWNtTIGfWE7nBMZKxj9mSJQoyYsQgKihmNvkN3jYymNwIYO6kV/MpHJHwj55BvvlFMkt/3t
AHH8MS5dUA8OQkK2HlvJduGrI8RE6+1v1y8VIpCkbBRK7Iv0cP+Rt3H+NH3N4L7TniHAqLOkb9np
Jbw1Bq0806WNFhr2wi7x6I1kw8sMKkG/NLxABFELuVHQDQB5at8YIDj96vPJy9ZMjk9m6vseOCVB
MRZzeGuY8TAujtc8aEQ+3ShpDb274KDHSUmdkPZuFebh+NcqGhvdWQ39sQ7vhPB017LeV1pVdUS7
S7Zw4eBdsx/6QDHgkwan8xoCVYraun7K0NFj07irPalrCIXGcpljaqongTllYnEwX8sv/R7OlxJo
MNau4n2L6Qrz1wKfYwrH4EXG0Sh/cz7VqIzh7V6oJd8IyN+FSQRBGVL4Iy2H1+wjghlFRHeOrPJD
s9XphPVswh3hqjRkAdGq7bfErJVhll1r7/GdozrKtf8Wg1CYoKndjOFQF39KkIFgw5rkfZu0dW96
eVjS9iu638l0lbyFY7JWpCQb5OBzhe+t6uz17uSEzvWlcHJwf8To8i4tOsG4sJCLQSA2drleOM6H
SAb7pb0IB/WyUJIpwUR6CIaiY9NeI36B5GNydJMRYPNMMrD7RDnQ2ju7OMEH6ehvvcwbZQEXN2jd
yusJu/l+m7Lc0B4F/uqokxKk+UCPbCQqtO27VSVfb297y4nUKfCqGorSsx9V9QaeN2aY7b1UuNux
Bi+yOcXTMAlExlOE5XriZeerqVEuz3WU5/GwEaclpvpf/pcxqHzTuUqlZItYwQGgzjqdFWs9g3ls
K6/mJT+oONJPuSWjqeHG9ASMDVtx+nfL5FUKQU7cmeJ+yDgX9cBOyV8UpYy52e1Xae9OoSoKn/Ch
o1PLWdn14sEpqRvPgXOFuBDIflDhD4OrXjwuW4UqzJbDQDFrY017vkbz+hHrtzUZX/oLmNVkLEfh
Cn3ImLTx5Zt3ySxKJr2BecdsvRT7v3QjiHXGAmboGbv34PJ0kxheYnUbeqCYGhygSjIElT0hLJhJ
n8OCa9W2W+Y/arSagwEr35dLJzPmI2G5Kgc/uymKeCG2tU4+8BYGRga69mhrgN6x5uUbq2IiVlhN
3gMRmh/roWrUiZO29NI8DsoeAZZ4VIVysJRInPhP4xEHhLQa4r5iyEIymBGvxFOthj+b+ilJfySn
nhI6SBwfiX5uHkqbQWhG/IqUSFSu3K9+BGyyMe1edu0FbaO9YzS8h1rlckc/x8dli6JRzZS3FEkU
C5epZGW4QPMHVL0Zdx4N87WuSpuazjgYH8OzR62oCapFEzFOAcvD4C4VHX1SPfds3rsPHpfXYFNn
5mjdLrgClOHrvS14C3vp5jsU3lmvrRrLXukwhBbHYG/4QhA17F7nY3ZxfT6X4kNY6b1gtpHcU0b+
m2BZ5CnkwnxpQAY1pw/65DDjZl/ElIr1Cf71GNIKUqBwLwV2aKpvWK6d5/w92f23uL2Xd9XjazqO
xT34bZyeM6vt6SBfpckXjBLfR9jsEKo+e2b5uVxH+yp6uqq2o8gCHD+KWfjmeGSy+K08t1S5VO8H
bVmNFqnmaJphKvUKH+brQPqkJXxN8nPRXWCyb6KoOVDoTl7SOmdpnrOOoNR/M2HW8zebHxQdz+Xm
+UIEr6mRJu6LvsNOKlmdD9+2MRtBg6gubKyy4hekRj+1s6ojbb7n3J8JnjaVKiL+gzmJlLbGEwfX
TEp65YUc3CE1H+wpubHwtnkyuqfuAZnnJUvDiydxHVZRi34YS0buWzjQK2/OzuDX0VQTz3jXVdmC
Y0RnuboIwHwKG7AniXnzTNRB5Y/jqm3FYBk9TFryQZDrOYcl3dQPODQj766QF+0zjD1w4KBVoRxg
4o8DL9tN7zqln/0SAcM0FPNKMA8Dxd/zbu+pTqlucAgu0ObHacqr88lUHfFqyjUOg0ynrGWL4+/N
rSs2/83KiAeij63C7zUeye+FzoXYO06ogkqXbtM/bwPEdZnCXwc+i+OhxBKkV9T0K/Qbt7gN8bC1
D38pm0/Fkp+lvM7Xu0AYdnWn5UK0SOrgYRHpaWcICg2B3vWB3FDgdwcJKrGybVbSFaN9w1O6Uxlx
QUvnXocTJtHMf1fYzjnUqXFA/2tfPomR5ByEU72HbhEbw7CYvP6YJVo0qVaqO5G0oPGtTOSARJUr
kXT3PhqktVje/e+4QlRinAxy0tVMMKBprai/RV/uR/hvDlrkTBE45ns+km6JDVVLOucATIYxybQU
D/0akK9qyRX1eGkOUrtFEPaBpUmgZ3rzA5LcwNLH3mPJedv9jLSaL3X80R/09TspSjBrm4GMe0/X
OiS0bvE8KoZeZq5UG2Ti57laWKa3IZAUS9DG1ft8tY22c/El3M4npbIk6pkFzIegwkxEQtLfR7ZW
SyE4EC+Ls+FENXpiYFl71jL0RX9bS+yuvbUcCcpep4xVMalGiKJ8DvhBfKCR/kwSh+cXSjCOMx30
hoAyJN5unAT7l84lEdv5a0YdUpaD269QiXGnJurVpt3zyQJOWmo5+5/AMVnx0Ot0/Aq39fv0qfKp
uioybYNjohVN0wqAgw5zT8vZlXiaNMn4BHOnFFqrRqcEISyhX06sDjTZEiC27X2oC6qxPK4lxXPN
sNvo/cjDxK2YdS0umR+xXlBLRGuyg5obaT/xKwx4vY+9cqcp56Lhnw0YFtBa27QTzf/5u6l+Tz4B
v62xxoOkSsfTtg5luFdamsV5H0TKxcozBYE/qHaCDd60V0mn0TpUdrbf4lYbyAYrK3qinNs4PSHA
s2DUXsDYgFh12FHffTV2pZsGlVx6WOmxAGo4DMaKeMiEeUj43t21uOu3ydy3QM6Y5a7JsRJwnScj
yxbg0QGyte3FX4z3EyLwvsM+PRNeEl07S4ZreDl7r+uqcI19iGvT3grTAPunL4wWbWMLmjWMF76B
tGz0+pyFj/qoVffgaU38LrWIcDE3+G9aZPUhoEhfHwzJTSOrWx9sF54KoTkPb6ReUOot/LRiJMg6
It5XIDHtaJGGkvGxULtGZF7Bv8uvx+MHBQx8muG40gm/4s/cJQpiAI1mG8BJl1wRaThHAgVtE1lw
3OhkjXBJGEe9NC4M1OvJby8S3mwRuVYzjyutUSjq9d+bTFjmQ5eO+4xChOHGmh8Z+9Jgq+GubOuC
k+xb4q44w091Uq2aXp44vcaL0i2vCXS9NR/I+jekdooxpYzpmffmLMX5Ziz6YZ6/dVao2jPQyk7d
rtq2q6pR8zz4aVa4KgRCrgjqjIDg3ki16cIwpuswOGAiWjnJRmCmsUEKtRJ2f58+p1choDpGGpVF
iaVOyBRqMcV+4nvcYH39VRLjUj1tah9VSX6C4KqxEVggf3E02qf3dCamM+YmHT6BzOgYfEe7h7uQ
Ui1D3Qe5IBVoKn4/47Dp2rGe01/BKgI8S69kvNJsJlO7goPrBuLanZMBoG4DcldbF9KpTZObO0NB
qvc3fM/KRflkp+lcDSWUhFemKnk0B023yIEh5qTavp3T5zjLJlHlaQCRXeVyFH/8QyMlX3tMX+rZ
ZXaARJhtMeEvaowOGS1/YqzQCELhNbSasJYgsNvSI0iQhuaXaz9/GrQDmB4URhr32V5D9SvBCc2X
N+CIrO1aWsHkcHqxbaLA9ewBlfEUN0jF4sRvv+TYyfTs56uc5Lmjwp4Gy2VtS4/FNIzjMqAnolq5
rlpa5WA8Msvb09P6iVMZ5GCbNJiXdmVG4sTx5ZsIuWUr6KICUwNqpGDsCK6OomORW+SdGF7s9yHA
IOJjNmedh4L9QL7rYMcg8LSuUe+W1qchxSEbjhltaricEy2TuZXhloCZhPxjqq7YoMeX6ab4E8QH
XaIwN1Us5W+o/CS1x0+Kp3A1qRNTweo4yN0SSxYteG5I2+JCGdu9+3hAJ7C3dVA6B+IU+FV4z/W0
lIhBXTUbCBn0nEQrVYBZ9ASGTFlBIIBAUH73ZaL2tfm64xBuuE/EtYJ2WM4Jz1GbA0gA+OI5BP+S
ZxRerSzy0SoWPcBys/Kkvgh5ECnJ3jcUqoFs4ftwAC8xrRhdkxQTQb4nQPb7J6Rci37QzYDYhYdw
zIAvwxwnC5hSXgxresasIxnagD6nJhehtem7k0GvhpfEMQHnoPJJI4cIuuRyTPSRhdbHuDMWkAcx
EVx0BnNE/TdGs8weldZINepNAO1DxMM8EyNO1UKcsQ4JbL/uVrs1nSWxtd//nsBbZKAByi2lsiGN
9/DoHybpDC1h/+eqv3lPmD7U3ITLFAFpIpBSzKEoYgGA8ssUri88R1a+of+QGCVkA/j9UGaihz7/
AojatrmXgJSJ8TaayxfQNDNLbVKK8vtYfghm1mDoVqkDgo3/+aNkMmt17HX80bsXxL5aH/269tPE
5UxWjoxrVwHsG1KC2qKAP7Wbn7KQwer/vdCkU89paqKmSY+2McORShpkPukr+WQvklaEo5af8FP+
IaZK5q7zmp0dqSsq7+QMOLXV3VGFPa0WNUljzFjQrL+kgok2EvYIoSaefQxm5HbSzuyupsTbm5Sv
nhBvGQZ91CDmpRIORypexPjD4X4PxqKiEfzm8BL5k7Z0qeAs1AdQ6x/pulbwLil8iWXCadR3JTAq
WqObYmEDF2GIDQtJVQzXMzcjoL9zY+dWPMt/itEZQ8aTEkvBqBXwYWRsbySkvnsnDsiOHy5KB+Q3
ZfVjbl+g+DyCurZ+XVLR37bwPGyacrn/ycFrwlcUWpeOrkf/GxOtmRntMbbiruSEw1Gt9/DlYqGl
sz2uYKzDjEfOj+FT/XpJMOjM7fahspa5oIYnd19eamaiyAq0V9A1BYEoG2GCi4hxP3iqaULSBMf2
d84191cC87Kr7/9cEQoqk2q6q9r1q1LzxyJ5VX2grLRsubVMGdK3N+KXENsvNg+JGmwvKjSiSFB1
DHlrl92lr78cMKyguhEAFSGAMKSJaoPFO44JXrgKJKEhNn/dVuJK5PSfNUimrfK+8Hs25rZAj14v
86I3a/TSrt8NYS+6pChxQO5GfGGMIlH2HQgmhy0D1f8DznMbuniaTMX+yV8Qk3wnUWUzFl1wfrK5
RlqZH+f6P6SzxnP2/R4PtSgc73okp2+3XKZrMlUTDbx4qcB12iPOGyTvf7LjhNzFICZzhlQCfD+2
KSYST3sLdrriYH+zBtK77hXK/frilNNXKHhjQeBzG19rX7oFjTCVbyMD5KNs+/CnluEXU7rq2wfx
BhujWgWif/lW7gkwocVmTlHKQppdlzMkjbauNCl0vN9KJOp8jtjhckaTnjT+fIoFL/KeRqYmevMG
aCkJEU3DWOa7eyw+Y26AFaj9vHJuq/yRNSMBfql6w8kMiKx/8B2ioKo6jVGqr0EgAXyR2SlvnMWw
pE5qt6TU1oTbCG7AgFpPJHAEhHGD31burH5vKCy6L/tqfnrw5IuyXYBOn6+PlUWzunHMmLvMAsQ3
FB/OzPz6chfMgXDrvPN6G36pXXwpELy76wrNWqnEQ9nbQyb1KQPaRf8VrGXvWyHUeivRupFB76mx
EcIsJIWbP0jhLMjg9WhWQXWC980RW0HGRvT/gEqe3bD6n5pbUnnrJHK3Grsb2xqWEtwhBruAjZHY
ievu5kKa/Qy4rKAfsxg2dAl79Q3cOaFiZv5vD72SOAcBVZgGLFOaRHl5xWVXhG7ubibiG8C6XzOS
j6Q/A7cyYVHylcA9z0i/5DVW/vVAqRBTf/a7uKOHdil5RDwHNNP+2Sm/QhZ8K0wUTo784JjHwlAl
oGh0/fZh0VjLS8jPQJLI5//mtxCWVx5+US7s61Lr+SFGXXCeJrMH0St9qeDlXAX+szcSGpezIYsJ
No4pLDmXchlOSGd0gUTG9bBj76JvCBZFDmi51b61uyDCUJXKAMIMIkGX4oEHnjyxrymoVbFeSRDX
zBA9ggY3xn9PKBqFxSMbsRIrycVQpkOfzmJRIZtcFRP98OLpIDWyCVzpMf1N7K5Z9WCIXuqIjZK2
hVf87ta+VqI50ltjhCMJwTUS5i58XfgIBPMkQf+yJ1GZDveffPddHDI1xXPGga+W5jY1kCWg82ds
G25wD5ijoskW9s+Xq36MUCARuNtkoyogccHDU4H9RZibR/0QhwW1xM2fLT8EawY7gM/uQUrAHwIf
zCurUJy0r7iEdRGpWxrzyyVBFPxCA5nfb83MUTkVTIt+KbbGRBuIfDU6qjgK9PVTuhpfhOA7WUnI
B3xY+vfP5WeW7GWUVm+sgLH24VY16gV0VlFZbfN8XMteGJtnW1ucNaa3m2w3OlD8ZpvE+CZMdVzx
hHIobeGs8UErMRHJwbXd8gRTTaIqf5WWJ17ch6+PRZA94r3WoS9Zy/nt6RkqVTEoK6r7Jt1FUhBL
vUTeUDQU1w3hop99at+pLgQJQvXbOTYxrcy+BPWCR6vBG1PT2kI2/aObkpnu7RmH5bh8/a61Fy84
VV/SMm29ZZ7YM5OnAw3ftX26VIrH8wSkp2+17xw+gqnecoUYV0B6owLNzQc39xnLlndsc3daKhXf
pemXV/ZIG2/D9j2IDDeB62AZ5KYg7wpVgvZVMk8z/vjrdK/QRsK0UYVZwQXlWXER2136A/OQLDM+
PWdzz6ba9zUoh4Aic3N44b1T5g2T7NDXZyRE7ceDVTezAj7c4D8X8QH8fLDuZI4rJqQ2PwE66VRT
ULiSnu0v+TQli3I0fZ2YRRtYxevkD+5tkUj1KR4e8iRNGc22bvDZbJYS0HHUCR/3lCBtRMkdEK/i
2x0CdU50feLGzeYsYgSz9z2BKqFsmgL95wn8poswcjMUSzoMdYZNwA7zAdog52qeP/VjeZC8+eVb
Wy3dIEmS9CsxxmEBVm59hHRrntM3DLPK1qv1nWS3a6UHtnd4E4o1WrBTz31dun25uwLZzwA7rL9o
lqySFxwrFh6whq4NqFE53a6rx3vCqtiLKECOEKZ9vIDTLXyYGGvs8jsY2CvE3xpOKMHW8NryvwBj
vzJxWX2i2oqBOIc/ZxIzDZHrm2MUDEsO8QiMDmOjMkF4W5qCHxl1Wjve0VtjpfSrkf4pJOE8OF8/
SPJtmDRjAleiRrDGFX0tK3NfOlLJ/7/wvSZ6ZQtFnukousr7yJPaX3oTZavEs1v+VuAVvhv4ejDo
kkxDz7P0/unx8KgqlO4lL9uwm8j9dZnQE1R/+22g4ayvZznOV4JgSNFjrj4hkdM64gioW+ERAiWO
1MHc/ZjeDsHhugKYSvZHUfa9xJYI1x7knNxxnhqI43uivX8a2FbGOyxtK8v58PVc/DWY4tR9maZm
OiliKFQPIvjpQC1NTBOpxNi2ZqMoW+ZT8ApEbmcZ3p8GqZlVkT3AlersEwJFNuqZsTG6VPXDIXEb
JWYZ+OvJl83GEnQ3CI8Gw7SPPMPjI73iufQcDhjzLS5+40dSPi9eARw+XY+OTVXpvhnTj/Ti7tVA
ZubyGBTLEV6jDHN4vrO05lfFSrzTPLUUOLA6J0YwRVB9+6Fiv1qkUKvDlHRQW53lDEQpXW54M93k
mW81c8e7w3ScbJQTwg8VQe7c9xbF6nuYsbjDYURa2gEF61RoO7Itr1W0+lA42ThJyoibdf3LCiBM
IFRnFetT9U3+95UlFbiM6WDUVW4OYu5dmOh6mF6OrlLSiWzdEA+PdbNYbMN/AdJzZEUR6hUmXPZN
3xdy1wK3xev+5Ug4i7d/9t1t7vwu9J2IXBRVhwl/5QP5sUEsWRiv4BkuQJV7kvZWQ0UQABENQnPv
zlSMkRrwbELZwiR0bBCikk0F6GEmBNE9eRtZvQ2kyb0OeaR4JIFm+AiWoaYwR+dIVSI2n15yeOTF
ZpS8miImVZxm8JNdlS6BC5mUewkJcZalzN3JeocWxYBUutIMoC4l+AeI03Ppsie7XNJxxmas+7s5
s6t2bOwJS/vWVrGRbVJh4RQDRC7HgeAJboARSiML52Uy2gOYRrwmLMuUPaKvKI0C1fZjnVa3x8Dj
qADDLOkYPhdCzw9O5mCbSZXqMByeiz8UysiPeUcMhs19hmepg/X19VD0rdOcIZKiJ9jzykso3JOC
E+l45YIyS0kdNKqArYo2de/LaF7wQXeUrSLyBL9sIRDqOEXrMGD+gjfeQ5vagTMSrHx5LGI9hc51
ObQRVAxiHCu9owk8ta9cksJ8cpeeE7QcoJs+c+zArtoSiG9E0Stj7ZvPbFyhFCXZUDh8f8hAca+c
PNPNG/c/mzxCr2CxuexbTixKNeDe+L6XQ08QwV9m6KmvO5eVjzd1EJwcBz6N1+Pg0DVLFmXenhsH
61qtGyD9dZll7itnnTQ+7wYvSi9Y2i5qxDIDwLsRIWv/+i89opXdBiEOvw0ScuDwfW3l7TT7NRmT
uHs3CVqM5UNov3WqwSAOW/NCh83ZEV1KQ6atGGxRpV+THgoYCl+wPVbD0u027SlC0rDjTBP928QK
ZCcVhU2+uJ2/eIf8ojKmE3C8fBBJL6wdtsRL45BXQcv5RhAlycS0lEPNJ/B0jEeelnv3BII7tuEc
PFOsbRDiCbuWwyM+kHnH2DHuaXUzWkQ/3+akX7Dr4J4Imh06NPGMiFS53ni559iwc+Z0+CqlLP0I
cjGvwVXnDqaEJqfwsIJUQ8qwGdBf7xIo5Icwdn84HAtKjIoPiGuEw5p6OEeHhoqqcYeU0EG0jbNY
NfUHF/qeANfGj/CDvCP5aawVLXjaB+ifi9tNDwpMclf7QXAvWkz/yDLpi9519PXqs1VPs8BR38yT
+/3GF+loTc5UFgifFwceLnp4FZ88pnd/mbxnOA7FW0HN9nOMZW81g0khwU3qBYjdRsSY5+aZwwBh
q+CM49iWnpGVDLFzDz/U9qyl3lpt/+cNbOJPSvd6ro0IkJepjVLJHGh/+NMiW32XIdXU/9+oFpG/
gHukgBv0jmR+N4W3uscvLnYmlfkUtJAoHMwIOUpppZldc6zbPvr5a8pmC24uaEFObfdP7dFUjZJZ
2M+J1xQbZ+QXaDRAA1YaXDEliu4xkyAPY/xHJ/idokIFCtFKfh/vcpcRba9dA6hbeQ71dHKM6FmJ
AZyQqCVsgIHJUF1ciILnqpk+uZ3Nh3W0PMk8uJePsPVSAl8huC51vZsDJc2IjsvODw+ppeGMqV3S
ygjZBy33tAWwEbPhxACPQQku0s7rhS7pF80jeZHfiNOzxJ7vzG+FbjS5UtHz5jZ6FcBY4O5gSPjD
56xSMI9oFx1eiGhW0DpNcioufjS+zOsaDGGT17ngV5ypYY0WOkhpEPy/X3E8hHQfoCyCHJSnx0Y5
hDilYcIFJrhhVOrHK71XBADsa/ZXB2GzljHgIConeFIIut4gKvEFiLGc/H5qSrfI6MktlttsXKZi
/FH7QOeqgEFtCAYwbzuvzZUECavt6OJLq0yVg2JDwxdqW03fe/LNpT5dAwTqeBnN5ldWhcK+sWPj
07rmNuw+3UOK/k05drvIuPf2mECRX6rQybC5sbtJk4nyJKbyaturV7Rrawj/bZvkGuyin001Zsve
raZZxLM9NUGIbknqWFR6ihGFwRyJnn7OCs0N9T4XUFTnkC8BYqCOqakzTVx+h813bUXn/dLiNjAB
/KcuO1WWc3g2oX/yP5aCRf11KuquNSSEmT1Z9/IyLr3gK8mkZFAAJ+fieVN0tA0umjYB1zowcuFR
wQ8SdwYj30eygkKbewBcBgX15x9IHM2mrN2d4Ljth6VLmaD56HyDT8vnxpQ+iApI6agBaYZHXtCe
K/W20/Rw/QsNwvJKmoksIVYS5o510pj7m7h3ZA4LH7iHrIwqUE/Qd6OtkcJM/R/wdpULjPhUsx9i
g/uY1IPiccpkWzDES8P2sTzbAM15C+XpgWE2aJnxHjIXs8kFu3FDxfnW4xviiMXAQs3LkoubCtL3
KSIpp+5x4XYgt3OcEWtClfMcxs1orkURyVpSZutufMVdPVnLAmOSjwlMXK9FBjQLtmXuke7eLzQc
rcw4ztIntQHAYQTD7tlD9ZF8oxU0MqwQ64jD3hzESjR3nDFLxMjy9eeyG6dukqR/22OCTKuwc2+U
V6ecE269DSEcfLlhYGfYi8RRzWFkebCYq0QYvYYF0Gd69IrGH9d7xo1Z803bX0/SyKHMCHHzx6in
q1N/7SuHjt/dvMg+Na2N8Gpb+R5EsaAQfz7hLRz5kld7ikNq9+4X3vwum9edXzve7VUm1lD40j1+
r7lIlZsiYBlZNtdqAUzKs5DPR0JGLa/KPk3GBD4zCZUOA1rqQkc3xjUOQqCuXVm7YZjw3g/i8fgD
ggb1hMyYh6NWN0crRhFrWVR1lXWw6+NqEYdVZOc6wo35u8IjebF3CHB/KX9yr9knQXqpIKYuDht4
aAa7nMWW8OpG7VzQ3NaYf6ZXDNXho+7pAWlxx8npNEhsnSmByJg5HxAgQ6KvOHIMajhIW9oAwtG6
s5Yr/GFW7QMaU/GG1lqbdu+MYWjnaCDLAatiF0+L2FBM0dv5px7WUivhkso5Gosi/4RyBit9AhG5
Mk1MFBxI6qyg4W9sIlLwoH46n8hY613ZCNEV3TIRRxV+SgQRzDk9mNDVejp5MHLN3nO/fDmHyGEb
cdCat827fyJhmHHBU8hRqMbGJI8XMJS6MdtzUn3+fNFCspLjV1E9sqBH9NOmQosV8XkGEVee7jHU
YUmW+D0NePH/R75Ki3+neNIgWz7Pk8+RA8hTwHOaBbBOhlkamp/+dZX0qKhUw5vRGWl7Uzig0Wfj
JMhvPJaYRqCB2HNza47SmBekNf6DD4SBPtLkl4iO2lAUygJDNBjA14mp1pXfMdiHOAXwcobS0tlw
r35z/9yjAIbxyzQ780yAw9YoDzkfCAUwn9E9/daDSLl0LJHW1Df8ftHXdI+cRDNVHYReidfjcWqC
ZkeSSnkYUvc23PRqcy4uHSk6HU5Sx6RiO+/pMfyc4JX9K9WbdGCEIXVch6YPaIV0F0HBh/F2fUTB
MiZ5NDxngrBjof2it/xNBFMP9fvitHl+AY55l+ecgKAO7Makkq6OlwXcXouuEtPZVQeMdpP/jqBm
5BVzeJZfHXRIIMQ7uQsHjRnjhZvqHyrRh/YIC8NXXhsf3A3wcjVKCgcnK8mhLzB1lZ5kTWlKeGgq
vWE7EwvBEtccNxoWsPRMYnqH+/QM/+stziMuS0TmppgVyPcVdCtfB7a9u04EApLT/hVD5974Pa/1
liDzWRROK/VN0peluORKjBuh14d5TNn86jpaCGU1f+duoj3k5UHkbgsNlSJ9Xj8ZdtJyDDSD/36Q
RvaMInhO2QW9Hhkgrg9LcKNR5Mke5E5XMSbjvwI16jIhM7vEGvvjYw4FGi9CojYikb7ESmF72tg+
PQ4KOrYzLxEpQpZAyv288yePDLOGfEehFP4n7yaPTbxxCqz7PLSs4wbP/Z9aMLyjMnJV/nJyMRdu
HMoTEi4uT8XgbIlkj2RQ3TdkbGDHGi+8RFzEzPd3mgKx/sEVj/jnImb5cq2bLgLHqRykaBAcLvps
MULPDHxoplVZOU36Hjkf9HDLr1VzE5T1s/xoJaVtAD2OIT32sTgBlk2CumA6ZPN4944I5rEWXyvd
u2q4kNhyjlV7GvJgQehtNdUgGd9Oxe8D9GmavOy0tBMwbKQKjZkSGce2WuTKEK6ooejZeC+Z/cAH
QgE9wi9YxRbf6xqTrKDmHNRgvCe/eWjiOkCuBC9hBiNQkuUhZ55W9paZd92OKtuwsMpRYZW9FPBi
k1DbXsCR54hFHpNGTS/ju2/jgOXiRg8p1TADAaPaCGXKsw2E0Bk/gUkOEKAnpaBJj6azFq4niXHX
AOPvnOc4kC1nLo6kpszHxRd9EAEkeHmBxi3wdb9ZYcDRPfSP27fLellc3eKPimp8ZF/vJS5ERsAm
4a4d0TAbYaliUt1rxeo2yGGK+8+7F0VpyDeSA4sHj+ALR6U+rDt+VRPBs+Qgng/3yac6Szc9N3X3
VBx0Ea0e+tJ1EpCP8yFp4Cix7tL9RBjK3Z41UMBJPezl1KAlTgKbL+7KkyOaGDZaS/K9GtVXjnVN
w/EgrI/y7XNrIlm0lBl2e9iDQ0xJ2o5dsNqbgts/73TD3lan+cz7MOnGlKzTMfcEGroJpwO3SIEK
sNXIvS9WGoAyuO11xNYbxcWaIb5uU5+QhZds43NP3jlDic51lG1QWzT8QKHjE3FQIo3iWfM5mywd
/nb6KVpJqifkyuhsuTFv4INg2C8xft5f7umr4V78w/aTai7IDTpdOK1uo1g3T3PBN13Z8xhNX3hX
jPk6YdwG7XYqTWqGbloktjhOFeTtwdZGvQSAvna3OFgDS/Cu2kLb+PAmjGAY772GDO16sNRL64EC
Mnwced/OoRl64JxtxxkI4THg6sP2hy/IYRpxQv0YUhoDHLnG03iJTb/07wrRA0h850y8MD6CrySK
pJ2mk3gv/bbZTx7jM7wq3KQECIjmcViyH8pGQL1n3Ux6wR2jkhxFX4IyUqXN7kMsMj5XN3BXBp8d
NA/WtTQViquXgZSeS7I2Jlzim4tbtV77tU1zp6YYLqp0o+wlYQt8ALAKpIswXuhXAJC6R/sAfjYN
jNBmclq+Xx0zw7awn/GecbbS9P0Ni0l6hk4Vpck7WCoLHJkfSEn1/m9i2VoBpStSiZxWeQmkns/Y
oYMvLQ4Zsj92o2Y27rsjF1QHuS77KJ87MamPOptTL0wajR5Eaj00/UfKGFdVsxeAzZnen/Mv9EnZ
xS491ENkOHZEclXEuGHDzEAPYF2W++XX1QYO6ISneACzoJ6KFTFG3wP6+Upr9UBOlffRBmReYNMD
udVKkxedsDgfqMNKFQnDbNR/N+klJ9hzHXoHyxUKe9YdlJUMBPfP3EQ/ohee0u5VQh5kP5RU1PA0
rncGhKUKw3PN54HDomO67kUyDnp229jO9PRGFzfPLQsHu1/3YECRT6X0iS709rirZWWPgOucPTyO
/C0HJqO6eXz+raecf2DSK1JY1zL6zwsB8sPeAsUlvLAmnb5jHgB254WLTvoIucyUXT9dPh4QX/gg
bUw4b46ENdAHl6enX/c4G+cHAN/XeCJuLIjdxHTHLCvpGrH5Y4ohrl0gG4z6ku1tD9t4jZ7M7AnO
bpf464Ez2ytoFdx0axG6pPMHvjH1jV23UriTJ6vg6slqfbfzbvHltY6p5hBqFOUIdcKpizq9bY+R
FnnvjQ03A+djWTH9U800xtGiwGrPDsspPcpJ/+Ttt79D6e+B12lSgBzeQiIKZoD+Jm3DO2UY618O
2itmy8W6Vx2gXjCDrGowZY7Z/c5HQXrWu8B5EIltI02HO3YcAq+04l4YXIpI5eS65722gjtEk7Zm
dGziJe7yQI9Jkz42ZFEYOy6QfFd6vs6oeEYq+yf6DInVnWXE+zepFrwRkekCZRraHm2LGrdS+Tgx
HkML5UFC2ypANyM3G619Xsh8A88TWXksnkV59uHrQPl6Oaydou7YhB4yhGXpxLEcjF4eC9ZdUcCV
M0DO/kbsLZbb/iHeev6vNkhvD/AhqOxLyt2cMxD2ocDLPShp32nTmL2v8zibeAxReITi6yuTAx2E
b6pZDg91vq9+8ePL9K/Fct5+s6PYDoD7CsPXBSwegUfAoQyHR08vDol+et6i8hcdhO+xQHa+hIZy
yEkS8q6WnOvP0lrEfeSSZHK4ayj/ohtkl6o3W/uzakSN1/0kE4X/w3PeN2Wws+vkrX/wp7cV1GBN
HJqX6RRYgDJwfU4Tl+LHXBCnvtevLGzutY3MJkw+0xrjouKWo/RWha6RlZ2qHoqLBBBfZ1cqXUQc
mPE25mgt5dXAu+sFXewCqEqjkaPtr7JjX1Gv0dksBwJhsuWWkklsiKQly1uN9EVm0RW+tYYp3cSE
frA8UelK16qtyMdppuAt/FqbB7KPE4D+PmWAJleCpNZDBUDiqMv06u5nn1M1pgYViKm3nwPGLF4v
FeJwTg4zl2HujsL2soDKzBM3Z7lQVRxWr5Ksq7LMa37eQAZL33fMEF9it09Q0QtwTOuoo0R3laVR
26uDY9Lxh9N6SOyoscUvNY3AAk7kgSjDMuAYNCUv6Lbfgq6vyxuQWIhQ/FXk262bdlw1Dhnbw4s3
whIvXd7gCVBNFa2ON66rjYDSZwY1O2jQki7PYMSDQNJaTvHdvewkrc8iAGMlvepeIGPTkvbb6rgt
LN82HQmbdgI63+Y6o/SWLbmDRbNzqX2A2R7/mls1k+9oZ2BW6zHOQCgiFYaTtsrrAT+lAds5KG1W
IJhsz33nRC4u5VlP7uir7b1Ca1ZVaUqRI9ckRtH2tv0FrRg8S2yNLNX+Eq2C1VRGM9HVtzYpkUDu
630Fmz19LacVW7X191Rd+Fuq06pUN+I8xdM4IPKOdnSV7zSRu/BCekGVPfQ+Xwu2vjPvODhe7JsY
2ZOjLBkGLkARTdpz6vrQHFn1zAz3z72DO5H8G3SY4FR4+vcAYsFwLsCt07DPVQnsu62IIpmu7+Y7
Cf/NAUK6KH0K2s9Kjzq9tX1ep80arxs8c762tthGZZ3bD8vKyNVdqI+mt9XIJ2FKQsiotmvpXuQy
fMRl7C1vN6rIpQ3EfPZAQDJ/nRxbO7hlsQIk5OkTdP1pKJhNC0fDXYOOLigmi4mSgRogojQAgj39
emK8OnivLLobqNYngj/7AgprKrbgDCBu4ycjr97v6pyz9mTlO51xavJSp7vRabDE3WodREifhtRw
Ns2rXLMmqUGK9FQqYgKZhF+0f8KQYnj7scgIUnr65sOSDYdIL2l90YF4NnL3D6hFbXUXXqGNiuF4
vTd0T5kaXv5Nu8BZndT8qogLojfWzw/MjsBmt+mpMKeSWrtg0Xs0Ovn6JQ9/pFUA+Km56SF+Co/q
SZZLat6e4SRd6pyW90s5R74ZLUVylw7JAlvcGf/9pk7LNQfRhuTMMSHixEZ5FlKwzwjqEyL+mhz0
ORbNgbN5bd/+ovZkWwo4XHrFBwoPEgpFzgQ1IeKIAF7uIgimVxxyEjoeKJJorA0bwnmJdM3V8XlC
XGivbsD/E6tR7LR9GO5HuYdcUTHT1GMPDL4/K5tGa+KKt5qlBl4+A7FqpPiVMCu3MSl6b62RXsY1
WMo9lxSHoHom3Vtq5enKdmNYDP2jztup8b/GeYp2+lIH98y98LdoedbEDabiiYogkm+JWBm2RnQV
3CMdWZGzSTcjUVGfOp9S2X3PQWoNwKw+nm1Lln4Tv4zFHQYB75JkVm/ewmdOySp/aEn57RNjOBsh
wLfxCVsSJy2qHrHiQ7RBZ+uJ40tO4gvjFDHy2UzvghrrRT+QLWoV2o47hdiTimgTg2ENn7Xd5Oh8
keFAOQpZW3eCF/mK+Y8tebvWClom5d9q151EcBP9TcnXLK/771cL4YMXcZ1v8vW5HaQ05J1foOAs
1vFoEL8Y1PrLz68URlK3bcxzaAyZE8SOv7UgRNtvCEJtUv+QpEDa/ygS1s23oWPYylFSsL01W69r
T/28mup7gKqyLvXJPfU+u142CLKuGwA/oRngceRmO5AyKnrFur7iQZm0DixCpZ5LYoIwcINyfF52
0UWoyt0ekcVYHwhnpLA4LuugythLhaX+oRUH1xU3NWqrx0WVdY/ERXP91x/B9ct/jESqepr4Qu9Z
RFdY1xhmHwF0I1dQ2szraXizra/Nwnh+pvzomqYUkyS05qgI3xqDpaZtzIqhHnK40yA2MaC8uEyi
7stBnVBkLBAskYnC0Sggq0DDwbyMKW2/npTdpqFKtGZYTKDf2lUiweW3DXiJQz1g+WY+IjMgIaY5
jyiTk5lfUuPU/C88Mw9cm1r7mbfkt/h08wyaEMpXNOUMlngsWZdfpnTnpLaSZg5a/B9IDQQQFdKS
Xb68ufVLSbAO+5cbdJAxSfpxfX96hWq5evFStdaPmZiDMqSGfWEQzC/nT9qQ9yU8HAX6I5qODbmA
5SnyquydxcZABp/okRoSkiLsxSIkpNmqYCrC4lhwAV5nWsXUncqfgi22PKWfBiQy3WGCknra/SWL
GzRLADkO0k9ExiTPTry0JK2ymK2AKH6l8Gi785rwxyOekd7cxU12FKONR7et2qF82cQVzfWLy+hC
SdeWpPL2Un6kw4eOHA6owayDd30dgh8diy40jSExg0WYBCl7uE5Abj1oq148rro8+nsj4qWZmap4
SqY9l2TzzL+/jAgzrXOYS8d8EYSWh9QNVW188blEhOkU2sJwnJIPAQHyBQRDxxLWrq3wyP//+Qcl
tZfMZeSRLVNdif3Eg1USUXZtUU0SnIVYW4lGdJD2eE9FvXgOXV8OnLwQ3AX9+k22LyWeQGu1dyxb
blTXNMgsM2gAFWCHQ3uq4dvfVeu02xS9WUx9iEb7GvDSOTcGc8QceVJ1sVtTvLrbmm1Bek/LdR/M
spgb0f6fhPfOj6GMDIN/IkIG3FypcM9/W2pnYIIkJ9a6zcjhbU6+3+xupFb+2qFD4yskIdYu+Lne
yd+8TKSVbPbXoRkd1fnAqxElg5ZJMNtR7m+A0CoejeTvuFTMcO2Pku3FeshECUhNojYkTSSKUQHv
xBVIfdzPtVWjgnWDz1vgjHW+YN+Qxsphlb/L6Fcz3YIydoFv94/8ymbcrO9Sewf07XkoD3BtLZ1x
TmcuohC/ajJpX9VafFNWFXu70VufGzohvSM6BUWOuLSeQxT4i9rHEOka2sIbTkawlFWobHqmDDRW
tevgbQDSBet2h2sT1gt5+Rs0G6VPk+sdhM8wmxH81p+77Uqi+BjFa7U1wxtN96KwBZoFHnuyJToe
LWteEnwHplmooUX7bH4xMwZP7p0LqRztBxcOIYS16hCUR2mya2ZZUbxfglr/Jd9aBY45lPWftbto
JBbzRBqkQOXOLdazD/RCpPKmkkl+xLBKMZLA2v3gMuXY5orn/tIJkhw2cTsx6USXfkEbI1YxAfd/
T2tP7IBAtW3a5VDLJh1Wo7AMj4m7aLdqfnyWUfiTEMPMuePrESSG45YMnTumG8zA9uYQdffcXOmr
1IGfpr1wnBVvQmL2IqiQyxDSJnuZK+rT0I9NRGd//rp7zapf4/rKtBLaeZrFhsSNfUfiIa3Wu0ae
Z7HQfpr7WK0sSfLo25zYXpLmEJVocRO7Yq++AuFLm2yfnAsIfkT8641xVccv33KTJaymsxn+4pC3
9LLJ0EvewdJfoKC2gqE3w2AXVs9aLi4mXE0LC2F+jfO8wD7Z2WnGwz92tqGcPd6Fbx8dxl4m+y2h
6hdsQNvEc6MxZvCwAsZHY5b2tdEF51Ul5Kar3zm7+2yqkH8zI3xhsULtFekkswjn4UeL62/bE2qK
vuaF4iRWYHNzA9seM1L9oYI91lOiz3U3RYbUaqDgCwCLceTg747Fz444F5IuJpeTKAI58ffELW82
OeL6C5qRiscTqGMS7e1O7QBPk9qDYblEWcmI9OWaUFgRH3H8O4TLMIADakKKSH7u1LCgQcjPehrK
lSXpV5CEMQ3bu8VsxNqqIv1pRS/2jUdOhZBZz46jPcYTvirjkH0lM17rs4wvlmKg/52xAAidGnez
q2OWmVkG2G4YxTgQLOhn4I4eNKKUL/N9kZ+Ydj+S13sSLj18BAabOVW7yAV3wj7jWNzOa6n/hYAo
ZhM2bZ8iUF7tYjI0uMBU2voCDSVLqro6ZUm8Dz5JxiyBv6pg0QN8t5Sb9ci4OLj6atfGtVwlJmUL
oUdD2/7CRV34pWZ9rvHtW3Zqz9vtHWyjbyBPULLx2uS9uyww6yBltzA6TesSKcX2/+kx6+8wmUvy
zQgqfnQCCYNUayePWZUTeZka8NYr3aDXz5n6OrB/taLkzbMMcfgjnDmT+3HTMO3HZN0Ks1YtQ6Mz
PBNA43bZ+VagcUlvrZHvBVqqteMkzPqkuu7KM0myvelvbjR6b/NPi/ypPf8soj57prLKRmqDdQur
aHk+UmlWVPAL3+RXSLnBeMrwsEKx9tMoe0rPYvN3somFmxXm6Gn4VbVXZcSH0Dv8CjFrSoCSbzp4
tKPkpnn4x/oxsbcaKNNMWyI344B0SiChTxeUn1J1rCDe20lm4I+cRPinUqR7lY3p8f9TUhbF6Rkt
2+A5Fo1qmvsrbD5Pslz5orjEcspjn8Xz3c9m1iTzGtiNgyrhQt3W1+wo1PvdcpWo62cwY6ZzwDSl
ORwm0vFCVxlDsAEweTGDNpcWIg48PD5qK/ICH9BwBG2Ia1kKI26u3quFC51pooIxIrWNUNMli/ed
wb4aIx5sFXU3rA9OdQ5NYK8oXvtnjmPGUy493uT9L/QKL0kpnp0dKXPDMwmyB5//rh1gQqzt/rS/
qXis7r52fSNQRGdMByP9DYMB+i5qvZOBRbazyTj1tZpeswu+YixK1khyerhVMtCFnSbTbPE4WJpD
sTjiQMjhoFc26H+r8niQrYunW3cit4Fh4SjaZvhE1zT41qocGw0HQoW9ulWJkWWZ/dkXPJ644uD5
ttsgObvlKghCfw7sNg4WyP102cZuHr0613egBjt0u8kAjpoXlZtIjM96OIXzP//fHoTWH1LySdEM
ipdPVwAKxY5G5cwtQBakcPDOF4mfyzeBoRrIDw1h6KMBAyXqPKm8gtZurEzuzKGQW3p9zH2sGTnN
Bq+hrsk6oYpsvhgO87lTNV5fQhypQ5yl0LyHWSdrWzk1MFh/x+0jtwhmwZbdfloHibZKN+s8tss3
SkwErP48E5WPneyuqCD9UdC8KZGEwkRDVtgliegZsfv8Yc9BsBUAMvaq3CzUR9CLFuqhFv8s3XJH
DFtf4y5FBAZx2gAo5vb0+l2HFR8Q4Ds5QUHtcarVQ2rmjvlgDBtlrexMQBHWMEadm28IqbwkUoXo
smzgP+k4+icoS2CNTDOjZEn4actuqudpL/k3bMCGm96moZp21JGGhfiDysXNbV5bovNAx4J6NB9W
Tut/VRnyLwlaxg263HH1Mh4ajukM7TnMbs8dx3HjS9ZVEc0dsizgpK1xphi30bNItVyfC6UqSk/l
RpHrVNmgasqMEMjZqq5My0xoHzc7IWGmrpL3l+EJcefyOk1nwnjT+tDhsFAD0SvjWw2XwgMZ7y2S
LhCJ2p1NAHAhNLCbBvI8qKthHcvZedz8Fdc5+T4jXpQUMElDLqlIohIxNzoRQG1E8WCH8xqhEoS2
KlannUI0eqeR+OfroTR4ovmD7b0+SdiRx7AahPFbHYExla7T2JksBjBmN57dhpQ4+mrC/y1X3Hh5
wZOqLWl+zG0JISJ3oXPI0W2o9s6yV+ugnHEzXifFpUFfBL1UcELOzkoGKeYEBZdtHtmTyVrePOfV
bxIP8YiKR7xlZXS3Ewr4V/upYpoQWdnNoLvdQJW4I9FP7IJ0D7Tn8J6VX0JDV7KqvufjdDCvzlxq
jRbTXdPXMZnlyDqpyPMLMFwDxhTJ3+2wk2mfMXeoulRjqRPT578kNKmQb5HNLtnqfMe+UP6YWGwb
qlLzs2TF/aNenx7mS1v7OBdblfMjSzhy/0yq9gD0C5BZigfuMWEjYGTFbdLs6ihLYmNpm0w1TmTx
ddDlTya9hHKVgF/qXwTOr8dnOnTP8eVXFL7RffBi0qqEKb5cPcD0ZMO8sO9j812VIfN++PSRZca+
h06vWVIw5a/UyM0mE/LuMzPiseBoyg60qKfuYeQ2zFvtj/rt6Nm2jhauHV62ugd5P3Fb8toxQVmg
w/0w2AfHPyFJjbOtRkc9fhhyEkzZ0oX7jCtGtJxN4RcC1VBURopRg9GQRcPmkfa9GcJ1AnNX+Zzo
yqWdFDp7Ax4AWzYFEVxTM4kR7EyVhMja4lxVmcJvCWCvxN2yTP++dLwdXAgmaSA1bZlL9azW6MUX
9kq6Qsxy3mgbzagJjFbMIDe0ZhsMSY8hSOC57EFlty/MJX96R4WzNmNGupBqz4rpygZq6Czq/Q5h
yR8/G7wTBEmsPz3O+xA+4kE07axDJ0XBgX6VC4vLfAxEaGodA58XOW+MSP49Xn9P4qDlqbbYhtdS
oRY5xReWt9TfEPd9vDBohEdCJ10QzSzt+BuBH6lzx5/kwAP4DxHY6hnZ+CkquhS1lNE7LwiF/0D/
3rZeLfbIDctMpbFnNrsn3tpaIL0qr5VVwCDs4i8wmYska+k98dsTEaQnA4aJg4CZmVEEtiM43ph4
z2qFUCdcB61+Y8r8kU42cFU775RpPo1g6WXcFZ09FLBtTD9MnlDqVMlcnsDJTQADVXa9BWO0J7uP
Yj1kU4Zq2uad9PaAau0uJHDGU6xh7bgBBKL2NRN4AgAoFhRbcTR5tJbJE/Mczkg9Fx7b4sGAaPAu
GbEhE4IqkvMzER8npBqMYmDjwGDhN9+FUI/9zY2FtbzTnQOKfGw3GWtrfd6JKzj8TDzF/sGtOw9p
Q6eD7JKIsJo6FxW/QYKvVLQUu61widTHtnpFHavQk5Sa2Hsl3a+9O7ZrEaD0T8E5arAPp/mX36kk
S2qXRYqknjixMUriQ11aBCVfPd59EQTw3ewMPe+URwDrFlwiAtqSgSfaW2lyhyMwFi4DVRDlpCqn
vzKEbqLSCp1bg3/KcS9X7vpP8c4AMJBFzcCa6yoGxBEF4M6zjuxvZd+4gb2WmfHGMk3vgywaKXk/
vmZ5WY6QG5vQicviKcxXVSu8vHtS+4v6aN4DtaW3yTyjJBPyBoUFnI3mQgiLO+hi6whh+9M/V/Vg
pUlClZUY2qMt4tTRIVwPr6vpSj+0COonVU1eWnxS5I3SG7qrnortZMEvwV94WBeCJbXQIvTjrBPG
qbqMQgSJvE25TQQnxK9Bos0xZBLwFlU7FopNzInVToH6GWMZMPQ9EPX4GR/pDXY3eHmGOTEfGTCO
t/1cJ/qNwmxH5CBCIgvLVfv545k7+S3bFPXnZNXnPJyLn0JUuZCnQR1JQDcfLukk93S+c2VHD5xs
JpyMS6tlZKYN0JzWSyeIoaqiblEC4fK8eHSO2HukDech9AVBGf1hkaU7zakYC1iEqWjVkAF0lMto
1A1cdgQu1zKEoDqFRDIQfX2DhosTc12RWo4Q1j3plP6wIdIuTc+NbGpeWqZ3Tnk9bs29MwCsMwiv
ekeHJ0lE0G7t61FIIt4MlTVkTqRg6/3d0NlF/ThT4kiruhCyBgDvMWwkl+QjxYWSVU6OBLOuaJ5g
sqmPED7f9u/MUvVS0/8VYAmH5Y0rN3EDnGoe7an42QNyIr/p29cDVu7MyNV5Mgzu69JLhrVaQtne
QUUOtJtGk5R16iXVGYIxj1bUrgi/AAbUV5+vwFPM7vkqsHw32Li3FMK8QqFYjUEDZCuzWWTiBZ64
AMKWV894cwj6ha5WkMjDj089VzaxCDBWlCHDR7B6ATJB5KmoxJ8DRNZ7cQMeEXbkbeqgKDKIurrx
Af0eyiLFAXaJmYuYI3/2Gan5GxEXe8CbKyHfO3m9u1rtQYP9sLMTzFnQ0NSsUhfcbv5OOemJ1VKt
BfIFa4YTcTGoiUhC7BgNqiJuiK4j7CTLn09JhvVhTI0k57VZefSowG1mauli+jCa7MdEX/XXSk0l
iOvLSo7rXsr8Y8oKLUGqj6IJVdCTNM0Npn4e1oH7spxsXjCRNHLnbjuRqjuuSIM6Fja3noN4eThL
OvhhrQXrm7DdtWZDzw9KL6a2c8A5+rk6aJZS7oCrwN2tqSbgcNblLGHRIpUcOrnviNIKMEXQYBvr
L0OrRDkmSkBRJir6t76hMQ7TATv3We0GBVNcGaYdsvC2Ja12JZHSLZXyV6vX9eGoWkXnniPuGdOH
vSmUWk8RLapDxJvE4tLti2Q/R7o+RLsT73gyenQd9bq8fX+DGI2JTdKyNZ8Zm2Kvss5ahOzu9SR0
OWe1ViKgzIcu2KAM0cDnS9VhhiC+FASTra81DvCPhRaTIVYUexHIfQgLa5R33gjSA6edbQKFX7sL
Ohq52icl/a4rMXgD00fnJGdK8AVXkwm3bF9WLHIBY7oqQfyDcCPOk8ute2lqYQLUNsMXZK7ME6iY
imzirW77V5RWTUFgdyIQi6S3CzcemC8v+Kw/3QNAMRWrTTxRUW3Vb1Q1la1x6G+tkA1HFyQaT9Ra
gwobvxj3LR5AmvldItjwgHKq9oSzuIjsKM67DjsINsVmK2POGZBWx185RMwg3nLl2GBjYX9akHej
05xUh6Mdl/caZJ97gxmNvuqfbG9sNFEFmkbWvfWvc/zoS+55y+HWgQLOvvAxQ2myBNhlKzZKhOX9
ZyhPDf8lKblKDHnNO9Bt3FlOJv8FyPXKhhQbCBadXqE0EpyZUenrZYepQIrBVVpG3/+5gmNkR5y5
s10JI1Yo/6KTlOD5xmn5t2dR6+L0ujWsMzMUjLiWPJA/ffGqic5xWafIbtOCPY8qXfJwHnW7DMbe
GXeqgl9hdiVYaibxysvKin/j5CA2FvcCm4sIhilSidf07mioywhQKCJUVrtQNXYCaCWtlB0kG/0P
f2EjPF1ahSNlRxxrEwTr1zVvs373LkzD61rcjvQINaSDfNUFCuZRMUjMVF1lZD7vRa6jWWbP41jx
5eaR6+u5YjKVEoOx8i8X4PHcNueD4gH5/PQUvYehiiQauWuWDDNGXwTtxu5cRTKVH8aiT2o2ThnM
pGlkxpfDbANZ4NWVMB3+rTL8k4/ZTEyRzqPeP0HSV+hBzSYqFT+6VweVWiQbls5l5cksqoQaHplm
ORFQ7zaFNIXqZlNX+mM95rdRkTZT2HRifLYwpOWz+z8mxCh7ZygGLb1IKUxw3vhwwhFqlOgPMaQn
T0MlzMuKLNI7ljgcruU5/CSZE6DKJqpIOzYiohEspzCPkiDnfVo7dfWJ65/0xYigKnY8Sj0EHjIq
Hly5pxwYsRnduw/idsUz4q4TN3DRJAhsRHNIy21UAYFF6/Sq0O890oLhxyw7wOne5LX2J6HuJCPM
tFgul9m0SvRBE3LXDNR3IyyAYvEHSXm16XGPWJATVE4VDI9Udc0ZxooeepWkBG1ghgdotaPpZH6t
/2s25d+ApOHBx1KT8KXCxkj2J7yrMw+cmO4T9yF1iPPgpjNfdxNT+tWO0gSgTAblsc52/dwaQyDf
o3lIOvaC/iWPRjAhqnkcx62J7EEklJTSLiVydH/8j82GmOzY0KiF1/s3UPlPJVUyzHw/iIvMjEUJ
ZREUfyrDeTMmFnBu33kb4E/TMSwO5cSB+HyBWAg5Upk13GPgKJTiUxzPJvTZE9LCpc2XMkKn0UZq
8A6w8CwFaeRN9KvJkm6WUIF6iTokMjZlPkFbQtYjC++xehgEMeFI/F1/EpwoSHMFhB1Klfunl1y5
1byRbHeD7thqjMQ4nUw/hf06O+I/nxsqFNT5UfR2Xy3vJiDdSuQR2PauKwIOBG3W5vqUB5npFCwK
v1yv8OTgoLA7B8WWHDFRUUhPSy1u9WP2pMgfGpoTZskFLPRcO8+YA61Y0N17OIsjYME+DQ0Qsnnj
9LnDqEWlAJS/YKfaZbsgutHoYFZI6L55WNXnDh+fn+hn2KL9Q8uEFXyiq/+qRaF0VugXN1qyJr/0
wuDGQuAeeZTK2pwQwS5ZgoIQeDF6E3BOa7xEdIKKqBf3uTWP7EPheyXWLFDLvOJST8Nb74ydAspH
DWoeVQ4mf2++mZQZVRREqpf8M7FYbPIeWthFvrOY5tDK510gtNlvgvbUKkLa0yopNyubrqYe4UXd
4ZjOBn267crZiG4UArD6c3cb2CSPHz7MboLFLS4Ui43aVUzAJb7ImDHT9MLFJtBM5byeCJ7IyYOJ
ySrzdAbR39LpVmpQ86as5mgEhO71vji41y9Ir3+vDD/QbojQTpBStwXHc7j90RfAY0BhoXWexdMo
6dVXxlq+89HEyvC/qUDfSKASo+zKmYPv+gxb89KiTLpVUWM7WLzC7Jv+uj+szJJ21FjZPzzMc75G
J05KtzBgvYArtF2t69Xu96+h8PIUDD0glUskiNw01Pq+iSiwqDXOxXiP/0uNyYZQcKHLaV2fWgl7
Au/XMRngIwp7fTnMpOILK9bWXy+8euOmjap84OTYp1w+amFGgSCKCT5khEd51huX6W6/oiQnz4uk
VIhxeAIE8nMBu9tsSdU/SX5aqpG5utGHtEsPokvHq7lj8SuxDNJvwq7wcDWuRtrRMlDJv0xWNtSE
p5Xao+0Usvoei3/77QYOFwCMTJURg7vw01VAFW0/sw0VFr7KorNZqIQjSCP4SUqELstUa0o6XO2x
wsRDHB8x9Os9+uRg6dYylm4fZgsk+Wy0l00lYo3wuCtOXURd7+HEN+yueKeFY0UydT08yf8NMZXH
CnL9vJ3sFETylwzsKYBaAo1ePOMo4sfkRGt6T0twVDLzkJCo2TaAA7yRZ3LQ6wDgROGBi6hpqjQU
R8iE5L8e7sZCS2RZ7va8X4LHVGv9mHSQ3J0mUI78VT9j8y7Vqx3evQUZq75ehDmdbdsYaI8vHBXE
E/f56+jadWG08KEDV3Q7kXI2Zilvx+hXbs7KQy8vkUHXoWaaTS/AEEuhukZd+/uvfKWuoFaSrPU3
dWuOPBjsB/R3aHBqbhf2JB7b0pxaW19uzd+KOQjxxeBIX7R+QMTgA74+PLUuhqbOr0Om5O/vL31B
WOsEuBi2olJAryA/BzeU3zjtmjFZNNrouItqhO98anXDPk5IFYeyp1lz+95EYy0/1tBM8qJc52gH
9hIE04n343gJY6SpfLAKyAjZImFYiBKVhJq+X8Nsuwwf68GU/uhHYCDMU0UF2ZyyA+06uQ2VSpkp
Qg8Zd+rHzpBxedXdRAhu/m9XDfk6t1VXT7DgBY8KVERXsWm5dhBQTiJktcRboIBmeqAbyOWG7Z//
k92g/pYduqAKByXBcJUMwNkoIqkbPOis9RWUK0j7gEGpZqeSknyOP1hL2tq5cXJPlr9NSoFnroYp
1rqg6p5/vKGehrBq3sR/zGJU7/oShRi+iaON912CFEFE3XMdsDBznc9SZP7BizVsf74uJlwvR/bn
BPgn8tuLrhfd8wNufj83ACn8dqxhGMZu0LDHNTVbesqIonitNXcCiFzpCuA7nnQpmojeYUeTLykv
6hZ9QDvD5n3ZHBlIwToDYAoZs5J+3dwjO5h9DgV1pbiFnQA7ymLkKgW7sGyQHnnt3PEWKyc5cPDL
Zy1YoAPa8U8HbdCaDq6P4G0kXtdMm3rAT46ujr4ku5dWvkCacc1q+kOVO0QYtpaww1lhnp4TiwFl
kd4CF10kVSgojcW+s4kZF1mCJMPEu4eYGOx4mDDNGB85dVW8plcYzGzJcjivrIvIp8mSpuEQ8xFa
pvLCEzRbRpNxLBuGAKKxLxOfpShdaK9Jau7MVlqSfaVArXXgJccNv3jXzmyl2jsvUBZXgNdzcJCY
JiiGYykQ7WMLE0viBpBJLA8S++p8o7W4hT4omwJdLjg2g0wUN6296/VB0WoWjwq5Vdn2PvdDf87+
+rpRWG5q60OfGGgy1DE0K1vClL9KBWjcICNGbtOU02CLX+W/sfm+zRNAYZMKec3bBKyHCRsTEoWY
A7+shsaLLDOqnYASVM/2DTF9Kn6h8wkPGN2fKuz7vClj0dC2+FnxCUl61+ch9H7hg1FgsdkNsy9r
K1acWmdkI0rAkDkRMTM+4GSV9oMt6oOpBw/KCsugdg/2EAxQS/dp2NHFj85sZm4SdDAlRCmFyRR/
lcLaSebeeevgnzle3Q81XAfKJA0tTGR1tEqSpFbj7jtjCD0tDvGI1gf6qtqfCELOXqZjgBRBNIpF
/8FP87n0VgI/y94Rsz08KW9v9BE9Vz3tHXLfz5FywI/tRb40ThFRna/Yc9e1JKvzcESfC3N3A1y9
HnnER5xybBsTH52p3T77bLUUsRUgd/B/r0aj1MrFYdi+0dqQm1cP6P3pVfPX+FgS32jo0iGBQUgF
98/QT5xO1F/utsh0TcGf8N9qV0JCIBMHFv4Q8ot5Bn3NBvDCguEUcRMySvQnykCyqN2pfaKdhLba
T7O1l4sRWRBeTyODnyD6gMVUVqroyK9tb/Ut00tHx4cYTjmTH2TSfdr3tqJkDquqrNQTl5PGi6fp
ZO52tFUc8HEwuZLSxFvQT8ARQfuEFSIIUHkwJnimjgC6mJSfgGQI5YxHCek8Kaqp/YFZSdsfnaMz
BhoqQDzEuttQIKZs81+FOA3xMl5tjyDq86rk86rmHhCFl7T+a8QUUr0fSPGUxKNh9NHJ5Y4FKhuA
b1yT9LpsYEPbMwGl/Y0oZg84M1KfvK/PrMR4EWB6zdC3IpoIVbi277w6iNwnL8+vyvrypIwmV85p
6m9k8sstchwghyYymL6wq/IydoK5c6oHUu0vNg4Jv/oW/VkGSGmwgiAAp5PTySzG2Kh7zOLG2gUr
Oiv6Y/s93zMAhnJwLGpbiEw56e6zlGTHdpNu3PMG9S42PKQYkXQ1nyGpA3JpqG5+RL09yJ+cMuAQ
+P99STZIRbSlbLAOqa9AAeca+TZl3rmNAfGR6h3t+JlI83Mc41BH+mIcQoQNM4XXxdKNAdkA7IkU
vThtOlims6Lo3T39Z6yZUbtJiAmwDs4xOHVX+HLr7iJCTwCV0N9mSb17+LJdgzESmrY8LnOqehJd
9hrMjqIbSz4Wz89bRrXK2TptgdBulT1mXhjj9rje+dYZIGXEbx3Ex1JwGY3sd8YrlMctMcxQDGRm
ZYgF+6o1qo2Fc/w7t4wksDfDWVwbPej6W5MCufnm9F5tzb4RydSY2BLyOIuB9hWwR2CkX603oLP7
5IcoQ8YXD8yAJO25E8M4AuP4nKmS/LWDzwD34aADsX1W+TBcAC3v1P4DfoT909SDpg437Hyow3wf
q6qRwpb44Wpn6ZiUj2AeYepEaJYAL94hv8+cXrTty0EQwQcuOHHLKR3kNW56Rkir9syC+ujDuHQh
n+z7AleUdyHLeNbnA/GADT5yA61C/hltrSkzeZqssMW5omQmheHUNSG9V+pzg3M0isGTFUnCdZGy
KWcmGxcB0h3O/psLhfe0WLHmY29N0hyuPZSJOSs8s5B4Crb+MmihlqqUbPjL29lQlSOOGyEozi2E
wE1vdoeTp97GtfBF2tBAGSWZzntM040Ycwu4WrL5C4Isx+N/I3sSqgUCB/2W6Yz8hvDQ8maW6KqD
wmxZso2LzlnhhpjVQ5j0eBxfJmp2IgcVFu4vjP8VdXtFCs6fxxEo1ffjUUp0YC5beGEHe1JBxP5V
kOzpHU3cQ72wL99HH+YlrZFp16UeLCSQwQsk8JtKux5jAQQjWXpNxoYbvhitIokWvgCoTXzbSKzD
UDMWP7dsllwsyVv/ROiFSBLYhyMczzT3S8vMxN1jxK5ND9NODlHAUDyDtRcM8sF8SAaDG7brEtTq
qIALibnrLJ2122p3r1HoI39yF9IOR/uQWJlUSB8vxIQeKOoHgcaszaPNzx0dqNlqfIgxKHovojnb
vcXitAHbBzn3mK2ExYynjjprqgK2n6KzsAWDUbfVs8qz7l6+rRGiXVWUQ3SSXOmLgxSKQqXNOF0I
JUnSs6tx0hQlWuZ6QpJ2ajqyiH1zWlIt/epaa9GGwt/NPybQwATNTqOf5UjoB3LIItKD6op7tzbF
N89varhAmVKPAcZXi5rakwM0QQNEBWQ5lzYI06+3TmSdu5rmKYhYFFOG5kA+fhsj3vHv1QlnBn5w
7cO4pNAkkDpGsOndEdY33IiXTCSEyBJgYqHqbrhIzyaQCMiVqtkg3ixPnqJTlIZYLPOyoMzcIki4
t2NngVPS6B1948kEpJ2NmO8O06sTADCb34pwsWVBZxwrJDFuzz6tZ5W21MLrIgc0mg+vGewEPcY4
lzTnIMEnSwgpfiiCgfU/5cmzglUePPqnuZcBggwOsvF74OLL+lGLpPxpxY32VZOMCL9iV8rg/P42
SMD750ZsHUb5lxO3XIAKvw7QkNYSMSypUigoSpJ7Hk/hfK+bJzVSfpMcOnpWPg3bcGfneqKRfYc2
HgfLlGU6pBQLzkqtbzodnFvdjHGgftbhf3EVBTyo2o/QfOYEVSYBkVlEeR6symqXZEOvYnlDrS48
5awWyDb0X3c9/Jq1wtnVsWB7FqBhawGA7+M8khtZViAhBHg0Ov2a9svOePp/A87KTgtQJkJ0biRH
T0axei8N7OdzIpmBowH5Kkjpi1h90AMMVmcbQqkeb8bw9dX9LBG2eSA8Q/G1UPzfLQbodFEqiyp3
HYuWoHfABPkYl/57uBu2gH321NUeSXxGUb/gf/uA0ueV0THEvMin6gbsmsPspkaPB/t0qg44+RRt
h7ri/YRH0QneCEDGNEjtuHKN4QBcpKenjiEZOh61laR8na1MgsXS24inaxjmxxJbZz5hA70hetqo
xcEugZTQTIqRjzVJ5cF3q3BZXN7/EaEoY/VuCrKlYQLjqd03/kyJUg/G4+tlNVlTqQqTcH1MMcmC
mVh3BEyOEaIoNTqbZAoDIVzeKtagcct4VcnrBpZVcGRFRrH4gGSz/qzTViiFPd3MpVJnnL+wzSrf
CY+PqoBC+0qi+gfiCckQpKBnS8uMh8RTrichdZM4bAeT4ER5VszICKdB8EEJk1GjedFFSY5YdHM3
egW5G8923zbJMfeuHt7yHWmCZKx/Pqaxsz/yY4R2IIiN+7oEXMySDqZiUf+j6elYyQT1oj9KuTS5
vf0Ss2BVF6HfoJGXbLVmmB+r4JNlU9yHLXgGRzAznunKxsnG1LcfSI+ZIhEf2ybbFinH0s7l5JTL
N7RTpsJIPTuSTfnaTt5pJcI3XlZr0yQtN2CLShN0QmoHt6HDxVHDDO3YFANuLaR9CxpSMuoa1DPv
HL7HxG/IEZFwJSzlQotZgND6XcUWAYwvVxNNyMc8TsqYiQLFXoKrFpaNUk5EJBjSl5JPF1Kfk052
rm8IwMMZoPwMLibGmaeRroIu1P0+LrLucJOiJpNCwefVfyEbEWs2YN54qEta6Y3xZwG+It7T5tw6
+YwaSuiTvPEBj8U19P6j+Gk0zG7x1yjL2x3o3lg7VJCOOUAMtvZ+9w7QmHyMa2JHQln49n9OLPSz
TPiCoRECqBZ1VFww+fqM9N8XYZHRpsE7Bu+RV4HTVWfAk03dVm5FqDKq5fuRrXSEs7RuA8/tBkqC
ZWZMbWqRFEkcvKFJwPcYyQgILWlBxJFbkIFbOuZ3AYlg5YCu+6jIGs0jlYl9N0DPE4WkeojadYvh
pemshyecuUMCQmeGB/0YiceM9Ieb6AsXk8Wxe9NP8mm3mv1laRs60EuX/MrZif4maMBoGmbDfuN8
z7phf1USV7vgDRIJdv5Z7+OAAG4bfrFkMHrsxDBQ0+MkFZfoOVMFvgtWcgFmuMXCV1FrYB5OlEuE
FfhKM6Yj9QA0OjKL4cLn8sqn8FiCFgS0Od0XpClJ0g4ln+jjK8EEDtfaHf+L/mb+jDy9HQfVmBtU
oLOCxLffEZrYLFgZPeXKxmWQq0p94jEWr45oVLQjmu3Xf3DmkTsGyMoxg9TvspvDniiGiNOM4Dt9
kdSBgA8XtpUxx8oxsZbc55zFeBL0msQN15YhzQIn0/tmCiStvO4bnQE4j7hJA2GD9v0u6o9nVZn5
dofGush/0NnlUywkLVV7yScJoCd+vBNdZG/wZuR9KOCKLWYlA+seRhJ9JKIimRnYRCrhsE7C++OZ
g5BLCyVPRv4qefhyG+GKeFGNxsTURGQB/qeEZO0aVXdRBh6xUiNq04/GgQUmswQaj2Y5HRzWVVfN
Wen6OM4c0vnQlyX+OsC7KGJKUp5hOZLcwF+PQHXjSjab5CP4JllF6pD6aGQES31F4A6jjvJFapVv
s6ywtif9xWJzj7/T9hDl52jMXOMRr0JH50EW3Ggy5cftfCWQuZspOyOr/0AbAPSQUTV2FtaH2lXj
u0rCxciYba0OgFzDUhZi1nQfNA+oY3BI67qgkyKahuxmgsJuLMTBWUAvqSlntf3nFGmfFwj9Yiiy
EemFQ6KBE+zQncEHOs1IeFj5MNo/H55xGvEZ8bCDdBEm6SG3vyQc3lUFGggAC9Jzb0PHZDy9HaV2
ugmNPRWK+fg54Yxopy2HqGZ2d3Ihgqr9xvbVgD+Yd4fNHKKRqweC3dqnE8952f+w0Ap0Cmjdh5je
s9Psvk5dxmM0EyFCOi03qmTTNpURnJVva0PTRT6kZb6D8cgucXos474OlCf/Z3R0raVZhVSYixAV
sCHFdB55cIXXik8NlGfBI/cgfPUx0arQ9R8Dxx8Unoz+mFr22tX0uJJ4kLDw/90ypdPgeUDUUKtl
a6Tsfw6zAzKs/eGsFg5DYrt17iL7i/jZgLBdYbgK/MOMkPfuEB/Kfc4lg8TmWYQe0RLoPwbK2OVR
ZtqV7auLi6mwAT094w+8QJp6cFo2lybWVVey9URehJUfCKcKBgpvgfAmpy+qi2vxpz2Cna4Tu+h5
KS+xaeqSfJpaJsWrRlJVAqLjbDv+sBDSbxF31ainC840YxDnh+or9CVSI/0Dg/fNsoh5Qw/W88MV
KebrLuvBRdBRqvi2fgyIR4zseIsv5TQUj8810tUi/B5S2tSbnk8eMceoDUtytZOAIr+xrlju/1Z3
nQCfcS/OkFb2UrgF79Bo7SiMedwhyK5kD+pAtNffMPySA+Et8kO5UEQ8DJ26XZpvMLzBM+uG0Fbg
rep9sossoP6GaaiuLGindEnJqyoel+PNH7LtH3AA1dz8Cskpi8lj1x2NSFlufl/k1AqnUZF3X9uW
odREiOOvcKUjmUQr9ecLhWpNne6W5o4ahq6ukZa5N4lp4nxZrBjlCqrhz+lo1WarX4sgmvrgh7JF
54ENYuadzKKgMcDqZCuUt7dvBh/jfHnBPJkX6ie5PvyQW5Oohyp4C+0SDJ6YxceW+apvHf6dXw4f
Ae9JfVfPyjhTUtLSAUdz2EvDKc4o/oSjLu5NyR4S4YrXL+PxVBnlAfn31OHmXxUTnYVUoMsVhP6n
34zPB5UuyG8/I7mUSPJ21gnkdi9udQ9UcLvsH2vDkLyX5tcwE494dblB80/f5Tla5TBOGGg6wBde
n9TFigJk6LoPjWbg9ybHj6zsNjE3DREJi1+xqXYbvgP+0Xuzh++p5e62ULECn2vCK54flMmOyKim
bkPTVLi4BOX3abQiZSRBPrjNNHPEvjt+wRRgExblnYyndDrDs/Zc2uTWR9VbYHTfJk3sqQNccLFZ
yCQ3qHUacDe/GQ1gnknw6V/odjHsF0oreD08Vty7yKC1tW0pXy5LO8cfj+4lx9hodCdF0nRK1Y4f
NKcqui0DU7R9yQ8qVn+IEbZiNV+8SE8dOqyVWIYorV+n7pBAx5vq/2tD6+FFFxrMd3CRUfJFv6eo
vZojgBrv6jCWmpjQ8c/P/QjSlld2pQVr1UJKWmKccoLl3lEdzC+4DR3RT3goNne78zUVGLoUQxIB
9CaM9bWz4ziAr3/WwsBjSe2nPr3x9cEQ3/WFfFa4XB5ZD1uDIr6A9G8xhSW0JvuoBaSh0nCukxdA
NK4uAjI37EA5451SspfU+Pr6Jvog3kcGJrZhVbntWGGCEHkrqQEnGdPGNQFV+X8r/GYEmBzTq/fg
xrjvSr6JdSXJlUmi/GYuWjfA24kvU4n1yGFUbvIgnBFnltewZGImrA2sRrDwnj01DC2+59UqilCi
aDnVDJIgKXbz/lAhbIcgOWRf15kYAeIEFLgqEKOcs4n/kaNyCY9gZv5Ofq0lF6aaWuW77c1JdMzE
o5UezBwKmXx/hg64oNBu+rAO0DVtO7rrn78ojjquY7nm30iCQFfdP8JutB4jNqRWBCP2fmY1nP+d
c9nw3roIwK4cEpfEF/a3yRmk0Ggw1hxlCfGp4GTPNkrE6tLq0gEpjMQQkHs9D5YFtKqcEpD9b15G
FCIoW3akTsyDkSVnqyNybLJ8Z4yUnNMHRIQ8su9cti4cHDw9TWhg5yDYZHhxVBscqAp1xnLtsQRc
lZWBasOcSCKgpLfWnUf3AJYnPSPS29pHJ9BtVmRIUWAIc+PLmzRi548P/PhhKrODcNQbA1pDOf/h
W6VcRor9ZE2hSSgilO3rhYm5aDvMxKWLhq3yeSd4/kzAAEM7ogXM0s1gYKesZg0dxUrTgWvTDepA
ycuNA7uT5YaglTDKr25luuSemPF5HQzkKex7ZAw4MBgEeSz1ewgQ6zxh0varwVv/D570WgdYxURH
ke20D2cHcmwyYmqkBUlU3Z2iKn00PXHI8EVSezUBHSC+j3IdIwMUPo29P87Fnyi3mlb4yPkDX+JC
BIEymsh1KXDaYms1gLioLdoxd3mV26hvdI44nTeCX+MoBtCisYKAecJv1x3cNqaYTE/Y3lcGSu93
RJIJgNUEq0cLnN2XBuNtOOU0jcAB43MoQfSaZmKODGdZx8ADOEllxAc90RnRT9aeD4E0yvUMb14x
BF/hA+llzGB08FgLO14uXgBVW98suP+Xxo7yRvhbb9LorvIEUxTUME2PGmCDpW5J6DjbFkJqX/6K
8ijdUEYquQgWVVOkorQlDa5l3FE/jQ/qmWFqyVnBUPsJTPvpe022eK3/Avc58nvlvgvwJNythypC
ooZVrLgc8vqlLr62tRVLfCjAO1wQA4orWacRdPMXf66sIfOA2jhFOCDWZFrgmhKwLorwbDaioaKx
cf9jP1NXpu+RCh7QK4jzJcCoKCxmZuX4qUFyUxLtLbvmEXF3d2Z7rO4fkry2vtnA9GflSep6NGeO
osGGC/GndUxGm58C2OQjA3glWs99KRYve3aPQBDXOmgq9TQSGvo+2AAmVyQngL8wAHTlfzJ4GDkB
cgeMS+KDu0pzEik9YeHQ4k0JlaxFXKQgd8qxKpEIFrTRx8P9HwEV245ByEUL51Tdrj5NuBw7BspE
0phwzTh011kBB9Fn5W5HHeDPou73nmrz1Hq94VZvCm2DD6exA8mz35cwjbxdUB2g2SyWg8ghS5/F
VwkZLG59cnu1n4kTFI30KuX4bcCf6VLdO6C6BEsJz0GdiA3G29PGHibLlO5MtmIT7PnrfoAr5ZnQ
pILjfnlLynaVnaJwxAfSQ/d/6SZWPgG89nt3RccdQfFkSUjHgyRClZ5gzgI3+4r381zsxJWogymL
GaJIa3XfBjSuU2gigsMnWGoIOU0uhcyQT9mvCISEkHAgCu35WktCL5P82erLXeJktkyHu/Sjftop
L+p4bvi0839/GFyWxLnkGolyHiA3o/4ouMroggigQRltcd/1QwXyyyyM+BOtzc+ExrrMw4BpQuiU
qSL6uc3bSYULWypnmYtI0msibbIrhMbYhLM5xpfQvYL6qy4WgxdtARMakX7CDyB4zyjKChc+ltx4
ZTotYCX/0xAPFF/iHR1Gyvish+T1umdLi2YRjxChubSrOe0pW2YOTbDfvvmjGM8U6AnUG09HOFw0
GOJdEQcn3+3piK8kOMFZSAcCOqUlUN4puGXrdRs/QzhWZUV9wGGTTdbHxgIg1CbmL3GBQBfgE/sW
vYsYSezbvpo00ZuNJnuPaV4zEeA5XiotwURDEgTFfSFESj1gm42HUur291NQH/WCAetg1FLPLR4Y
GRJloXGOi6hUhXUFKLP+rHBh/cXcOLhZ0QOIJwI/kc95EYZWg7cPoz7H1aH70MjKP1Vz0oDfK7yR
gnfxBmfn5pahm3sVGYaKalwlNSctao/tgsz0IWgzWXCZ3cNldPvTbO77Cw2W9QdOJ41RR3k5i5gF
5UXniyZH3laNQjuE1ueh6+vrQ3WIXVuTLdKM/tw45LYSRg8YnRqk/LKLD0T7oAyKmYJazpwJFViE
97Rz9xwExC2xFhbVscDYIXA0aV95rOdbc9mUGXJRe2nK3z7KOG9AnmK2vZwg85d4Qz0UyyrO7lIc
hRsCKPt1Xtzh6OtfHbPcdMI4MnvskeFUPHzebUkcTMbjiz0be4UF2G1FwL7YLyW4Z7l0ZczLcldz
7eCu6GYMF0MfkM0JKXfSadc4cuE7Pu2vHOTFxUUsSYgSldK0ZhqD+90DYividsIFI1QJCr5TSx2r
D+F9N5ojweklBRRHA4x1lASScRKjUPdQlhrKFOVO6kBWNtOwwhVeiWX7jwK620QlEXN4FWr0Nsqk
ddKFvh1MmWZikU74hIE1g7iCDwTqYbhrZWtnfpyB3aaGn/dkS0+vXpskoLxO/wOC2evMxtFlVg6g
UkvIi7i5fPnihMa2/eLljxJL692IDDL8uoeo6n1frUkjQKn2+NBxwdvv8znad48ElUiJC/btzPJq
QHuj0MHbIAD94aG/qw4nmrBpvp17aAQMWroEM8mqJLpnCifNlD561SHby16ksv1xmTiavNSBXLSw
qnMesBE3K6+ODfYMog75Fl0hUyTgKAkwUEJJUZo1GpEX/AmKdLYzsdmY9fSgP4qKWxYoJqhSCfP/
1bAeXavdYQ15HuX+DhQ7kJT0Fiw/Hon/LK/cVbg/YPXnbAziMUS0r422/idFl/lpnssRDMIxlucf
ADXoeuAoRk4Rq0Xgn1YbY7BRDES/RNIKpw2/lYjxSmlBeSR0YUqNh6aCkK4ivS5FJq9g2N7MuW49
IE8D/sXFe0JZbGn5xLFnleSPGBqknjKoBIrX9HiU4+VA2fQLE9n+0fDlPcg1X9zApz5WyNxuYLuF
mZq34BO0WU88nbP9+WpMsmnDWB0npki2oR0NX5yAZ5LQHpmlbZzcdUHtUSF6wD7AvXn0pJmVqmHi
4qBc+KRhix8/Sn7B/mnaOVjTjth6bkuITc66JpWmCPlF28CqKgq6ZB36luIfk0ixrACm4/pRAwFT
xYiWXIG2nsS9nvatD/5PGmkOpEl0WhABoNBWWu3IKzu6mAKBmuSYAQg+7rgkH1crPLsQnftaFQQF
kCez7qwPIes+uJIyr0gpEYk8sCKyA+Wh685suuFZ/zqGt0oZDPO60NLlRwKXjVGrv3eJaVlDCHUa
0mA5lw8ExAfZD1EKnkyt/lbiO+S3Ss0abTraJHZVgFVEg30FfMR2AW+gOjbVu14JNPIirGSV5T+T
+GXhlAc33Ka35l1inhfApnWxMDaiNHP3mIIAsp5WCG32dp0PXRuGK6iMzaaqKXLnt9AOfP5CHUU+
/6UgpFCapaWaZYDn3uuDWOpWxujAtFHRHczmubePkbsIKGjFRHqVOEvIiuzAPtLGwFxTFMHIugvm
5oInxypl7gL2DpvpImgvMtZ4hZh07mE5tBA157ZEpWMVdBnU9lxlJ9mYkfT9Kz8K103Jrim84qjB
7KPqhbHhzB0XCBAE2uj7AZ6TjL3vigKoD4HFpp/tEwo3sGjSI9RcQ5c5ZrSBhN4zugmH7ZwlHPzA
Y/ps1Nb2S54L4mvRYSlitIuSnxYUX0pNB2lC9IHXXThGzeyDl9dFRtoNfyt3UqRUn2Ceti5OR2vu
z6OVYiaWTkwwhoXqNWHqMsewnTMetsxkxC1ES/BxBNh0FPaZyqb4+/SnsLqNvC0VeKma2WofLqD7
QlmQadjNPp30TNMJM9PseEVoCbXTwWeyeS53suw58F/pB0j0RuRkqCFttDklXde3aouNw5kTG9LP
g5zXIjPonYYbuhboSzfUFvkKqYeoLGO9I5MZorlSCRHGfOy9mOjp8MgVH6pQK6NLqDdd1oQ6RVkp
+hjrU7tAI8117rJNub4KbwLAfM9ayVfn52HCiwHiE1VUja/VHpP5KEo8vOUgOGkuPSN1dbCxLCSF
qPeHoYRyxx+UTY2YLu3D/dOLwg12MBDd2y7BD4mBv5zlDL7L3ukg2bpO8u1UYAvnbMKsLtaxRCtH
ie2a+3JGHQHsBIY22468738y2VCeFj9jC0bdcyPzyOhOeqWOMsaQL8AO+r+2k8T/FILwrH+v/gTz
xm9Xh8/x6bL5uQYEVw+mY96UR/ziQgreY9BdkEu62KjCl4ze+Rp+DzkQ2z9ZctIlaeK+uOLXJTVW
8ctkbRIobbDpKNOSJeTLaaCUL+OMAvvGsUrKtQ5dW69P4Gi1S/iGtSiWxq8HiWHyyHbE/xsp0bT3
SdPNM/dumWOm/rLXQ1XrCwdSGGIMIfbJI7X/uhedIEUhii5vQHY/idPrw5e6zog7hCpeZX9afY3E
aWXMHudg/07PQ2xdiGNzyjzaY5G+iDPZ7Ha01DnzzLVvccnvKqtVBLDmWHk9Vm7vOVH/zI5P+F7H
ET8iJl4Uc8G8FjZPRLbuZrBWCAFl+kGY1Ov2u+PSp4op8VGse6CGF/dQVQzz7co8VxaMNzmQpYMD
N5rjUjsunPqDR3jylE3TcHHAXsWA/3NqsUh3AX8NJDc3zhrjGngTyTa2BuNjDH1bPvS5lS6gOZv1
MVhs9HV/RQ3f1Z0uR5ba1FhKqrzXnWq05yiASjPWKaAr29MH4ZTJOcvC5svTDh4x9P4R16cgdHZb
gMp5Ed2fMS5qwVF4iogj+VoHZ1Z486YK/rjpaaF92ppiZxxD+bAgQHUb97Epoyp6K3fxjPMgyX5Z
hKhXYP3x8LYmPUY2UAh+Dik4ZpvJjXnque3h/zR3SM5MsmOoNvW33jz+noRJaKBfdq5OYyIeHhHX
57t5GM57fSAe1t/0q3UWNw2N3yENtK3BsWYV4tRadltsD4VcXIlL3VmaSYu7MdH9JQFRcMoZRfGO
3X+aTky21YSwf9+5lJgLtbkY1w9mZ7tnkL2Ja/l484xl6wvv1Z9Ivltcc54gCjy6hUDzuZ+nclVB
wKZOTOIT5YxtH7FqjFFpYwL+FZ0BFyeJaQ428drpp0XqlJ5lbo3gkW3vzLg5T9CyzI6zZq7UHS43
6pZsjpUDGACYlOtPRWDsAPmITA9dQUs8/jLAm4Xpnu51VvHdxiVjlanCv72Kli3PkXMyTXyopTIx
SnSO9fFAFUzfyTrQa7xHUAXi3NZL1HqBGBtVcbW+liS/1dmXP0DWGt8x0oNI7rgHvpFJ9si+B9Jx
cn9oAdYfBaWz+/1tmPYMTX0FgTAvfppl/A4/o3I1aIttfQgSOTHS1aDH7Ho/jkQm1HGXkqgFcsG2
GqCRTW66HPqfAjHfrehe/2IqOlet1Sp2zpKmNUWybU378X8LUS2HsHkwSpICdTc8gIyqwqamsZqF
hpEfCGb5RI7u/BRqfZtUOLg9pfFS6F9UD1/3ToGRAO1tY/b1sbc6JDHrnKwPcjiUWCKcp2FdQCSa
2ClM2umDFK27IFQqw81AZfLzqR3k4MSX3/afvdVvEu+mkM26hARqRClOANqVqwe6N6Jf3i/idVRU
YxmUin/2zF0qLZXWKIpJ9fFZFHsCuPaEYf1Y+0o/ylL8Ep+xLNF9JQPjHGbJX4LnIxNmKyQBcO46
h/EqF2RMNzbZLzeHS4ctEHTuIRbuKvIPhLz13fxKIdHQETBYyL39EYqAh5ABBmIXCfqZFC9YBU+z
d4uHqFCLzWHbREmAmSpfhMGNxqlj1OqQDrl6qv+FzFIaR94T3RKauvhUmRgHLweUgubPx75G8m6f
cU3gEO9gnTxRzOK9y06UxoHpLzIvn5eVTiSrF6jZA7PG+Slw8GyFlQEd7YKsM7kHo8xOnHVsKxiB
N1oM2UjZuS3+RQoeAKggfpN+aUE7K6Zly1lHkXzvpYDO5QDa5aWGIi2WKD4Mturc73+TZTF5fbTB
ewNHWD4m0tW33OllUbXj0LhI7sUFJoUWe1vnDxHqNfGBNiIHEISL962Gn9/M13Rc7uxCKk11n+jq
FplahDPgc7Bz4Csh2Tj4GmZshFaWBFsa1Z2PooTwE8vWEfIXgg1JurN9Eo6HjAG6EPCM7eVGU4EA
XoqjumYr9mOekvhO6BQnFJnJmPeLy8nKHElq883jrJXC5k14nhDiCc9uhQObHXkLZZGvCtrnQXs8
+84uAzrJM2FbgB+9/W+EIHZ0DpkEkldEN39kD0iE1QFkww5WQxEv+UTBngNKeKZvtvJNJdyajaGz
i/G0yrStpvUsiU9/NIpndXlZuv1qCy20JziIqCu39b8dlSO12F80qYmqTt3jxEehl0VqrMo/qFAX
hUFGKWWLjAgFvFWN4zqNlXBfQSHhXI6G7Uzt9MnjCOv0ZeFuDSh4KcQSftpxjZqAEJO4hZUfs2qQ
nhppwZM41bXwza1dUEEQaESllc6NNIjriP83KCvseHyqvgwkqjxfZ1N8qloMOb6LzLMxx4D/Up4L
JIgqhvxUqEa/GGdymyFXdW3U4vDjHtF1SfD7t/NTp64S3jonUGwGCtqClx3m16JgJ6uK3QxZPU5l
CYR8ZY8SB81KJfNHXlXP7+pGnhibFpZzJ9m2rXROaHMn9uO8kNWKjdrDttjxY4fnu+9+ZhAAPYb4
ouTjuWjDp9kqBkxWq8eOfThjgGS1ZjLuIirYZujhj/Qeh2BsSu/Zjw0s8g0WshZ5TJcJty7tMhBf
3Tz90qORIKIY9CLur7vS4LfriScbwHgkuh7FOp4oinRSHO+tPbVLtq8zW8LDvlVaS+86wtZJPjtD
RG4rMcfxTeqRGBmfeQc6QkPU2oG/+DXbbm2vp9Xs+I8cjQLNSjQ8k7txibGAleM9u21OKa/CeKfl
Rb9M/ubTmKFtVYcuXVuONadHAjtqf+9twF0OpQY4BJ+Xe+stf5pXNYP2lBQ/zTcJ8gvhrxmn3dtP
joHKdgUtwFDG5bgU7aW76mQ+VEV2vNEXYZ74NYvMfOb5ay+LPBZPXEV+uy7xbOOes6ztMXkReDop
hOq3dbiw6DK0oT/H/7uQU4Ndr4gjcMSo7ezaMMfUkytPjCGZAhFjBLpUS8EpeQ40+uAYLJVIElRE
A0Iy2rZHEAcNc4kQm8qs4b7UmMGLwijt+CX131bnJCdtVX7LFn4emCV+O/8NaWltBlbnog9nSdOx
Apk532+D5p42q22mVlvPMzugq51CwDeeuUAn4RiHdXF/CPeaSlrCfD6IbYwXmIgQ1GNAqdbdwDGZ
iBONUKgCr1ZP0febtjoKa8lYLU8Pgexn0/IV0dCxoBlkHs4cBF7xhc6ezdwXSVsJNMq8qEufHk2N
Lmxy90gcPHwbJBHGkLmjZM8opDH3I6o3i0s0P+R7nLcWSNSN+SUsIQQSyFq0AcSlY4dswpQ3L9iZ
a/OYT1yr+QWpIYDI3lyv87aY5MJcZNFtPA9uv1tDJoD0paxppbHmHg66Vhvwgeml1v3NukHIfrRC
T4tl5I0KPo1Wc+Bd2MWaZKVGELZn16CthKWxoTmDlexkeVP37h0wi/oCSeHpaK+0o//eGNzK4Y5F
6dEDALcMmkpaC+Il+WMV+zsHaqiGAxJveJ7qnNP/VeQJ1qUCYw/KAWgzEth+sUk9n8caJlIyIuyv
n3F6HyxTy0atFfpK4Nhd9RI+6a5HoeNyQLZHW1SZOSolfGVkACKXDbcHIsK/s5XWYwqm0JnahGJU
p3e7qlmFngVcwLFSZyVhMWlZjvkOB3nNS7/KCgsOl+/6cizbx+NYCULPhdrr/cNnhBXijUz9lzBf
OCxWjD9Ct50w/nnnUsdylMK4O9xID58wHcLiui3o8cFFNQu6n0FUEMoiFL4hA8WRVQ2k1JHG0tyM
3fbkpCkTAU+LYdU0G9/8YJnMB7sHEs9zGHT0dxBDbtD92oLFxa/Wiq1UXY989bZb+Rhv4XY9BxUx
dD7Q7vdfLp0oZ/vMWoH6cEShQmTKcxePmQzOAMDLYgztRQcyxIOrPpl2bnPNOgGkdJNNfjmdwkjO
RZ4GQj1YhrG5YFkcDCozmKBhrTHdWzryqktX+lMv7v+fORgrYpp4jLqo/+Lt6NWnFmOuTJ8GddIa
x+84fhvXmWBsB5bKzOdyhJMmKN3MWbBNy7CTpyuFX1a9VmKl9LdgaqCWBl7RSmbC1JqOOUczOylH
+04CQCclH04sTnvp1fAJj8j462UIlFUrN/UJ8BhUGWVcmpkBfh8aeWADbevDTPjtHqMLmDcNm+R4
AvS8u2A/PX7hzwemXjkCFujee77jzZ9U8RISraqayYwol4NzwXYvFDvB0Mw/Wu1hl3BwREAtOvAg
XMxhdmm6IIsQRzk5ic2NPmSX+yN2526LZS+Abq2DSOzVDWZydPCwD6nWBPYAUFBtAU1rFvr/GyVJ
FSRYP1z+Otc3IY/mNne7jcF9dk5RnVfhgE+WLjJZbLX+J3nAMzg6EaQ/0vEmiG3BUb/0Le8Dso8o
qKyH976U629t+zyxWcPYXQMulYF85rzVwhEslpKzPFv9WL0HmXzwNh2UiC+YhlPd6x2Uyxm9aoZb
N+pmylyAAJm/JtJC0mvISB8Z1nPFpP7sv+u1kcYojLFx2WKIe5d7RhUc9XBjLLulcJ6ML1mRTfMA
l4iGaElWoOlZ+xmlKfp2CMBG2NpBPNl0e/Xt399sqpYn42c3Ljbxw0zawSwsj4RLlgWqeYYfSMS1
nh+OudFyFd0Cyn+C+mLJCXLqOGqVEN5CcbEhagQUQF9KlfQ8d1bZOP0TtRXdAwrJn8ZuqCFZrVia
zax45M3UhXrxUI23bn1I7xGWMPU6fDFZ+LzlO5g3K/1ux9TlSQ3+mxCxA+1PTv+KYBLydnFguloE
z3n29mCU8+Eh6lKSSwdMqxgCVovWR49As65YmTKnLX0zAgJOK7sVpq9h6NXQUdRk+kumAcvVgz+Z
og2JWNIjn2Vb/Ae5FUotADBpXt0Ksg+8B18tLtYcsi5GitLSJRB2I+eG2v4W8aFr7syAjMmcFJ7y
lQyDHe/Vp/aSTL8hDKT6Y04xv90GYNuL/G1wgQRQoRGsUgSIABHyG15ytZkcJfxo5m4WiXRkiiUC
TIDIBNpzT5ojZmqEyuVtG7mqz6b9TNU96Bj+MbhOZZNW1dEFKUDRhoLXqf4Xoooq+Q1cUjbGb09N
Iv+QbeeBBPRUkm1J3x9KFZK9t5danDkEWZhC1TmI1YEII4hO6WYX4UYaId49FuNdssDHkGgkgkY1
eAgc5VyIAof750sdHlRKWcfPXD8VAVi29DNHyMqE4+jF7xLIarirAPTb33iubC60SDGEPAWrwgU+
DC/dGKL2sp01iyvUiPmyE6P9qbK+oVULWmdQjyGElbOjSbKC4EbNYQu/hI/AmxxlzOdYW0cOvDVl
sB/cLmANYzE8K9YJfBo4VftKFelzi+YkmxQDi9yxsN7od9jVosos+M3T9xRFcmIMWHlAAnKpVLK6
ej1oL1cnXTuC1LBtbBUpEPjK6qnNjoHWfyiWw/paHkNIdnvTUj0//eCKIgoBIAIqBKZllw2r00Cb
TOmmO+ychF0Qf40xgtSIaaxydHgzEPhjtRNUM2p3BfD02eSCCM5NGgPj8tUP5KG0h55OvUiybFr/
CGk3IBCfoG/GxrCGRsc/6W6nKniblvhhH+wZmwnXxDpccINZIqRaPu47hy5ljw2qdJ64ioWwtIvw
py1M2cdBzp3HfNtp39IYODsPtdjHJlTwvZN1lohDRHXJKTfDMvRbg4Kg+/HTm9asXzvotcI2XV8r
Zd4cDVAIUrde+fn19u4dWJ7F+/i24x5epoihwt6cuVHCauJoZaMaiJz1SB4/algx4PW+PfHUY0W3
KIMQ6F1YHQJ3aMQrCgOsqezbvp44KPesTFaayWn/deVpteg1IYpERTkAhusGPaiNktcxlJ0Zn6g4
4BXRwzIqfkaFjD6ZC1RZMtCBN4lBpmkSXllrgPe1O+Hy0tcOc+LIQgenWSDEpyAkMAr3AHeBJ7cM
LtCOCYMqeXnu6BK22HvhNqMR+SKYs+q6WLko7EvmObSlIdxX4gmR21QXEAOMCdGr0k3Kz/geBFd6
nP1hmchEVjB/c29O+aMkWQDFYisoLPYcS3uiSWydVdXd/6tqH50H2wi7Nd8hwuW5OwbfDd2sQ5eD
bOr3M6UCdNgBTa96ocqwngHeMkYeu6ebz0PaNUD04nriY5ICRk60CXGhUY4BD9XHlt6P/XsaHVjD
6tRZz0BiEZh93BnipyNsHi0Zo4eIURxM39bEPMrs4DvWxBquZsMXDvOcL1we20t+hxPW8vOxsq3Y
TQtKpsXJmKGGATam9koNtETWh4dIT/v8DwSyvRYAFrB56grH/+JOMHsI+pZrAMNSUzCb7FS0r/02
qHBBWfcE9n1gN4G0UPEcyFVNydS41hqvnfGyq0XybiJgMKzzyB6VvObP18BjyCfmR3GaUvjIi9i5
Szbovuy6YsKFI84bHaUdkKdh+eAwjG1MLthguQoc5dbxCRXZe7nM1VMRHSJSS51IKVuoxI7CQXjP
TZSTA52bhmaTKia9J/yHjd6vLiji3jmFKuRDDqKHepkD0jSJuHA9ubg7Pts/G36tQmT6hrDGOc4s
dVPq2GKv2D+NpDFk13aPsWdZlCG3Bg/H2tsikvVJ69r8vRXI04h3od5HIWMZOL6aehgJz/4pUnJx
VUGV6NdKcgub+f+KjjujFISol0Scq9yDsxv/HpzUS/GWEQtmUZ4PAHCVgyHg53JJlXyi14ds+kXh
Bq0nufOpABcfeSrRos5/kOk4QJQV4ISunnVZmL1jPE5RGrsUA7DlnkbO+4q5rPl+cE4b9AneAtJ8
738ChjFTw303ENm3DpAo3ksp8FKMa+DQrgqsMwkAD4aQcOrRz0P01IaiWXO19D+U5Bo/NJOevz2b
7mDM/Pckypk7PT4ZkIVjT1yPJVDdNam87RvedWVB3BMnaEJHRzMKw6Hvf2C4X+opgoWP3EJWhGI2
A0cvHX1IeRbcrkm5KFSz4hoHPvUtPlM6U8odqB0wJsL0bkJKLF6zX+zQWnFYfNmJ9tKKEAGSiN93
tD+Jx8Le3nEwpqAT1PAg4VgFdVyXU7+lRevwmhqlblEu9FftYUcoiE07rZvqLFrVzcoZwQ5oLC9d
3a8CDte4RbSkSEAa4wHn05w/LM6yKAYDg/viIoIBUaDoWt6Yef5LW8QrijgEteHu6DFVGyA+SKEf
OIub0eKPcnH4Mx6lRWRXYoXWBihLwxRkfF+TvHLcWGvZeJNl+9j2E6guRm5hrF0Kn1Xt4+N+TNXW
6l7o5ZGdLKfycFL9/h/QBKW3eAFtOl9LxONtP8NA2QJquxUlFKAomrHoTjxQKILiMyXJjcuJm3+a
wV255uF9/5c11zbaq8I/aUDag8q1jx4RDx0SV4IML9otduX8wnIV97MB9KmktGOkfjSIrTBk2rzD
Z3ox3KH8FYRIeqjh+VJufut++ElZwjJaosKvonRoOGYVs5PdBzydysB/cdnagChxyo1DXS1gafxz
lbDpE678OpSclQ8uKCxh9us4dti8eBO94Tc4CiJr82cfNULHqo6Dc7jX5hY4Fd89gU59dku4G4LK
FBCAZLRlrQcO11iZ2a7llzxT8NNwb3cukKTysp6adBcRXzTLw+gktdGGqinZtuoLb8AWhGkFeyFt
nx9jgSBgTg3FXhNGbpCLL818H4i58HZ6CpN0odl2bE8gXrSLkglUSXmgtAVM7Q9X0GdtnDUMrQX8
nnC10iyOezJFF57c/UarZPFgikQe0t1vyFLq9JOK+2f6rD0JfCvEoJWsxkRxLIVDZBixHU6L2MAT
Q2jookO6CuQEPCyqmukhqtztsDQpnDinHlo2gfFS+Zm9DBAitk3Krw57YZyHr+TQY4J+DyXfNZ+h
mh76LslHeOFKhStywfVoP/eQiPNZaGEY1WNCUD+yuuA+ttjZSvbBefiI1lP5Yrz2mlMH0hLFPtps
/6Sato8bJscZ1r4r5ua1pC3CajIFjcAn9bMELitzgH5yraqUMH6u8IFM0qozQ5CQVi7edEckrgiA
BmlmsOQMOBcQ2l35qgkcVV60xn+9T0+ntHGTVcIXo65tumY4T85+yPBKcfeBgc7HOXcDlDN1BaZE
ORniR/kfgM9SsKcez50/8GVqby+X7ooKMZeaYht26/RT/32x29yZ+zw4DxHlVhwHz99Aet956qCq
TVpRQxPDOEKJ2MFwpYqGOQnp3yaVAQuxpxHl2lNxgqUv0qfSwayP8OPZmvTKnmqogf8rOjjpeQDx
cBbCxAzyy3sSyph5JqND3yam/V+n9hQSZ1mdvkq6Q+Q5QbWmTOoESHTD0/vkJwmGaQZRm7h4h59v
/bWNtgiB5kEt50jW3KoC6CGLhJVaTNWqotD19OYMryb/sEeV8Y8s/aNzJ4gpU+hG02qqkNIHGyYx
qvO/KPpS3nYzdYu6yY+gScyLqiCpHGXM8bWhtv2aH7qGcqrDF/jlsGo8i8v0A2F2M1jXCLnREbjN
Fff7TD3/nxU/C7h6rZvJv7iP+AEHzjQvd6xXWCpiltIWId0Soii67GAG/noeglWQPR5Ji8bLbCGB
SjXE+bORez7eUMjvrn2R2pgB0HrMaPsmKWzNo/vDr/roJZ7IJxFPdninSeJwN3EWqqORmnc4N0Hn
ibGhYIJTH9fFCyCvJjQVBVOzM0X8GgF1EJHaZ+G6XT58x7oY6XBuPO/ESDjCOoVZ4PN2+woqJg0S
4bg14IjLSYpibz2H6o0vEGMY5xXAX3UXZLH5cGqXJy8z2b4LhfLZo0a7CrtlZUL5KzF8rP4tMQ0E
sZJgQ69gms69/4K7w+PA3LG0icVmYyF4zSTHJa90WVt+Bx/t12AF++NruTLFq67vn0oV6iS2xBx9
SkjGB5xPiv3uqST07FmwxIT3sQcvYXxvXS+W6ZWFdfg2Z0B2xbL8bmfsE7ldPwSn8Hl04NBvMyCL
KJ5+7c0t4g7utim3qyKLtTQ2abLLt7aY5IiIw+7Usf4Ve7VYG5HUbkWUUkNwTOMcSUYGDrxYwJcI
00hsKKJKgIP8gTtdWUUfM9pc8z3syBK0KP+u+UVdqrY3FwO76HDVVG3hhzr/M37F2TMDlf3QE9/Q
0dmOKDwys/hD42JDEIfsWdn4vSh4sHjRshc5i8UIZv7R/L9CSTcBOO6YV0jbvYBy7nh9UH62crSn
EM0ceqeb3jUMeV8PyTkXB32NXCCwNltELhNQlE2Y2ffhPnFy18KplciRftUxaSK/FxrpDqwndWfY
MvGVBwI16ceuP3ol4bU3d3gWtBfTBMrg2pEtkiKAOAfmTFF48fU5BbU0sVGcFupXtMh14wMEXkYr
LfjndFEx7d0JGbFFKqian2LNOr38SN7ru4fNbFcAMkeYCguzU8xd0siC6a2Knpu39gk/GZrf1j9K
jTN+bXrxoUYki4Lk8ec3DO6bEgw+0y39K4CfXVghPTvZA41IG10qvt9BQAN9T89qJo08VZDmI/tL
JLcv0ZEgavzG2UcdUBR0pOpz69Xe2KJb/K1B0aVwqdLdGIuF3oXEJqLaVji0Xfn/Rqj+PcnFX8C4
9UMR1UntDdZnDVt5yMi+CADc4oJoK8LsWE+p/27X/ANzW1/MHQzrqNlytaOm1SxEetiHeJmkWZjV
7ImaUsdU1ZEyTY1d9Vdbkz/87u8kSV/9amfed1ZLqIpB1DkM3h3DtQz5GFFVaHUtzFPL2/oOsY2A
1dANq0aKq2L5HJMl5FltUfg7xLoKtwRYHmLsuXr8HoMG5kwkCdylPuVcMzF04p827wotsHgQY0gA
q/g/D/d0pWycTz/lZ91/pbZ0HN3X6G7yG687lsweyHRaP/HFp2FhlCbaq94HEMi8bxHd+y8k8hKX
mxhoX8kkLD5LX2oN0RTlzZTJUMn28G4UgT+laIii5IXm00kG0Fa9/o18R40xgNGZccEyXAZSI6lA
lxhriRm8PuZe0diMDabbEH3kxO+kkQSdiKYLtW1x9R5YnOO2toZum9Hc5R8FIGp7lINs65EGh8Ri
Sm58KoCWZ5PU4gkC0Yo50DkfgDjgVR15b7atWRKT3j45sR4dWtJYZU08XzYB9VQgJeEmDR28lg7o
Fx+nheCmQp4/PP57xyj7rSMPmg5z2rxaINWkoFUrIlg/BhsGLhS1QYJXMz3eFGdV/B54CbBJsvQo
DRvd2WA0v4aKEs1jFvPX2vriN/qfL5xhdKBabE/TmWT7Zy3yufQPrh7IxQG56ZdlJhZOUT4cKf2s
AYaoK+gw3K2A+QSf/v69pq+Erec8sNP3+b70YhJywNeR5lecna1omtWrNsA72YtiFAEBuvclEx4I
t/eqm6ZYi4W3hMMqlGrhCrnFhVDUbInbyCCJnDLVJRGKDgIAJoAN4XL2yl+vBZqgTyoW56qYw9s7
chPgQQ2LVYQgqaqoTqgG8mugfQ1hzD5O54A8zZC65QBG76+Qoi1X9Zpexv3J9yY4Az8EEsC7QkA4
ypVcL5c314JqRaORQfj/9tp3IV2gq8VsY7oAwDHe4pRo7tkcXu5f8pxFrcxmBQfDgEW9GP5Axc9p
uwKjvzd2l16BGSJIdQcSjW7RtytvNXdTvJPhUplgHG4vey7DXRW0H2mNO0pPRelrnfsYE+8eBIBg
LgstzY0/YnYE29O0MPw0yb2lCZDtpHYBCiesSiHs7O42E31BXcmKm8Z4mV9NVsP6xXmCEVnXjsZ+
ustU5acO8ZvEF7m5R2RzoZJkzw/AfNwHt+3e3qxlLRbImfSW239OgPAem7IYduBjT2uc9aPrajLd
BPPch4dXZzNcvDOSfg+66krDMRrv3YZqHYjjmaJwAxDGejry77I2s/dqx6qFfoH2sWbzcuxAHtOl
TKWxUUdm2Ltk8Uuf7E3fmhODFahx5QHlzQlRS5m15XShVk805XtWrG8wUycQy9iZAML7Y9WqZI8F
WwvF9gEmgiMAc6AD42/13E90rpd+4/99u1VFb8t9lPBGKw1kyQ54NtyFl7fuQsFRWOf0q2F38WGe
DKs+z1SnGqE1vg7cLQPUiF3Ul2qdoUGV2tFIQOPToT0epYgzamWGz4nUomL462XpY+nD6iomAlei
XKfJ6HZadu4IH1+97NUA+4DJ2yj6CnY/TIKrsC9VOsocjgxCFIL2tSLGhvoigSnGigUS1f34R11d
jzXupVEpbheaEB/HJOvyTGk872h1RwuSUX+WxirhNRY2CeZWlZ9DQMBcwSnxt8Ri8Sy66Hb8QDAF
cWQAmY8LGqW0ukzjhki3cN8KI2lL2TA9M488CUwKBvL1MTpFclfT2B5ZATzpxwmkEPo/7ltSbaMB
TkJLRnzTwNCwXXWhMQRXlZQsjlXyemLK2jXCIORKyFXWyEHtVqJDQE7m3WZ4m3+31eSKpmUWUz4W
mUrnAVdbkzC9Wqve3xygo6yqoUCWp1QJz9s2NKbMUcW/ZUVYu+yOE308IfwqGnzw5+NzHFtMZsYY
9cnb6FoqDsvLzoePSLktoaukZc2QJk9+1Egh6glbHoyY+ENwSY2SpWH9zpw6O9fBRYBmuznRD7WV
K9JE1xoP1hSUjGvX9gx3n1m1lWv2y9Lpoqtt/NTBhuIIJQtxIFXpOpbevyI+Ct8Vn1b9ZR+z7ROe
Ok+4t8icCterhSO6ZjijpchsJZ2LpBvsjeyv1MgGIRE5vAg0TFb8K0/3QyQGp4/CQJO3LTXCtEQl
SGPRox+jA4KT0NsKkUrmeNbaMk9BTrtSCDLUhX91hWsa0V1UbwFVNJ1Dk92w5O6gjIMmAg5Vgc6Y
xVKvvWvpmaYkot+ndu3JHmKeJPK7DpIQOpW6pejIo1MRdJc4HLl95TPYnD9cqxEZR8H+UPA6YoLX
UoadXrP6rtDFk5hyH3PqsWSU5uV0uT7X+Mx9XIkNBwF7JCoPHTP8ki2A8vAVJlnGq3KpYtudwiH4
i1Ix/16WVKs12jUjxGOKeFSCluxirEtG2ZiG1dxtzJMPYkTYFwOu/ujmblXTyD6hxHTkESq4FkHf
3FQYZQ23ffzqAL/G0SzLNJNO5s8+ma2FPAR/2sv/fiYkOBGSlR0n4EDwI3OeTZV5Tr4s4EspjsIl
mEaVnetdJy0Mu7XXOZgJbpHO2LMF3I4M1OmY+91jvUlCvQCn4TOIImaYnanusfKX/9ysrWKxFaXU
ErOCGzm+YZ4q/hgB2+vU+LU8WHrbliO6wbhYAsL5v4hRcfxfTFTcPAI6xRgLURDai17JwKhT7Gmb
Ehm/7wFspN+Pg2aEKkxOvSTe92pzfEdgnPF1erk4AbZXl+vt1fWTFkjuVw55KKRk5+ws6P+C9nTy
smrU//FdhxF0sAo1pFHZjhUMLytIxqHM4FuKQpV2QXXPsSoWWNrWdnD9JxYQ8fpvMzU2SCKTSGcL
30pmf/lBrLsfo4kZIWKOlciSS5l+DnxAhgzJZ5YnNTaXK7vrh+xfsVOA3TyteJJL/9RP9xwpyswM
uPaATJ84AptGmQCShQaQF6/xKFy3E71VN0S9+ntqErmgso2ergqNJe9FBvJVOnzICeSpLaZ/od1J
6ptrHWiri8GaLM48CM8r6KZl0buTpIxk8NdxGqX6FtsAYkKsxefFJDDK/vkb7o1T4JmvirfilK1M
YopaRLyF5HmYhat+K25BYpyXTFdHZ5r3vEI3LjftzVbrr/423wpvcDA+aCr4a1u7ZzRSy1vjlX+S
6W0YttFUDygg6o5PWYjvSd0UWSZy9+Wr9fVqx0Iq36vr1EWDjn0NRWg2ZGSDywgbgWGiRvIP2b65
69WSxxw4KhD7y1vWu8AB+sT0LEVmoObCtrzkJCU22qROJZmqx4GxcLPq8kkjwF2vKdQf3eGzeSss
w9+mcXj0123jTZoF9WJvuCeQJ9egdWWU41IENcw+CYXRQ9pZrFEnhFfk6PmO3BAVL4pRoYgSAnWb
6k1+PMpgY/N+GNRPg+Iur4zrZqZVMDqd0B259aQvQ3fz5mjqFenkyjhd8SVlUQEXRRratQeloOb6
C+zWnxG/1WKRwXCn1764YXro1Fxi129gvfudGnGkERnAp/EeL4p8Tj6YwXSfKZC1FCHPrKJi7fUl
3mDtme+IFHwh/+7i9QyyjmFW+NWvp4q1jY2NXPps36MBGQvpjSF2X7pjM9qCPrWNFVR/T2VblhRo
wNIlij3dsvYMzt5uUUQEOIdnGHRLbxUhDr+bUO6PjD79+/4JSQzS6OF5ntO84t/NM4khOWP690OC
JfFb+mNJYL301ZOE6iUso4LYcMgkma8vqJLbGRrHhOQv4Ocvb+sbe4NIvDmPMVfdxk/6Yz3Pl7Wl
XUF9t8hKtqtRoqW1Dj2MVN8+jF7a+QLvEORLnyxfReet/iavh152eXX6lcZRNSznSq0jrcKnPjlL
pUmlqZW70gVM8xjCYvScGdPucTRdyo8NsbPhbXTkplnPdzAt29tQ6KM4W7QVC+bTtq9y5meT6fAn
ej6RTaVLiuUkWxfbXcByuqWV/DQb1hWum7mkw1vt2uX6trq8p0OTvqRi3x9oJJJuaVNaiyqHnAGI
2Kdb1HE7T5l8ZtHFBHXfFHNT/9K8G0pSOgsENYLWsX+BB9xl/bG09N8Yv+bQ5svF/q40js4M7Tu4
hAVM9lq1i3Mb9RXDHEBad0HnQ1LXLddwvoarBMkV+uXPW30hibhYPJQ9U8QQgkkQQ8oulpTkTtK9
7gDZM/COfW27nAN+kD1FQtGKBo2XJkje054//BBpjM82/dd0Ei6cWgc2a5UX1HnBGJT1DnHMpXKF
WbKBCqJIUSr0O6Akx3ia77w4c6r7grZCVg6ke4Q90qW2TYBUf3w17YOmK7AVon4J5HdnGdotacmP
kP8q8yGf4GTi5kpZTkMvI2Jou0XAl2fytjlC31dBqiPqTM3oOGvDy2/e8iG+4j3cCV49+py4f/N5
dffipuN/18DYKHXxm61gFQ+AjU76kupitOqC+vPjJTt8+zF96r3DpHghQD7hCNuZGt0Lrkt+Co2Q
HcLqSmcEBtwV1Qu2ZU/hx6///kiMxww0jWbJIyEpqCl/d8AtY7+7AaWW/RU1LhJnF2AkpE0xXn6M
ae4JppkL3Z15yfXEAgQYxvJYbX8o793LByBYWdCorPRR7Q+8dadyH/9eZxwBdHg+WCHWpresOxLf
bf/eJKKL03qooBLiFnysgafOQNZ/rubD4QIks6HYx42SvOllP0r51M/7+fBqF2kcSwo4Kq+hoqtF
Awn0ZhksGT7aWW0P16+w8MFKKMkYKtYp9kjyNIUU0TXIZuihriq2XuH/QrvU/qGeHmmmuK2t9q27
7KBgmLrD5yV6UEoWmWp/RrhSF7YQQtaF11vfLWWBJi99JFa5YLE6r/prZs4ebI3pnEk9OLW4esX1
ayskvhRsDSS6EyJir8/PUuBEoFqBUxALrFsYATFQ2o92Qpb29Vf9WWcTi5Ij4akzgo0c3N3kU45L
pNiglHCHpqgn4sjMSv/07ZK8ABTyr0MZoFl5nDQcuB3CuiBwGdswr8Z2vysLFr5rcZ357QTGKRXi
k+8XXRXHbqMZZwwwjqvhKqmZv42TclbIxH58lK/PS1/Q2FQ1HP8iumSMvn4gmk1nt95xU1Wns5/E
wLR+2Lyk/PPhHOJccYLMqyGFnC14Epp88FkSfnIjDpM2ZdHc2vxWDbOrYVEAyeTN7eOV9RhKFbOw
JUVLzsGcGqErbWlL9bmEaf5orxryvgOHiU5DEhQdvDY9dy7Nc0GN4+yZNR3PmRYlz/8Jd+7GydjP
52cSF6YU3JZDT3fVUoOtLfS91cQZNva+ynSBR5PeCOc4taVyMIWrTTzdMOtpVrQlykKAaFn4ptDZ
cIeIA8us+lM+7xz655217a7ta1vvtBk+vCvHZvVGRyDSro7tSyA/6Dxujo8TP9yAbZXBAfjHJ3J1
F4LjUXyfOUZrA0qs1fJV4c9PuMzitistYv1zdppzUOdp30gt2SNPgDJlEKByt0IIz7PkpILkOMrF
Zb82ixVM/HKHg+nowcZovwJ5+fY0U+Tk3KMIYvaMpM+di/fRGfdkgK4pemHWA/OAgXb64OrH4xJd
UCtjQniOZRRo1M4EImp+ovRaK5pc+J9PV7RL0IeRuDlJ9WSRG3r7ULeW3vZ/JCP+jLQiL1QoVF8s
sRBXs2u+RsaavrYEsxHFjedYYmXeyO5QoAbd3wOjLjfH44GBVYDXxvXJgwmijSKteWsw+OdDifL7
Nab+uXS7bboeslu37Bk/M/DasOiyZ7DuOv5N2SLvon2BeV/jc7MAoZeorH4r4mSJps7W95QUEVxN
8ghb9Ae2FfY9ryeYVjx1l/kYIjlFHVlBa7dZbRsb5dSp+zcjxpPZIHhL3rYfaJSGDavNVSPw6Ejq
c4Q09RkOoJEyQLd5mytJIalyRNLZCJzM7Fywz0UEjTP4mQf4SLJ0NQmIzZVz7HhuIun5Si9pKYp1
hCrqdLb1Lv7tlUopMAV+kqNhqz+MsmTxnzEd/gX31KgL3tvPQky9pNHSU5bRHJaVbAnNvt2PBfvf
oSSPSeXwhVA+gkeKtN1Q1kr8i4Yg7zTTWsGj7XuhZQeID3aa208jOJiCHMN7i+68ZJER59SlEGaS
eUA7LOsFgSeZKr0QiPmzngC3U3oQjqXEdJfxa+i9FTgLjxqnJ4akXRpylhx1dfqglv85Not5vbbr
Hsofq92rgFCQPHqzUaj87TT3QR6ZkYrSZ9yG7dn9pARp4kXMWbzhnrGsMhVpIOz03iykb2TNARe3
6cIYm8WkobNb47Wy+usjNsLXMIE/80149Gk54DJGwe8YR6ZW89HMiP3Sbv01scPxSipbOm9fjOzm
0XEvjWqOJnLaLiKDkGj99WdpbV9qZ3XSjP5AfXFzmdq69PEAVDZBhCh/7tZ+g5tVr/sHD6ETlXf3
er5y4TcO7b8ekO+J4Wnhin750Yr94/lNmKdg40s4g2ACvqUJi2tHw2vnws4r8qhw+mwR6C7u3Apk
L6YJMiI0iHW66StgnVCrR2m/AjWaHff6lm3V2bBk/7eOPHvZVpjHGUaVw2gulC5+SwaIdrgrbPys
N9Lbxd03+GJSVU2dqmeG6BD6lR+zMVyMSrIfQyfoDDy/twO9+uwSrF8ogbfbKB4aFeJowEXSUDpn
OpjOi0oMNl9ARB86RDfqreOFN8XOuSa7qdtLSMaihLFbQ8X2xifR1fOi8wEXEtOe35w3nM/YHAHA
733byaEH/mPhugWjmZ6C2Y04wCMlogCl/lxfqZwjawyjt0KXWXOiHywWNZ1WzLmvfV+OH2mRMiRD
bV1nk65tYr7L2VbOZNVE1+qiKpFW4pPV8iI3BExixAKpzVCKCthZjt352iOwLMBiq4/mH1MB991W
ZCHEeZ8k3ZAKcnc/WqHmf9CGXhn+QuVsEgMJO2f0LES+6ngWun7b6mSoBTGOLJluV3eeP9BUSWkF
TPo3oDLvNb9oYdsrqk8VHaBQW7O3QcTluLjaZRR6JQHs18gjrkyqZdA7TiARNEdSw+9W6M+87uP/
f+BxJ5eyZ568hhxBTfKMbpXnQxvJkwr0XcJ1R9JOQCFbU0K/hN8irUrzAFsDcvQXhV55Warn3NpC
vc/pC+WTQjHXXj1nOsHB+0VTGkc7QYEO2366+1ibXVjOepIzqh4sXsfTuvrMvlJVoFVDgXZKnKUz
5qToWCeBk/sqgnfEoxOZKfhUR2rXSJhueKH3NfFfwr2Kc7tSC8GHEb++2XTGsgDSGOMA07BWwxZO
oQxcPSnSxGm/bUxrfSO75ViEmleobs6otITprumMqpF6YNy1at47XgrOxIMBEvMN+0tZfGCynMok
5OXbvow6AUaryNNw9ceUSUWxzL2ydKks4TTMytPrDEv56CB36ThiXtvE3gIO92vP3YLIJ8wBKTgQ
6M/KecVarPT1a/8hpEu8Fq/WXQykr80am12WOzfZVs+yoSNVprS2/X5UH4yR8It2M6tdmf+hPQwW
m1N/lztyYLA0QgPlM8FbYvpKC1NJeLIwxGKhAsyd72H69BJz85cmk9NxYW1M+e+Ho33I6m/t7xqN
MOoofBdZr73+9R2QqUpaGynS6HqLkgbUBQ0HuJM3lfI0z4OYZZjshC2JJDa7/jML6zPPYT8ZEPsS
NODayLUdz5kvXvZa46J4GVaxEzSVfHL6SIMu1ucLh4nb452sbsGVRBRDg2qgDDcqGN+b03/0I2t3
FEbADHP587xqilHVSr7jiJN/6HY5giM4+03tOsXz0skoKCd9TBR7qPYPPUOUAytjZZgKWE37xlUu
edEbUOxFsrkGVrotgxnDU1p4icl9TgNH6oPIcd+EvrQ4nGFmIsa9eFMgU2/HAKjtG8EHmnqrbU4I
9Me9Zrv2eoJquCSLshVFn2EoYsGgx6jV5oLzt2yBXOabNWNU2i+zIpYiXMjd988OofKxJ0Sc/ZeV
sThO22fO2GAd+Mxk5jI7yV8bdpldqe+vDfrKkfNE2yXjP/60syuqEZdCg6uCjpAACNBtTNRKFElL
w8aTI2/XIFiIRqqfXr8B5r26m/bKorE37oMM8grS+gYYmGEOslj6oQzzMPkb4+XR2jsdbfjSOzge
UdSTXAraWzpEiQdyhpH/W/6IeuW3A/bgGVeqbStimCpRhCkhJacYtD9ajbnqKAL2bichbamEjSxg
nxAw4NMOgQ+cxLzIOBbKWgD20S3lhsgOQphNvZnQHyrURspjPCvcbZcu4961dZevxgchshbhnx/z
HRrXisdHQuBP6du9FGi2nxKMbZ5MG2Q/LwsS708QRmgJaT2VQDsge3zzmNXUtbbEcA2C0xXoi89S
livwBneO1BurbgvdqKzurHz2Mx37hoNpE6F/VIEAcNeH4CU+33q/Pu7ov9826OvAWjvELhKafmsp
68a/UK0a4mL9ZWqvn913UFbF+W9IhyNozbD0r3vuAFK3956aIPyXAK2OtX3kPMIfB3EPE9kN/93d
FtlFEBzCVaZ4exXKZRzgJDbmJwuwNHg0D7qxhi0P7sPSIoH7YutHnsfXr05s9NdWqaBTNVPGcSmT
4E0p/1GuqtyPw8VXZV4CIGOpL0AJwUhzDSXkFbzJd03DdRR8Hy34CLkw6TVIPo49r7r3k2A4jYw4
JITJlLHLzZkkPYWpA5WCgDtAAVKvtNvfzbRw2Hrq3iu7iL73JxfxdpoOMoJjIaJxw30KAYP4/wvU
kuEPV3c7a4dKg457umQcHqwVt21yqib4KdEU0EmyZk+i7/yuW2wdnO/A9foNfqTv0lzDAx4gaJE/
E9VPijRXKPOcMmt3U9OWt/OCuaXANBpDQWdo+3KfeGNFcFs9Ge/azyov/Cx20vOsjoB4HSP2leHq
XUV+xHzyiB7KGN829w3SVgv6TQqy68ssiwbjrykR37ynKZuGK3RpwOVw3Ez4TdvGqWQc9hEhEQp1
pMem5EynkwFnPygnTXshemftm/aCllgLkzzusDDJWevk+/2AGUo3l6JiOqI6SNXvSycxMR/rWBht
BTQ+xvBHsuDrxdkD4AonsjbCb7H9pcRuAFwHuhdLmU7uimzgm97Wt12WrUjI0Uum8obgHuxVXtIA
6z4hnPuZgAT9LJmOgUcfRT1uais/5EFRuFQIaYmvs7K6+J9JVk8JfDyttlWzcsKdkhfERjwC9A3q
OoOXqas6auVb/gKK2GmcqebgWyNcntkU97virrCFEMdNgxChx6b2rzEUzASWlXyZu/1yYXYhAcRM
PtmflAtnlqaSS0EfOiV9xwZygBXHCY+TwXdC+FEJ0UzS9p+IIavKRbt9F+0DsQV33V70tKj90j4C
NMdUhehFGxuayX39mdFgnHkQxbpjhZVHWKBWKwlNRuYvTEDq5b5LtYwDmd3kpbObJKoZxGNxQ/xM
uyhoJgSmkBy6a4DDTRS6MWwbTs8wxJ/+EeKO+oilDWMt4dWhU9p6nGzbVtAUjJIMWwlbl1ualRuP
pbMnstCLDS4D7+yfk6p1upnLqWxh36X+J6ImpwcQDk1MYGSyLdB2DkFAIWzRRHdbyVbgvrHZog51
TTENTONgqbWmpCQ8RBmM/y/glKJeTofzsVUW8DnSu0C4I/w7ghA6Wi01EKaNV6+hrZvhFEgKZRBU
4PL7XfAJ+mf2ty2XitLV8Fl/yuWpobBJUbMgR6+ytqYWe3JH8JXjda6Mq7JTB8f1UZk/RsTUi4kh
Kwbd+5ZDcNYTDaLC+xDA+QLQNKqPZyK9CIToFDm5po9iW783oblbeqKTpoqgLRfvMKw4SCBRsG2C
cy6KkJjeH5CDkuZeaHCl8L/F/mtZl9afEOS/LFmlnvpEOnRvbRBWX6DJTk6lf8sgswxG1+qlnyEF
KG1ynEn/E6p6B3TU8d3kAzqUeuLGjvFd2kWSfIg5mfMVkoMShPBJJRBYZdWubpRSpU56qUCN8v0s
kE5Iv1wpMQHz/iNQkWUE2Vpg2ufNZvf3sOuU8fcAhIzFsRvzXHLHdCBtXkYjFsrrbr2jiJpRW6PD
gAWB9rJ6MgGh7NWrMwyLdNiaAqtA/m+DVR53ouvS9jzr+AwKc3t6YJdh3ZEgd5uycIwZjlZB6sLm
MXYbFe9oq3qf5Dy/k3+TFNLv7PCbxH0UUcdFUBujVhyF/1EIm+yKmGfNoyfH9zvLJzFur8YiPHgn
D3cI/VlfZqoCPwjfm3xQ8P6jMHkXYLj38T/DOTjU0Wgp0zrChedD6yybLHnijyw3H0aAMlS8w4mK
ZwVQ+Ixqa+m9l4XlsbGarJLuja3rAUhAgc4qbBbpV0WLxLwDxjrd+RTpTLzAjUsojrtKMJNH2WQn
qn52pOJEm/kj6NyORT4ct5gI/1sY1a9gG9Co9UQLZKA3fVQvGv7JXxUAjla347X7WbGlwLsGSWj6
JkVuDqNFDFniCt1TxEZnbnhoSbVjszy2edazA6xOEiKxn0ybcsTu0Q9it2tbA2lSZSpW5Nv+xQQs
zlO5MQcNEVfcKwQmoYmkZDBSupVyDc+UuLZw3WX0t6RnXONS3GDr1iIL4G5uBCjnHJNHESuSkMVG
iEE8M8yGEFvN2qfcitNaXF/1JsuPN1k8LBoyr8D/wuz8uk6ZwLzW4jf/gsLF33f9ddJSnozHiDNc
F91ROwtaeW/pY4cwebVePmbW1s28+KFUP4Pbzbl9AHzUKpoWNVRZYh1axbxzr3HZ14LxnvSddbPq
ni9sUAAecOFcv+7fWkFVwszBKATsfiaZF2mXTOIeAg2bSYJ07okUeXwqjLFDv7kdThzXDLmVF0Hu
v8MrqBCTjWxzwFRx9+q6gpHLacpz7OzoFYogmDPK/t9dJE6bb/QX7gn6yItlftW+La+UsLVekuLw
htcVkYvKBj+UCjwkWOw6As3EmKIDHQUuKFVM6CNR5I4PV1X6NKppaDAtKMcP7dvNAD4zXWlkxUFN
mkiNnbK9dzOqPUA+49aT8dgexngxuiUhCNULftpGXDTYTyJgCCZRrB7VH7LZUGTVkzLsxXO9E4Dn
NnrEa1b791ClOpz771qa24/FyhRusQmka9tCYVAXZLJw0zN4mShG5hB9hITdpGqNtBllWoKDVVwn
7wTzYJpLTe07Dy3UWw/wX+zIxMK94ghOgS/iFlcnq32d++5EQOb4QPLuNV0un43EbT/2u/ezXtyn
TsmxMHGZy4kDgi+mXpKPbCW8Y6MlNU4JGCwSPj4eIjg34Y4sY0Q6lWf31PZt/Nmc1EltUJs7Ftzx
E+E+kjJta2Ir7H5rxVaIsiea6o36WgNVVbMbpmXGj+nLMY4glSpYUgj6M98VmGL8yc4l4NTx7Ixu
Nf0dcUrltk7iAKOESj9S9ui+QedlggXqOG1StzqTOSCrb9Hi8urkXkZDNqBWSoUIhyQ9e4J9akAd
7C46Rvx6hPgsA/0Cd9ZWrBHc0+a9BA6zg2H35B03kgxYftV/s0DEi3GXAxv399elljd6SvnrybPM
BImH48d3yppUanmFoUOP/fgfOCjUp5pQrAccVZAdKJBo+Ua6hZodKRyDSGsySWrmUST0ub6XfnuH
5gFMjFf66btid/7h592DH0FsfM8+5m7p5R57n+nT/eNrEXAwLFgdCYHb7NHue5YUpw6ea4YR4vX8
StBJzBjbhcGprnZr4Tmu8C8qOXGz34vtWlOLgdqJPAu/2qzHtyxNGT0f22Qy6G+KPgIgPA5p2YTS
cKjrcohyuAGejQvQrAHyS/pDoMyK6FdVwcDcA4Qduva/F/PKgbY+zdEiLwyWqAABFjXsJbbYsF7b
Y3STFzRsKELTLHXLShpN9LAdK6GOZfklleUWxKubq7EnrYo6aRakM7SjDM8N1BWqH9sGTqQeda5s
47UuwoMgEJS5kfDa+Zai6CQzLPNPp+z9NGB3hQhyMXyNUZyR04mzHdnk/kNeixkeWPP9qaTlAara
QSXTgmQg+srUI6aRRXYygXHDBLkBF6D2czNqeq80gvhrPUq5O6lIvfH0dQmoYk1OwzwFl3EgwUxY
tGHdkgCg76Yea56IzfOoqjo1S73Ajp6gR4B2kjqKAA43mQVMK34h/MOiTf35+v+KIR617Fb2sVOA
1ZOUvzknBTvn5qhto7QZgfens/evKfIa87n8H5Jb+0fq13ymtfees+QO7Sk4pK6ggO9Bv9xjuy5S
BjhoL+gdR/HPzAPYiF4Iuo7jD/a62mnzsvXlWp8Jpbh+8wmkWx4gNt9tEu7Lib+eWbeLBdEuWi91
vge6vKPmfK1IOMvK1yEC+Cee6Nsz8LRNnsETMHNko57NQwnHyJW9GjLxTS4xAnlVFMRjGAjWwePI
z7IXwAo9pjKql7mKOYgWXkDiklodSOic0xi+rs3M6517t45vSGqp659KJuzYKLuLcuSiIaSwtMnc
vj5ulEF0F6TLgI18bZH/704I3k1abpyTHaATdOlt5RwWAW/PJ5YdoZ8APh7TKbLJJQJEvQNE0imu
hE9mYEM4QJJmkHCdoYiOdcuYOewLJ4bPIg3rX/thSwnU+WPfgVAFImPUT7DRbqXN1pMFHKbm1t+Q
InzYc/dzYKluoacCXIk+mZSEirg3EPJ/9sIPTtnCY2Ek5IPl0FOApwJG5E8r/oxKYTF3q715XNMP
bXxmReTEYNEK4LTh2fGRrSel9IvT8/BMdm60fkT+M56N7UNisUMHLYe0OzxRfWubEFFis+4ICj9Q
C5hVfPaIbDpox35MYcRwOH9zshmKs2XaSc2PUT5WYyuwpG1wNc7dksNYJJ58craLM+ycIFDYA3+g
vuPC3ZiYYsVq9wBrOVRHOvAl+VyvGcqcLL0gKf+PKh+dHTAHkyHtI5kqTV7okzjyofj14D/k0fAy
cbxRXWjiwc0L8u36MQxGxd8SWhJ0hmfG3sv8Lms1tnFlP5Zj/YTkd/BhztawZMAC2kzQwkv5aNsU
IQ9xqJQdGb9mUj7cGb/Y2py+Svy+2r4uUkVjVcV3onVgFozxiwm78oq1NPivszqvxHD8abF//xCP
6T8/UWuG3IZa2cdkijL3lcyZltOWxffWDijFHklV2k2G1IKR8EquKdj1RNih2bYk3oGwzR3TOBxt
T6yuKJz1ccZoMI+QZpzQwkZJUMFuZ0MfF57UmA6Z48C5ZJBaOht9EwarxduVz6hwxRa5ufCI1hBB
PWt+8bO9WPDBb1llDYwN1bjXJpmwCUgvOchPJikt11JtnRjcIUkWvwPVBGxAnCPSUbpMN61TMAvk
+skXYdu6NzIcm/NF/R5GSAkAVNDrkNPx0zFW+2rqID3vE9OjP20ZMdJLYTxKnO+8dGfHG11P/eCP
DUbsa/o1qE96TqXwk/xf5ATZqGScD2jd0lL9kcqLw4P/JxRL/jBNQubQUXA450vURBnjcia87CMO
GHR9NF4l0i/94LqcKZ5ccqMf93urgcTBRv2QLuW+eOdCjNyzYZ7o/nOu/U7/6kJNRtNE0yAM3dp3
q8lB/ESmJy3pXqBuTTqKOYPmkkK7W8iyWAZdoDNHDn2fLUZyoqUkO/QvLQmC20wdfWslaAr80fon
nLn6jCc/jNWCt6XC7OwN6Kl1K6k1tKfabayzLWogmd0khdLwSiMaOw/QS1u9ACYRy2Y7VsRt1oR5
nqjgwlgO2xvCdJvBU6hcYcFNxCToYt5IIaFw/k4jumS1lEXZYiDyJemezzwfpg1WT+DyV74Jczbz
M4f2rgigRTiWMTYitZdG+ghjCS+ePmUZynWo/yjk7qjzmNFiA+HiJWUwIuNllzf2j67OdYGi/+lc
M8K4yax1O0GrQdWpETrG5ZSunUp+Z3EOaT2s1QVip7pBDdQuOsGOkxcd3A1wCI5UTBOWVwR5ZeW/
P6ubyXUqO707Hxz9AK2Le7ysuor0HxqEzIg7/m0ZeLYLtUxrDUWT1uZTVybrH8dmMHe2ML1SbeXD
75opvD6kOyIbZyG6nMgpW45/bSWCpE7HDytMbfNqeFqVQ77sGR9bPgeesx1vQW9y74N9XQF4Zpuy
EGKd6Es0o69cqc/NSUrgGD2031rou2jNXlgTdWicJMKjrANXoxSKruwLHr+qBWdfLVQpcJDWK/Tf
aXE8m3sApkG+jraIjY0xKoc3qyLc0zv5HrISmrOc5lFlmHr+PgLAlKv1NSlwt+jM48VUi0Ora2kV
w1gdFtBzumD3WMDUr4ZMQkTFJexSo97AqKAlaHIhzLhdGhk/jH6siHXMHKRVOd2xP9dv7ZjkA0KQ
z14WJbeUuZ+JK5X0uxUum2D43TQsHR4AyNcozU82J7RD0vgUT6+XyneZ/jVcWocRge/kpkrHf8yD
GwukK9XL+GDlw9f/FE9bWWNy6Z+0MoE0MwbiP0JVpPJlWLvlpx4AIp/wHckekHFLO8Y5oGRDroBx
QmKfe5j0JLDlCI30tg3qpMH+MnyeTQ6xI0pLLcUmDwbjpo/Fwivh+FNgShH5oWqCIyw5EXgIO/BU
NorzsBQ3SrGlda4K4EDtTJGqI0HvNr6U5bL079QnG5seCbr+fgrG1oUWmY6IhV154ALAO7uW5+6e
/YLwvlWmncK2CdulFwrSDVBmPfsr95227zyZUHGSSnPkl1wVDyu4K7lrnGwgZI9egaHKjZAsScnX
ed/t8oAr8QJlIup9MEfpWIRJUrEsRvofBpX6sE+1UcoeuVGWHD9MWcSw6r0DJ8HA+yz7e1ssnatq
46O+XioRX2YgfyDhfYb8K0d5Jv0Hhye/I3m8yUkWPHQrw5KZsnbPaakvF33Sn46yVL4GHyNeY47u
cz2MBWzK+tu0RpdfU85zAa6k6sbPwMbQ9X1E4/S68ppUb3fwEnrOqhsskvu2Uga+OoFXSVLxdT8h
86LdxwVPVx4vATlvsbbwgUev5QuoIVdZtY3kaMM+p4atWiNSZWlmI8uoaMcc3Fwee4CmuUKg+lEc
M0N1Lug42CJTSD2Jg2fidCFwk1sLeWSa8aYRvnr9F3Wjl0qLXvYLCwzo+7Upir9bFcuQ/oNX+sJj
eIkoeu5glCXgvZAuGSop/h55/rrCVPNgAZso60Ef6ezhW2bfyXO2lcQxY7Av8OHkefhQWp1iAg4O
nOE1T6Ly0Xprd54EDBP4LYqx8pfgnTu5FZH//MgSlooYDi+3i5BAnTeR6WU+kMk6VAwaZaaUqlPU
9mtSG7Ip34fex2R6fA+qd5fa3CAUjMG7+yedzMXIIkG2I5RbyAyIOeXEgWKNL6xRsGBppoz3UOG2
jcHpagRvdA98GHxJganxvUhZJpwZrjchAlXUmvCdav/rwEMRGiWRHlxjMakmL3NJDqR28WdPex+x
vVQ4BdhST5ckYbq5I6jcRr7ooYQfYE+GEiseRFnYecHndoRNMkC5+JmZGvmq6OD3R8RfsP4bBYOm
e5H2rcXh9pIgErmmaIh5e708ipoQJGRdIk+DUrE+FShGq+OQeDjssGI1F6ID87oVRRb1op4EAXWx
/B0NOp//u98XZ+Y5EpCw7UDiv46VV5+z/zV4tqh/gdBpTn3qjjluiYHVYlf9cu1JbRbNhKxyYWQw
JG+nPeh+r5HjGISvtrHl/kAGFrdVpUXYEAum6xo4RWh6z+wkxbTFxrkBE4roEERKb4yWh15jYegO
jD3eb/c9elorsspnHwtqDa9+Yhg/UBbEKXcLjpWXUbBR3b0Gb/Ojt1Sn2E1PBEGqN1T7uVq6DhQ7
fvKAWHL2rOLb2eFIb+Nb/yXjyXdWSN8eCYIWzoiQW31ZFohv0DkNJ1ktK2Nk5aJvIx0Es4fD6X9Y
+J9GzBWKrhq3O0UM0EIfDQyh5QURcUVvsWJfnuvLoVWZWDoyvRoc5dUjnnmAeE+Pmufvvpdbw438
Jm6G4zbsbmVz2Vzac21cKee2pkBfele3YKnu5GY8BO/BTlPi0KTNZNJVoPm6PS+fCAO1PG0VEZhK
EmtPRRyLeVjw3Qg+XY9S5fM3cYIz/iyvM7/0DSwZjdFPIT7xjjvO7NKvrgrr7Nh5GnT5VivwFO6d
YASV2izlWD0Fl2Pnr/L/JDjbZ5z8KY+xEZG85Ipj2IWJ9+46xGOfcKlrTSxrvfGCeE8B/i2jf47c
ugyJgqx37cWAzX9NQnS/oKr3LHUrLk5TY3FEGWx1CLxhKh22uZpNL0LmC1UFRoJG5bRCHz9xnF98
Sqz45E/KrVd5Apx3w1YK5Dir5RJffRRH7YrCjun0lud91SDpQ2keApIcqBgNqr81np0ixzZJz+Ie
825RITPQIudHTaJGCJjy4cTgvAZQSvxw55nT4iziZfcLpilMim98SIhKdTd73JLmiKq68MxLqVro
jwnd8QRTkeh4PiGJbBNC3Y3q+arjK8nhRIeDU3WVVLFAEUHYc8XXBzwGWyDRGSEMqElgPgNjVnYi
QXmeVLQgZ5XEzY7iKjnaW1SHznuS9lj7IGfvsV4WQQ+dKo4DOxnoNP7G/w9QXHcTl0jH7v1y/P5z
nqX7tCsTOT516DOxHGmlSrE7ayUMGiacKU4gTRjz7lAp2lyvva5kmjogNstsEz7JjP/luAq2Az5z
+k8rNYYj+HFFByg9X6H9KtQOZ9p6koSGtk+psKgt2pBH80D+jiGUM+lmonG82N16x7j8NaE2Toqf
jjAAEO7S1z2NjKCb37dSDCobTe76H4TZf0kD6bEVGKP2B22iGlE1venvprbcAIjp9MtJVv+O4L7u
gbKlsT2QYJprd5tny/+g4Wg6tPj3dLjc/VGQxYDzIIZZIV8hFFWHQXhd1WfzKMHUfOvnPMBFSlwc
SOZwYXImxVJSD1wHHwn/h/gwmp2tc2BDyoToqUNMZ+5MU+AjXd7cMRu9Rc+0R7KEUnfonzWkJBBE
OAvmPOWrNsLT9xKpKoGdq56YJtjkVMkRIDUDOznAMTFCI/FNU6F8FVWnkyjhtPr9OG3lv1FhHk6s
vKE9caJkcp90H1BimkJgTQm06/hmMMUAINxA87kq7PNNka+i3WL7bVQ+TQt8otjOuow2qBf7MaX8
3bMf6IV56oFcJmq0vZOEXjk1k4/DUiyO1oyfquim095RpJCrXRs2Vm10uyVD2CSJtz8lqTP0Ar6B
WggXTR1MdNPg+aQ38glCIOAtuG+iIksdq11JDH2nCHENosJnp8y/SjBwx1J7Il2uv6VY6QizIxom
DXi5BtvbNz2LbwFbwlPIIeudE+b3rC3z3irX+D96L2YfiFTjS+aFUaGQNcOh0KaVeYvabf58fyj7
3wX15pIGgV7F95TjQIN/174OY6HHyjl270hAIwkwdxgnFq1v1HZn4/DWcqf9uLAG/vNNgR9ga9BY
VKUFVWIj1TPodz0woQpWiQqYCc6uvqkfCaETjDhxk2kJNkaWPEuY1qMftlW8n39UmZrKKQyEaqkT
PB298ewqLjVwmzmmllbIC84PqFXhsylvTLsm76NJnxVmcs2bksD/BkOLFBahtuYfsz3OyIIHzrW8
ojcK+E5qCort4rNZqjCagfxbh/AC37SJYk5fMAhkRwu2rPddUqSBe/m9yAXm7Y9TOxJThVYi+NDc
Z93YNb5+x2LM6CoB2HAPwGRj2tjRM6V3UGUevHNXz6aaBKrBJOYyA3tsmuute4XdX/eJQdkLIRkX
cY2muxhXX9bxD87OeD1xpmgR8vFJeppI+wyhF9okbHClZpvWyRrVivgPTdzY1bK7x5dWAbDR71rI
pXjhURzzqtw6als99a+T2R7CLYCzvM5rchGoNtKL0wcOJExVT+WOhpcvGCUps1O78el5rLwTRGe8
mQgAUd9+JpBm/DOPq1mTm2IcNiVVLFKBnfYP1WhyfYkiWvTKUCdGQfFhiQpwEdTqo5BwC5Gj4NGc
2ZoLanQzWCHESONBAziwzM8V8P8BhPkisOMtVTHji7uV7kGrunHyOEKkpIrnwMAm6WC8GcrDw0k5
Jak8yK0NSBYqIFeRY1FgwxyFmgTGpdxch1nTumWrXeVbIe/7HjjUrEHJzTsRU4zE1+6zoQ6LRd0d
9PFYg7cKwKx15RDYwHZ6JOZdylR8I/tHHJ701TJIIFrC3QN+qBZR1Dpwn6OdFBLhLJVRtOLjfp0l
/bRlOgFxL+TdqWGa7/gKnfyvovSUR98ZuaXVFC8qS/Zmd0hTvOw0SarkDDP+6u5MJNgEcgbBmqw5
5ggVwCiJrg37fTwbVU+3f7SIB64PsoeRupwbuuRGBK5KKwukrrcbiSUbmTI34m2tWt6CMSMCauST
tD5wvIDmWoopQmk+rHUu3jeo/utwQOqVeLBFRT8BRD/NbEuc9M+DFBplvC4H3mOtFnwlINllnmxT
Lxh3cOEkO5ygqgct8QgnzDgEp7A0QKAtS2O8vxPcyLKae1/7Te2votEw55BtBWx9j44balSwco9a
j8igtwN1P4hBA2S05ubJu7wqJpvdWOaPiG8+pT/vV0GP613BayshUQTOWii3dICXnhqhK5nqoyO6
kcCVOK+ONzMANiKlkZ2GnugQW6pVp3ZF+9lVzMWppzPVMQwLArySbS4KvwF7gLbkuGKCSnbgkM8K
R7phg2NWj9joAsG8NiwRUtr1Mvad9oyBjINc2B8cZ3zx8F0U+gVhRymkgY81LHXesu+82ezuS2cL
Hx9lo3Lk6lYttOnLpt8LD98KYzGqFsHOmrpAJa+bwaGexSxnOPCgRuB7FcdsQ0I1ZRKrZ52TM5NE
potegGjr8ynzUoFkWTUzO8UWvwC2ZC3jwg41XVxoIvtfrKhbev9QsBJuT9qkDkIkXK125aouAEeh
SJq5FSbRCcf7kR87NLvSj8N4IdvTo/22qXG9AieCb5E0J4uP9h514LwHYxxiXV/nsYf2bEmsKjyX
OnSzKR2grgZoxdKzs8CJVS4PI5m1HtU2+Cq7oUgjyVed6lBiNRcN4BWdO0gi5DhirVtQAgguQPxc
Hctf2rjw7eu1tYOzLqnxiVX6IHRR3/JvE89+oKpPsV6jVdwnUBgqvyP+YLSydhfRT/l3YfR/rfYB
Q7p+dix7Vae2PGMe2e7Y2Ss5II95PRfQzzZIPc0g20OF359kcXLuiE1PhHl9zMJVHXXxJ2vXBFSt
+ruB513oeNzqeIRNBhKrk83vDo7Hif5SmPXbPoNNHD2qMiDyLbHosIA7KE0cLbmUIabLIAxYHKQ3
h0QV3Ha3f9YsDDG04WUwp1GWT+DBoJAuUwi/uRps8762x48yWOhy0XNCqCbNodav/GugeiXssEOH
YNqY3M6+chLCNwTuDEU02MvF39xHwo0RaPfB/pAxoTzHlNE/P+RPZaBUMtfyr6fNrAo0h9hJv4q2
LKUgWfgl1BKeBxGuAzuQ6yptVY/gQQY6ksp2KVS7OmUTWVYDz9mFAAYP3g1AU8l6GmQbbwNfPqQ3
9mCJYPGMgMpbsWINmluLiUDz3ouwhusFozHsGOpl7tiWNwEeJEc5+IQZhVx+8Bww37v+WbY/TgM+
jtMfIx0L42t3sACbujm/SSTryR+kJbQ1btx9BC2ZUTsrPr2fpAshG5Ao9TF3KYLXEbZ4JtdKfoEG
iJ+QfnTt51v4Kb9/rKyMMLNU+uIloPnIZui01aVEVCrrGvTaITqvzhhVqxjgIyplftWjY6iGDqpM
4Rl1HpiaR4kRiOOR7laKy5dX+goDsiEq8e5qOb6zL6Jy+81PM5A9/Z/U9z0CM6mer/X1YxjVZmyy
hJT6D2NiVMLvWs5EuuEalgzQ3TXmWnTnrECYQJkJsIqgPhf2OGnouqIc1BwBSim/mykhdmOYHOzm
K1rnl/GezH2+TFAjVFY2o6rCdVsYnTe+7e/echloWgAJ/Lfwsev020GcbsAwL7F9LX0bJLbBKKVA
i4FbWJnO5iAMY7gUvVr/hBd6j6Ikjhdgxsfr6iAhH0OLnkHDbfA69Cn3VoKbhLssFzk4cti7kQcJ
Bt0CjXM2sj/cpRUrMQt7AuiZpgj4KucmC3vEhMvMg9nX+76w5yJT/T4dPPg0EsSJk/bZGocwvSft
DdcRHfzDVQCox2vkpOgBzL4rQymfZkkygJZ1WdZv0ZD6HOidfjvlBGQI2wNFAhTGF5xjzO5e3Jcs
M940v6C3tS18u9xxu09lJThX7aE1uvlMqqMmB9mBCMml2VDNde+hW3u8KPEBNipLZxCzwyLOv2d2
TaapDgS7wkG2A6wL83jXDfCd0lgNBrCMXhpNLdBN0CLoufIlT+kgbKhJC62xMJsjQxl0DEI59lJc
UzYaAo1mHWqUxxrfMeEQJ3GyP/Ofb3+OnxQJzy63Y5sexqR2HxT+536crJEFnShyeTTLyaaD6G4b
FJDeG9txdNzzriq9rS/U3EYNmAJqtV+VAN7Tckb62p2hqGTXnR8DpebPwJcoczZNBD8JgLA4PP1p
a7qcAq37OImXs8F5X8YfFxk8JhIO4u/3txnsbMjKgCm/vNC/AD6Sr9Yq9b/mQufKsjWorrfew5Ti
tiwy8pm73DEHo7YTnQL1b8zQG46XciQ4vxvQF2RZJwzUZNVLhdNt1hrIQy5f1BcoH2HzU8fVWTQ9
QsRuDLO+zhzXlBhA6HFKxHmsKh38tiILrnVuroylIqRe+gnbI5g40CVgmZrOxTkMmnwqz+gIcc+m
ke0ClqxXr2iBcTIlMiejSlygED/kZibZ1le6fC2I6CFNLtXkqLlzLnLKkVQDvgQHtN4nBGfEb4LB
VKF2KjTtREPX4Ucd50lKmBuGNmpn31lGGEjKAqGU48zQMoJSIm9/GQueNdwKlABVTkhEM+9eZcdM
BRdrPlGOfkPfAP2Jz2lTglbpZZ0Y/1lkV1ttXaIb0hLJbKykCgRa/vsjFazBqH8OCNDZWdLXHtzw
8BPeS4E1PkwGdjPtfjlaYX/pW2RJOUuyjYayBcYUGGlyAF3ITAJ8DIO0FlSNlBWgvG2yg1UYi74p
FDSETgZNVRPBKJ8aEP7GpXludNn1QKN+ZwhRQDc5XvMu2fZxXl+ZcPJdDkdctPAG4+0vWLs56yMZ
gu+AlHli9tKFIBwdplS38IFYMGyO+CyLxztHeyuAhiIoGVhRWDGacYN9eA88zqkDNNCVKAWMoNVC
MrAI5cnMDjayG3SsBPX4rFFPAG0yZ54bqg6LwdfLrueVd01V0USUyii5mCOVZeIPpPa1DA9xKfcI
rolpbCkoNaZtL2WOh2WAkbxFXEe1+LzdP1XbVxYK1ThPfh33xiWbMGgznMhfDXBr0cZm3bJ22It9
L2jfXCS+lhp+CFckkubDpnKkEgbL8EH6Eg8TyO58pcAD/kh9iXVyIPABA/wWVCWT3iD4kLX5XuoW
+vBQzejo/qa1K6fXRVzD3HrE8b9YhnSUJpSTGcIyjeL7gLasdY4kUE3GQyWOuh3hdoC39xGnf1dF
uybB/cQpxnrawWoIHadCy32cZeUxzatoouhJCSjD+wP+BfLNG+oX+MaKtAaAbQxAlMM77w7ht+EC
8F0YsdPg/WrBQrNlcvo=
`protect end_protected
