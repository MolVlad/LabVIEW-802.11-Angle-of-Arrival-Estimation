`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T+AYq6jdTkwmnYnYzEwrlmS7+eYso/KKkvXaM35sP01c8oOaHMv6MfMJDhMg2VEY5mfkegP0uBfW
vDLGzYx3DQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GHSQM2Kq0tQXv6iGsZq8LvJQ7hIMWXoYBWHP1hcl9XutQvTV8GPEBc/FoMbD0tPqZmtSLey6cvXG
WjmzESaAPtIbWAenZmbzDWl7lJQ0J6p03xqxF5WpV4pVwgeFUpZpbAyn5f9vWoobmPxJI7HCfVRk
RRflNdDAESktMUYJBBc=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p8NehnUSA/WcV8CLI6l2P4VQPi3t1SLEYPHUD532eDsILRUgdPzGTOX1QThhtBWJeG9LqBBEmqAD
aawC+k4d2wmRyYro2vekqKEFhbs4Rzu6N9zyDHYeAQ4ApYITlbACR8m6a/9BIQvFbxEff5QFGTOI
4UGRPZivqssFxtWF2cVptbx8vKg+vDpCdJ9nDD0dA5YoxiQLFtaXlyFsHq9MG10D/bFbzhW8oJXg
5MgsxPfbEqXSYAeYvnqsH6MmjVGfT6ygBSQrYizT5UtvZPbn3iauKRVRme4PyFt9jdYNK84lSU75
PfD7qRBaKWrty5zrn1kNZr+goeqgtWwi+z33jg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VgV8zSUJkZhCEAy0PTNxsP2xwepZb6TGSQBWvdzqr4fGy4wRJaNzGRivGYeUeqznXcqW4R4vqEi9
rSCY3BXfkMjBNT2tDMQo2SRgFCdJ5orNbM2qdhLXDxjbuxll2G/dunOAXsYfqT9fyDtN7axf7GAe
LWB+r0g1usjtxhj5NorvN5r+UXUkvoxW++n2Ww4dyKgpVlV0BGvDvWioClR6D/T9jYsEfWwQ7fx7
cMy3eMjomxoVfm+MY6PNl5weWu33b8JezjUWz5Pjie4p7dET+WbMMBZ50+3PQfLfR+keYBrjoxoh
K4Gsk/WuCU0Nl1Ri7ctRb+SjvNcwRjobQ5BRkw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bE4aP6BYyj8zPr3jVkLfUL1s8q8oI1b32n2NUwJpYcvjzDEFN/l8QTe53ch8HyIvFN4tVCwpBevF
CcrGZ9kBaeXoNyJsUcZCTUC3lIChRuWuPmC9IA6ax7BW8Dl9dGo6acHrkDJteULKQ78jUJP2Znza
3s7sAY5y65moq4mQoZpL3jBHXb+pi0oHwxH573abgp+k6kbOeN1Rx11IYqbFL0/u4RLkHhyjzRkc
Zcr4wEGwVLrfm7ugP6qSW8UBgydDd2SiouJKCe4UOgUZ2QMu0IwcJJLhdi0S6pSpty3dkoKxaWWD
NW46tj9VQhFuyElVXRyTA9qeANV3I66NaH1GlA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jCLqFkVN6hxBPbzi1lbz7a70e+1hEdXrcy8I4/0KWaEqDygl4NI2FD3SU2/qgr605SArxqw21T0H
xH3aj8O+D1BoU60gTDAf5HP410nDyFwz7w8WzFAvdsg/r5JMfzjhvVnQUrAkAushF4HDe3auxPPK
RP0oIQ8eoiBEHiwbIq8=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cxvvzfXfuptc1Ki7wNMtIsbAIBiNxcofoeNcpl7yQCWTin0ao7pVlcc8vp8Z4T/Ohn5V01A/UfMT
0FzBilFbVAvcue8kCkNqz9GS9j2iT3vmR3dqzs1EEP9ge980sfKsTlXt8huDPS8WwHqpim/V+5Nr
acDN0cpSCbwfyDpECiMh+h3pJc/sTde6A7SANSkXsZltS+OPuN7mkINbcWbxo29sVzxHeQ4lGuL3
T4d7Y2ZWyqQIby8Bbs/waKQqPk7+Faf73d3s7nZfz5HMxuA3k97CLo9jc9kE17fu5aVJEx09Xl/G
Y3J8znC04I5VwGdaOdQBs3MHsb5S74vCnIIC0g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125840)
`protect data_block
SfYr0kFnzUhc/3Odn0519lylTuIDjHRatrJEJEmTNjmPESoSik+yPtZzPtJCSnH833uUHxkcfjEp
guEchf/6/6DHsA14ji6r1vtaBUEhwD0nLCiESM28rgDKt3FkO7KN0BPvOlVBQZnRl7eHhfBfRCbW
1NJyO9SoJ/jMPswCqzNEkUCxpZUM7YE0lipgSvr95mwWhTTJKTqK1wBUTW4zbIDWbCq3tOPbP8aL
NqxS7OStnAMHTq55d1Qe3A2pwx78ddXoECuBhBa6ifIcFN174ZY3gcNoP9t4CJ9d8r/LvyNGa0sy
V+KEsD5aoy/pHtDUMl9FTLJ7pzvJoWtCO27cRfLc/rjxzH36QdAwV9dn+ZTZS8Xh1BPg/jT++jFR
ncNr1CwqdZzw1zXRGHDuQSZVBlmdPSqHgqoZeuaGCkkJEN4Tw3T3yIZpzLijxpTGUWPuNJ/bApvj
sby9luiV7FFeOXMo7jLQqxivx+BN1j3cPk2bBRA4tHU8g9Um7XfvAR2j3qBnq8pSi0ew+Ohp1W3v
EbjtJB/X+NsHBpts5iOnC1JlZGGjAg6/Ko+eJEmVKNPNfU8MwOl6HjUoEtKZrqEHYWt3aCLfg3Af
wdXOvsdrFmnbHZCHINpivFBrzrYDA+F6BPuVgxy8DXNhBfPQBBP7k92oiutqMngJ1MLEwxFJul1T
VGzlAyNb6nuHn9xIYvaQkEvw1mxpni7D6jt5EFvuDMkpbGpwPKFvidcjUGGm0AGRNDaGeMeH3plj
BtIQAFqssmLMNln69DwpCRcAEEwOILiKl1ln1j+xbqRo5UP2oNJpSrJqn9tGUKoerhjKiMVhjCvd
O0YoP0ExaOyK50g7RappBxpqnIjC75jvVx71ILD2/0Klq706EQ5JMNczv7G6aQ9Xon+pzPuF3KcQ
54sR03MVWfmNC0RqCei7n5fPyHe0d6zE0ktNDURDW8VN8hRBpATSywFqdbBq43y+ftZjwxXl3F4r
qakpj34Fc1yVfPpo/Z5BM+wVHIEVw+XtCia1kuz7aMCSsTrK6jdqHruSAHPyhRFn1AcEtd+ETIQg
qgiLDkDkkckzvbP9aiT6eOfUvkJ/5jjLHS7zR5R1ss7yVB+h2TsVLivyeztcHNN7jDCcJEZVGj4M
w1ORN4VVp13JlQT1L6Tl97d7+tD4yUq4YReHDwBJIWn/VwBffJRU+ZFcwdcdEgLJ9/WPtvw5EpgD
wnkUWFBfL4gGNcxdaDw/39JKJtLg2VDiaPLjZuv/PQN3a9Zk7NB+FECL+E5ygsujCjGtmWyAy5Xn
bnhdsLhDPZ3ElmfT1EEFFnI/B/fR3K9djtdPQSaM6M5/nrUqWYMytqc1XBye870Coc5bQ+1UwHpp
b0UjRFCYmzwnXMr6tfrkGqaj8+5MWuCweRCNitoxlsVHbu0ZrhIEQTJ8XS7nsQn8rgE2g2/3iRfY
hkiarbxtxvNGS73fhHfGGaqRLXoPNaJZ6ezYjn0ucKaUBt6TDOrIaMcv2HbXT7u5Gufc3o+NeAMn
M7qio7gPGiGjV+n0cpjHIdQU0gdj7TPvCtjX6jmHK+5eMBCex787UuLj+f3qNtoGWOWmE4o6CwYd
lX2NZ9j7eI8X0KFBEPz619MvM8nVspCTMHJDCAT2yCecKq1KX99KPFCWGFo7UUbIvMHaZ1Aitmzl
oDQ/jx7q5rDhQY+OvC61fLiXmbttUifeNB8XkipvWxkcfMJMIepqdYFm/DO57JfltbsMs844OTgt
R26xb2Vt05Ge+0jVI0K1j3zqKW4lvyXKGOb6oB+9Qer9c3AEWInpgO5NQrQZkmli6RmvVaHl0sKw
w8YCXph0HmY01g8uzVhVEvhE2g6tl9tNE+TMacWMdPA7KM4cUbrQp8Rb2kApah8ZAE2ODbB7Wgx8
8eRY1LOMYeDqWAPfVVzZNcpBwHtFmN/3ig8vgYg2jJccnMBIccqqOnQDirYOEGOIkckeMLRLJb0A
zArsiV8iiBy6pmmCbNxs2EMiVjt36abA2QOTHUjn0bRQnc2hlb3nZvEFd7ULwoIoMmZpb6mYNIXL
Zb/6xgv+82oZvNH0606G2t7D22yWt+nIhb6jIQQ5QWinOS/H+HijH1c6DYwem6+ZK0plchVY3Tvn
+kx+CKVpUnXemJrMO3/8MQ1/G5x6TvEgHQlsVjkFYZNZo/kyf3xKT+qMvC0YkXNNK5tjVHKaFPNb
NfjOd6nyfu8Qax/wfbrJcaNTtNIX+BU4ILdE/t/4p1iSn/uGKaw85H0jRuA60dGX655vZIB7324+
7GD+XpqtpyOG+joxwvRkhnwcjxKXx7dScdk+4t130Vc9TiMOGlBngFYAlw/CfB3GnpoyJWKpXXxR
xSvAd/QNje65paZHB/Ue+ZnHO2+qP2uPZzt12MVYCpClc1zH4R2LqrJ1bo4qAE+N2Kv+Ae+jy7Nl
96AVgeCSvFgbQXOxeBdvKit934pg+Uc+Q38MWxqjx/7nJNMTq74DrxwXol9EJFPrZZK76ICcBMiQ
ylaSQhQS6cZWflBFOqTS9tfvA9neqYKAF2XTFQFUfB9Tpoaz1fVB2ivD61j8+uOkdvDr0xZjwudo
G7pkgkWxhOE9I1op6KQK3Ll5Hsltd9zrfa0htl+advcfVP9xPbO6g8DekkGUGuHnk3q6k1ZwTRck
YZcvh2MDoa9hpGchF+A4WWJVXz/GT9nDOXLS5i9dNhW5ftGeLVzKZ6hO6gZq1BZfUgk5Qn2PXPGk
gOV/lkrTcClfzoDFBU69fz5tafIGMVNlez5ZqFH61NIxtcDUDCdnsMDT+d+zlKLifZfqNkt2wzND
jCnAoYw4as+5XXsHvG+DXjBfJKgjw1iTa8w3Bv0MW3RxK3lApAlmvDak7wqdHwE3C6D7x1wBqPQr
5dAQAh310En8+uOj6Z5hMGLZqOga9nf6uvM0wmrF2o8aZc83D5QImCMnI40tSnPs/GDVFFMaey4J
V5P1fAT3/4tze8+Hq5hmzGEohJTe97VeNj6FGmlHfBu+aqjEek6zGv6elUEvIuQMtdWXYeJSSUtx
gutYxpmJgjrZouEQpkAG7quiPai1zTpl7hQN18TqNgJQwPC2mGN5goK/wLoJWmmHoO6z+PFY32jn
N0s5QvXp23inGaSpK++j11O63F88ySIHBSrzj6kP8Crj+AWy2O2/U9s7woqN5mdvw28uMOhX6VfJ
phYipjGE4jndTZdoLdRpjutcST3lQo9MA8fV8sV7YeSzIylGCkaMVOFZWEJMcqN8t5WtT1kRHDfE
mrC1Pa25hhhBNeNQ2PzbOKoz4xYQVlecReXBy4vFSsU1tk3voqg5gJAZB8g0oJ3vP2TXL/Fn+P1w
aC83k7z6WZWqTrtvfEGHec0nAk+0Gy1E5W+hPWS/OrNAO24BHe2MZa7LQ8SuUEzubKR6bytz5R7b
uOkDLPV2ySugSCAZheBpEZXUbST0Wmk3dkvqB4269vnLYclLcfqdpPxNvgUhGWK1GB9lYaSQbCfe
esNSTzE2ACFG1AMyMhpKMdbeG/+TW7gC8g2VT8GtSsdV9bL8tOMouzqrVrreplRACv6qB4Oayqyj
LI/GKcuEgf9cFksiCnpei74rRp5NdM0F4LbM4JpEgfuDqwCmC61uCthpD51dmfudZ02bTU/DSQjj
SY0lFTEPWcIWm0AAvUhVOV7qIt7WEQOxG5/+JlJrGhqqiNmHgc40G6Xt1w7sqs+g7347NgJJpVVo
NEYlHjODnMs7IOHFpJX8tWtUc7Dei+ZrXnIPt2a1ukyFwjZ5aMtdv+Daqk/GznExxCu9qz9FjHV6
uH7IrGMvD07SddRGIGSBfuDEVh6Sq+XrULwvTCIaiTErBmu2nvO39lyGcIcCioPIP8lWb5kn9BJT
TD+56YXAsgeMiolSLdr8tnke2JfMhlGAIw2Lof5h2kiwcz16/eJ8WPwygIa+dPZEyLqMB3vrj7Dm
pVoWUV2NjWcAHRCZWW64ESVXhTbtVa62rzycI9l1w8HQAQKf17xe4cy0JhlOpvlN8YYWMp/Kltag
ulsnlxSkaOFL0p7A9KZmvX+C7o2Fj8WBsevKWUrly0IMDLsaBG42WLbBO6N6TIglX06Kda/WUzA7
P2qWfaLTVhrNW5lCl06+nCgkOUDsziw7Hz2LDULrQ0eUHsd6nq5Vq0KavdUIsodbc4gsrHbnZoi6
aRD9M16nAwSJLu8DoNfdwvUtFOd/nccBklVZs7wi9R/6h2vMsdTksqT8C+nsVePq6dRNMF0zEvtn
YfQ9vUhwvEVakIo8BME0mv9N7u+0+My08/9RYKyycJfNPu2Tkv+IlymPuTzlFQkrozsJrVeMcRXi
mYGqXdbOwTlOmS2s9bAl4nSu6jvav48LtS/XaCXIX0i67IdknjwX0uvtmis2IgrSoWfNwo3hNY1A
tH0s+9bwdmJH48oO5Xfp3wlzZUATQh0mpmbRqe8mApBnXrnct8fnoHVau/pMeeDBODjqNTqZ0DPX
42iY2gseM9tg9vYEILWPQ2o4iB0/tLbnwNkaImLiB8M73y+iJ54aJHet4UTbMexsKVU07gDDrnhf
KbrLUcP2yEm/qq8Z3IJNQxJBcvNF8d38P4SWVmdyMEHNiBGPayTt4QQLrnaCOF/yQUkIKTi6ljy5
dq4R4cvg+OOXkhfEw0Z6NvhhuWxCW+oMy3mgjdnZ430rPZTubjvclqoo6XW9bZFpkUf5f/81uKR7
KPcC5OmsN6tYAOM2lDWx4DoWg9LZrD/SzG3U+6iEfuW+g3HbOK0w5It0uURNiJ0JMz0arxVYM+Hf
cRw/LWM6Mowg5ye07JdRyN09EwlcY4HW6gguv5uGEvvnbJt5j6E1k4VyNPRJYq1SLxSDQSqevxu5
MPsM1p39Ftrf8D5CUpoRwlBeGuRKljdNIy/YCPV+IbYcI0zAGTy5sAek7tK42MtS1dMLYCJzVLhh
7aqMD0ZRGd0UgfLk/CQQHgr3rqtkBcabu6/xKlPBJYmEu89bKzYH8uSJNvN5a3uYMKekEmeRcy3B
54yhhHh76un90dMdRPZSP+B5V9p41W0kUO2OYQArZLAfV88xDgkwLiY+u4JFL2zSf9fGl9SYjPhh
lpzx40eVRGxdb2BdGdxaj0HgonXTB9ZCtRQRbXLm+/FY07Gl7zm0sXptntHmV5RXO7C0sYXd3D4G
b+4uQ4CFvq6B2RIGYCajlpicyExb9HLhP4JKbCEe2OjRaYL7lnJynlZYAc+FgduzGpIJN+XtJpgD
dLyiydLpW+1hA+gmq56dF6qcZglNot7w1tqTv1NROqMvxud7+0BlpOdBGs0KnlpMWa7Z3sIRIMbA
cqTN9Ck8x9xvHHwhXrLiHUdMSyReG1N24dGUSVraSxF6SiKu2CStqFatvFYngokkUEG5jkFSxvk8
eiBp7t5niQgl12KvlfHIHemb9OUIBF2n+RR+4rrjdOazRhRLGx8rrXwPQJC1YfQTpHzT/k+OX8c5
8iAOCe+4VxXDVL1/K2d4xb8WQmwtN7f0xkQKq+91ncQw8BUZMCI07UmzSh0AO4wqi1YxojXixz2u
kdI4b6H++uZHDEUIeoazGX3UdDxU4upAmYiVZDYLVfrn6jQ+D6i/i9MNkQnCW9FUtZgDP7FeK12z
vgIjI5OdtkfysiqygKqWmtRgCkKGUI0G/Fx8eNBApguJ53p0ptrvnQoMJr6OshMSlFz4DzwmPSxv
JpDo1yCIjzEHxwftmAbDNvDMhuTRYQJMn9LKY5ctqbX7zxOkFiYBKEEMXKcg60oTZnT2oI8pVN2E
slzb7gMC7QOKGgDau9SS0lJ9+gV0mRKQUusufRBIr/GYOXoVBDpttiaURm+a4Hh/FGUxHj/GG/nV
eeW9+q9beqdNJLjcWgnnFNu97tL7rCkW1OVvJCOOqydbhZUqDReY53QDUb18I3qKMaWdTUS+e6Mo
Py6o1py/6Z5ssiYrBggOecXR9d+177wBQnGV0yLwJfTS/9h+Nwv5EydKLSNv33UQ71K2txidypzu
3rOGN8rlnk5e/LYoHQVKEWdx6ITkGVqkX9YYf5CLIAwHkOZvHKshX8dkmcXMQNs4KcI1bkj6zpq8
vpdTqjz/6JzUKVwzS+rQGh4l8sdkTT+SRnb9kcBJkz2fL4AKh1Ths5lXyXgtZIofN587vOYYIfXo
vRlp02npBf8Ni1y040Rpdfx83AJDw9esObwfc+RBXhY6PnUEIMVnvcCoPnzLqRgT6TWe4QSRdpu8
xQPcPTnrKWqxxwpeRLRnhjcdiRC61Ax37uPCFDAqfuGYfo4+vOTA4nhMjKlZAGH9ZSNjwc16BMll
EVLT9wR5Bk2/TtAyuoV9VfdbV/EFc5YQqChAmTUFQVybTQvH9vFRGAHlPUA8xMk8GTUwJMbe+mxt
OzYHGUvze5jUXsos3t2ogQgVbRYxUUNkmI+wf/dZMqqo7jT6mkkLJziuEzZUT/8zxdxdDSd28GZj
I36viSQKMSDtuqJeIkrIqee4fuFCnY63vovmsST61HFkdh47dk/bG1rJOiXKm1c5V64UaKvaZdYx
boBXtApA7n5yTdt4b1/w881WuCVP2+08d3SNm5fIlTayEIa3z6MNswFnE4eAJMQdyJYHkCQ1qn50
EgV/EMPkXU1hAshOrko/wUfpr83GMANSZD6ZYdiwZ7PiFZt6wkUrKf0XGZv48GhXdjl696r9A1yA
MI98JaAANB7oVFBlJOpOJZgYfwxPSTMc6VIqVSHnYG2Fcc9Ceb2txFMPlydggu8pF4Cup2+88OuF
FHMYlPbo/homSlv5+GREBURy5wQispaBPwY2eNK4u1w3/kNHkXfPVaiRFgSMdSiU0k7KfdqM45kb
vBjXIP+/eWxzm2wzmspi+PFdM8o48EH+poLNtn+NXwpS64QAOJk3wqVHy1BQNeShXUUOr7X4BhPx
DsowrlrrueVSFtBFmFCl+BsKdtf8SMt31496zw0rrfg6jQ81a0nYf0DYIsHSzhxhfngI4cCoOzRb
fAEUkg2XDJwa/B5tvJoiKIJqEW+KzMcDonnQfLedNoDw4/S27FBZ6hp22DlI4JaX92kyiHCkCwlm
1Zl91QNBBTdCjaTiGXlsIQrelGf3I4xib5hfOn4Bo9BVIBYj8Ppy2JExeNsYOtdcG9geBUQD1SpF
gFr4pkJr3jIYvIbFbTz7zb7y+dPT2Xt4EVymLbpDF1NbGzyRDgWi2ZDtGh0oUkQj+Tx2W4tIy4W5
CIprJw2aNfjKkBSQmil6oslOYgHBtZBxvmKRxx+LWU+Fib/Gtv8iYIML3qB6m5qwKvRJqQRF+y9R
5dnKUi/hfFnsg6E15dqoHLAYw1UYofRTveNYEDHMTT+IGtCis0eu9QWAgi528w1bZZDD037qpIH1
E4gV/HmSG4icEt6/w4IWjUhebMIrhBQfvTV6gL33KjJBJhjJ3I4nMhRImzF6sfl/hairNEhMPKMY
BBmQH2V7WgBrBfQKvNkFGKjDVUNTtxWUPyF4xTSDmu1Zxxy+Gt1a6nNGnhj4pBFdOEKgD0ONXUBL
NeNb9aYUmHGNdslaAKqOGcWcc60hVO05TbjMVbTmT30FrqbSjbaPUpB/dIZhvLsFBQhOv7mdTiCU
r7lhU2KhdIySSA/sILim7XJ89brB0KLcH2K5jCHfTRetjITloC6n/S3LztFKxszzQ7jvn13FL48+
zil7e26vyFNZbScAhmPh/eOEwn121sOxFaDGDBWlkN1MwnyThXqrdio1sFd5nZ9nGJiL6XO+unXP
UxuBN4sugq1H4sWwCkaF9I/mQMUHdH/+2t2E8djyit7Lqu5OWZY0ICAPSnbf6AaLyoEapUqH58Fa
wJ/fnY4sRjnqlTViGK5WwSLmfNufuYOWT0QyodVM7dcOw3AMnLQ/ssOS0m7695tYBpxlf8FR0bq9
QUcBXlnQeRa/+IRbbsakhL5enK05bDw4XEGTuLRhAlV0gKywanP6QI1AtSPD4QFx9LzaIuNiX6i+
wVptrDtfaSnV4F87C1m81vnPQvfctfiLAAcYhUxax3a443JjxklOV2rpub3sZvTvkWmuosIwn8bi
YslaKi9rdaFwsdYosKhZibDn1SLnb7V8jByjVE3wzYPe5U/NwHTuWXP2Pgnh/dnGMFjoZZ/PCeTu
TojTaiZRHtDMa8iIaSGuLkCSCDHWR6JR4zEA1aUqg2JOB7pTmZNoLNeQOKw4Q93iWb5K/lucQkFV
fOkXpUnPy4itH9hIPWO76aUYFZbF7ylA59IiHNyl+0sVyBKcbnc8f4rtrncTB2pO+1HwP972yLDO
SuBNjTmUM9wT0Pn8r3WIjF8EnnXnXDYfMbyYVjb4X398KMAs95kgRG1qFovvF8J+a1NF0seuyeKY
6E85np4bhThqdKr+fcAVB3GGd8aFPNmlcqqjFJ4zuMeFt/o/ec/I8wHnnQMzGTdGBqjeM5sg34VR
/hc3KjjL6VkyzPhfMSGLb/d2TuR5stjNczMivV1kDq+drQ+2OIWzCVrkjkEodul/VvyBxOwwRPrn
d8IGpi2z+cqEp3djm4KDzx7cxkUmLXx9/yNRHqMl0I/XwSMQeowXFJoiY8IDAtMyGFyL2n/Cie2J
Z4/s8dQ6beO5IrO3YoHATTU5bqgFSuT6eCBc8ncOjyh6dRqFnq85sfGYrA1UJifibLaekYFhyap8
h7yL1h/hkhsJFxD3/QBgm3c4yiQCmyVMwFCCUGI2r3x1UZsj1Doz+ATzjbHQ2N/B+2I7gY6KNCeG
5TbqUgaSEMH2AiAsemYrhIRq8Xc8kEyetlXyv5sjFfHUtUQI/VysA24a9z3iuGFFhCko+CGClMlc
wNhtls+PKHEsNsHrDPB6jttYVYs7p/hNug5S36lRuPgjP6AdJARuANKd9k93MDAyzqjWDPJ0kHZh
CHWeuu8a4NhuGHhHr1J3xlLrJGeDu1nJXDTqI3BAUSw7rdiTaDl6PonEYnOgXtTVmHYG7V0c+BdN
Tb4Fa5GEP6MlRsreeL4KhUToB26AO5uXBjWXvhxOdYt9GI/8SZvKf2QhogpKXFsEyBkXobfiNUV8
knFFR6j+kwehcTwiplhyJF1ba+6wYFiQ8yMm+oTIejZfoGiOojHetQU7ENPRfoar8V+O9p6wmjEQ
PMjiwcrJYfBZuQxMBV8SNP2YweFLMnSF6rAX7NPJZvitH6LlQ/vHJZlP8ws2Wr6biZet1wPZd19s
K3RyUXtdNZTC5ZZ29nGX2BjD3WluSWk/ei6oZeEgC+3APl7di34MLmsCHyD34BX2qGNdeO2xH+A9
+3CSqjDs/VrQt5gJG70HE9lvH57kCwtbVj7J7HnrIRdAaxXdDFFGxhqX5u7Ga14ONvYR2E5/YSzf
NdBSSLRDkMAfFbfLbRmNcn5mFQmb1xYzSBpBGNwhUQVPM4W83dFY2+eo8zlpmBlA3UM1Bnw5CGsI
DI/Jmy+OfjIHrkn+f/b64mmz2e5kFUDHAi5N3YxiIHALOz8oAWU0L93eZpiFpPW4MHaL6RLkCq/g
VV/QJRe+HnSUJuh8adcYtA4xUQ9H1VWXHq45fMSxj9sdnhyMSHQyOuQY15YWCpGcN/oUZKtqmu1e
LS5sM/8whXfixeWtwLPe/1l/tAhV/zRqoGSXrbIbP9WrNRyfPYrdK0uao8P0yr/D/aZhRKevKDx8
e63tLzfheby6c6OHTsH9BwIvhS6rKCEEj7LqTPFlVpbXSHkCqggPmV27ZkktY2IbpCN+jjPuNSpQ
jP5rSBFwbDyA2Z+SicfKIwWgT9vdt5hrn+/ODAzOruyxDGOA5cWtGPtIzbAIl9dVrZY420a2SxzU
eTOsysL62k0MMALHucLAD1u+LPlG91MiC0vEZZiBFFRc3yo+cIqVKvcRx3MzgCbkITRYTSlcREU1
WlEs7imqlFGiSgx8CmxZ/PeFfjz2QTzt/c3LDrb29eIrjFY+eJBEpSY5MnEQ1qT8nDytE6q0TGn0
7rIXq25R5DqYrToiQQvW6GdJE3Ufn3RXYsWg0ixGXljVYgB4mzzd51Il/9eHqR40/J/9A21izlS8
1i8H6knuVw8uXgB+z5S0xsYPX3xIMRFFn0b5N99aFbJXXjBpxzHQesQt0GEtM//6tHlsyD0RiJnx
R6+VUCLE5034qFGGDUiIliUBvB/KvsTN0totkf87t4aVd1dUNCkjH2Dc/wCmAPmZ3qbyFvA0HgiD
rO9RKvKWaP1aP1XSLQtTb3bXmQ/fDvCUduXx3xyrVGFnvm5qkGj32N74SVwY0WG7Atov48JQOhkK
oYxIyEVqAsBTru2xsrjjANbAWODH7GzzbHr0CP2R8xg8Qc9afcUrR3WVHP8bc6Kq4sSmZkgx47uM
wlqP2RQgyVfc2K0D49PTwFe7iRnBKFdllA38LrgBtFD+sEu5S47xdML2C/T7GgoLARazoBpxnoWW
OsIghnen35HuwEWsQmQixCYXucZFwWpvOuMd2aEmdlVMbWpUz7JKHrFlbFr6fOr2cHgfuDKSz0OW
lXebzyuICuSuldOSMYW+0o2eI41dazVvo1qlUIdUCil+kwTRo+VTn3/kxczQkdPVS9TXxOLTXu70
w85nVM5uGH2v1I8aMPylqTxRV0NCpC8bCcbnZlgfwCsOvfkehWv54fo0O+WwgJMNH8PfOWSfqKvt
f8hTE8/YnzVGw/fJx5kV6nMNuksO86Qnb0A2NBfRvCZO8uUTI7jTcw8MTbadBmKc5aNay9RZ/Xfm
6sye9gpuRuoysvHkysaetRDsJJ4pgcjGBD5v8z83ip08DkjT57zreajBZl8HGhukHIDilvu8Zg11
9RMIKPteJbaNDCRh2qqsB3d0VXLLyQEojMOMGTsVZ1RUg4So0Hq7Ny0Qn5wi77CywQ6IKKbzBnd6
HbktMsZTXtsbe8D4SA5AZM55AcQqRvbOLdDmY+zZMwpIYnuWRrIzGbCvXuw4DE8iqU4zEnsAVMkZ
/mRJEMtMWr8PXJ0UMq3/MhKaT2JR1fw61PAQPWGLEWStXFmYIWPOCmq+63qz8I1Ng1EMcsUdqXX4
nRFvnUdG7LAGgeH45CUtIwIrRDvv8YwAj3fglUdfuJ1QHYruK0kpGB/z/u5ALbKYxE498XNqRXm+
rUWGR+iiYgFy8VujVTaSaVA38p4iEJkC6dg8M/2SaTV6pntFxxesO766oXHOQHsP9psbV27cIHxU
fsca93/X4uBRr8HlDPb6KqY2WxWPWcZRG07LbcgZ2sntKRntcGyTeygPrJQz+IFjROJ6JQIReZGv
LZ5c3nYBYfNs2CGULLTw8ErrXvRhcMZu2vC9olDwHfxnNdmfk5wdAWIR7hwTHWIIWFawWdrxtYc9
Mak35QL2c1udYjfLsDhvD9AHPIV1FMX2MYKpdrfW7KZrN4Q/5IuBF6iDpGAptctgjHkwlR5yuAmy
uI3Tauo8/wEMcDOqaPn7udWWFPMdKno8nLi5g2gG/u3kGV7XTZOr0AaLvgpsks+zKBguvjnpyfnw
qPggn+EKBP7Ylho4he6LeglEfov8V6n/99TbbF0txPOEPZMObVuoBEQC58osWrodSf3khdjyQROh
ZdnfqjrlrU/fpqBnPeY4StI9/0/4ozPRnXiGARonhE7uikGzfuZVVu1IUTzFnULo5iaf2+YdtMc9
i8odJWFIoB2fUDu70xT7F8fOOOq5uNej+Qr14jAKaO1DsOIWgIbUq9NcCLqmmE0fkDhOZo/dr9+C
OerNEgbdts08G1SUJDhruxQXzns2HIS6Hrz3r8CCNigK841G6DUw7m8PANw7y2MN5N2cvM0JiWao
VfO5xHsXiR4cHygsh+e/01kPDM+Y/l5AKMjwoLF2fjGeqK81gu7HPducWkX+CjyitwDXT+2YVEu9
0gpqhPKq+MKZawNUrrgHV7xpz4DNU6ND6WY9+8JH1fLxIoccdjJrwxiAqhEccTi29jv17RtMcft7
EIXALjGy1Gcz1UXvu5XKabdzqhRXFNb8dH/T/GRx0ZgnWCS25zXlh8aRCr9g2fIO030/ocNgdvqO
7GP3W6lyFeYyw8nAHOhMjk8QFDTy1QCfocgt/XA9TqDMI0xkZWZtfkxmpeOtOAjv5KNM3jRT1o+Y
77DAUOJiapn3itCJdFoCFHTH9AdsJN0dMokR6g46j3c9ber/8QxKeGSTP1GI3tc5MzpTD2kkURdw
efAuzMG9bJ8LWcXH3ugL+ik162WYUk1bzslV5hCGEeWl5ji8r97c7SCcWzKrqtqUQ4DBeeqDGB5h
FX7Jb0sZi450pJJP1Jx1ZuiLRUUime1eEFx3NDJnD5A64yONeUmm8cyGw6ww7TrqqavzyW/WM7dn
DIPDGC4aG6Yqeg9p70PY0n5lKSaI+HkGcBZjqGHkFjuhjJWPyakJ7GXmbb1lXmgVVXs7WUMLrxp0
e3IymtuPThJ5hr/kMmD86RuDUpYI0nYRA2ZT1NH4lwMvpx++nqkuyb9iLMsWx0+clddbqZgDL/Xc
wPHXoDzMp8cCnQaUFyRqbCLT78YnX29d7IE+bYVv2rnTCc4HbYV/qfLjUAERpYGWhTmT3sWBFC2k
xf4ZbtajTI9AwznFyebsQExg5DFV4mEFYJ+OVFiLnP9T1JcOzP8ikaGb1sV1dTJUTE6XWQCvoPXp
3bqBMGWHBCJIswPSXXPLqy5fDZmLBsjvXUEjHTnvd9eQXhaD2QYbJuY/XankwLxET19vAWhFaZJ3
CIuiu2dGZ6k6IKe6U8rfg9UhDRuzVHta700/paK/I1OtwQTZDdljefj5Fu7gTV+C3Wz7VV3/m4p/
OZWFq5s0ZsGd43YCi/uIBKS/wKB3O3wp52b6i0IbJ4vgOUtVFl+hXzTNnyPNQ+iBWRSZa7Ag2tFb
xGag5LQplu0kVE/fSe6jFxvuL4/us3MT3chpZ3PK4TW3DqSFRzprHY06FJPxtP3XDU/fbYUZutXH
K8/ix+2nkjySRTLfmvY3Fm3qgckvJ2u72KhBpPOygB514GFCQGSU3PvbUJGS7nptDA2OPnIlGAN0
VT5OOtG4GdOF3k918VCXsYCaWlorfS9keIFeCgmVKurCMDQ8O3iNpIyC+bMCDh5dClqfe57t0MpP
DzD0rB8gsuYi/D4t8or69MJWWF6lJ+IM7Lo7EOBv2GkUWZegPoGiANwgJBYfej67tuOo/D96Uxzu
Zj3qHSduplyDnwP0WtVMFAqQxd/D8RY6fhzDhhW3ThtSIuipRTmicTq1Ik1PvGcLveMSLBd6PQfr
INGZesmr9nFmtSain4Nfa7tQTX2Fu42B2WAf9JkQ+pjmKiR92NnkvbtxkxxZBG9Aytgq+RD4HSpt
jV52J2pQp9/wDnX5MDjbRE7Xw6ZBBb1RCW4nHNIB6qEmA4GgW1mIJ5cxZ9ZQiZWGwQLUBRsgMPbi
aeOoZ/AEBNJErme2pKDBqxhl9mnOENtpvLBZYBlqoHVMfjXpNBAmaZU0d2BYiD43NNnCxwshzjIa
5ungfSQ35uqRwK69Oj8TtPwW0sk4D6iEbbKZ4zNcweq1ZViYWn1XClK4+mpXCwP6PiVzIPin3Pyn
anNaebGk/oO2dBQ2F11Pw2nZ+Jv1OvMqosNbVAK1McOtq2XUFg8kiOm+bPAm1Hxp5uoV2qAE42xn
W6hqOIbQeUT/Vz6DjBMQgB8nTqfcYmhn0B6t3qs0acvqmHtGL6c4qJ0mJKJEZDCj/u3pvgfV87Yy
474OIEVM3qUsL3rKCpKba/wYmteMYcYxtHqCqCd1/wqZYidTYzcLHVcfncfadboIfrcuY9tSkTJM
E286rE3NWBJRxCplxQ2jxn+c8egXj0xJm+Wlq0tBHP38AApH01ibv2FZf5utEVkvgCu8UkB2PKVT
/PvWFgm+H17V0lhe/ebOBWHWMZbfNPac1cPgH3e1ntORs6crWO0rGl39M/IWfT0T+fK55Qb4JKyy
8yr3A6pypCAFgjwtPBQI80Cc3Kd9TmUHVWOQoHupKpCe4kxEjJuBQsDr2Rmg1ts0h2A+mwm6YkcH
ItF/OVkDqRUah3u0J5PWrAb3MYO+LEPsmGNaLkjICRvphSNYQhDuT/7nuCtpRZcXGa3m4M1csueX
yJ7g2Qj8F6MoaHqnWd6xMp/Xicuxh18DXS6f1y0C681u1fCD0l6VxMwihLfmC7Lyzy2/kMHvS4Os
rvHbQSKqH0O5TIHOqg6uBhH8kSW9IojF0mJh+KBTTns5E7j3zCLDIcvzmMf5aM4eJdKHsq9QaE+n
hpApMtRtfeglmG/QCEqGv0Eb2iVoxPswtIaLqooZ33e/J/bYvW9KPQWWoDEVmXr4kao/MWAIwylX
C9MyanZvG2c+tqVBPuOiPzvPiJr9BDHf3UMEJUEtBOBiWtb1ghs+Zdgeie13TDq3IMlHHoFXAQ7l
BWc++/Zk1BZx0woD9+A8aLnese4TxScx66Q2tAKjCn2zwcmHc2K371fapi2+RMRUoMDbYB+C0f8i
sU93F68lYDAZn5mZAaOoUUEcb6D71KDEk2iqrU/5yghy2KBOu2FCYk8IIM0G2a03SnUzAAcSxFAS
QMC+OF/HXREaOdfl4s5kc8Ru8jAoAdSeQTmjX3aPsoXOWTFq1Op1e4e9LY7dIbmjGbUYUYp1oYFc
0rzK6AgllITxuOgG5R4R59+rc89wjn/C8BAmeGv7H3FVqrD0lM5ix1O4pS2hBKzH3GQoA1QlB9Gu
yQ6vqZB13PXGz5i9Aa+QQ/f9H+TwGqUczRnkKOuEiFlJ/mQqLDsGRb4K1EYxZCnELRv4GyHTiTeb
xSmuuWf/U9/mxNhJxPsaX1+iG0hvM39WBJ7dgWnj99Eq7kNmoBY3FP4+GiMalsI/6BErkhtjtZAM
MeX4d0lCbG1gVKaj1BZubW5gwlIbHX6/H5VB1OsI9u7PMIAIylQmlXXKO1bGIL8MEnks8kDM6zri
gKs98mhKfMU8sbNdISBvaMD+HIXs3nDncvwLApsgBrxxyURRqiLYgBcDwEdSR8pdL7uwv0BdDWt6
xUbChPlg1gOTsLV5Qr8Ltw2AxkTwZ3ozBp3NdaUk+FW06okjMwgnsZ/u2Yrr7ZKTdD6JVPd6xZEt
uI1Grsw+RHVNIa0i0FTEtSBYBNY84kry7um0klD3hPkwXLFeElrjY8lkdo1+Ox7rqsYk5RvIoG/U
9nIzMZBCRtrP5lu6e/Kpaw0vfNJVArirykwDse0Arup/ijIp2vJZlJGVygIE3Fws54vR3JR03KSP
0s51hbIpvqLU/DLE+wjnK/94FJaKDJGZbjt+xdKI2U7WXEIZIdeV9gFMVjxpVOIvfNH0RG+cSE5E
YGA3pEOcRq1HMVnlQoPnYyGIAKJJ94hmKmU7PlXNSI13AF1H2JLcaL4UR23kR+kmImUPs4iLgfQC
G1ZoC+fPsP/wf3zBZh8jKXVTcWi1cbdcEyLRsnxH+I/iuAP5zOoAd14c23JCBP87E8llzB9JXbxI
GS5KFQUO98dlt6cYw8tzRh16Fgyh8kdih/Cacv6rwayQLSkZkK7FlWqVgNGYXveZvYCYE2IWJs/w
KjLaLypCqJU5jb7PevZaXtCpoRKMQ3dCQ5M3oUVR5BSNvf8mlB4x/zGY7lQiT9m5onSDaebd3Xue
GhFwgKq/lNqvriKP+oVNx8leqmOFn9mWxkgoC2ztZxOCmgDhhxISjRyeTlpt/PJ2xKGHCOTL1zc1
LuK7MJvRhHoSjHztfuRQYv3YexT9H84mqWFW0lR7g3hTlCEtXA5FD5uDiOosE746NSqAk9+30dQp
dO+MCDUNEFM0qutHoXT0CIBX3nirM11y+vJ8o7POMjRhj3k66r4rvgPbwzAmEEislz58+WTEBS5K
P/dTowwQnqcnHS/hbMy5O7guJ04X97ZCAlUhe66hGC9RbTR9r9/KMJ8EtGJ4L8Pj+QdDbt8ycR4W
8Wf33mUu/VwvooURcK/hibLNVAYsd8zwYq+WGSyHpwHhtVd4htWL+gy6avAsnkb8PW23XweV6v9Y
rtu4XkILY2GRHmaQhyUuVM8nYwezk7lVEn3zN1T4ItaudIimmE8QKX04fxyiRKsIiKZKK7FBwR5a
ZDc4JJXCfI0biyQ+RmyNw3CPQi2CuwOMsdREE95IkUNxJAGbApkGN0rPLWMWJuvuCY1Rr/tKnx5e
1yBH6IlzVTCa7e5YFJsrjtutWWHYr5eBb8InMYsK+yoFTXpYexRmeA4n1eY0Kqmt0L/wXmI3toGi
jV0KgHB8APLyDflxw1zFggQBYKclcA1v2oza1jEUFWf5cOQxpknOg64cmoxrmDY7fU+N8esEMeJu
GVyqPSy3L3limD/ztl3Oj6qyDfPGFYYvhPb7YYmT9fMrm12vTF7l73nsovE18/yyynbMOpLCmSnp
2aEeOcUm5VG1GA/yeGL6l+zvL8GJpiKcX1FF1lRAmJdP3IkwDlzPYGHRA2LrvryiI9/ETlUxBtl2
XhskP/6D+6CIsVGmDZOlW8AGDsudiEox02cbFCRDHmvSX5084at2cBfV7canLj6Gp6PScsxLlA/k
+7//hZ7JmliIygtfMGc/LZ9hLJJmdFWfh1q+5Fmfrc6SX962B2g2EhQCEmLw17EScefDBkwHX1gQ
L95xYBA5uYqm0Q71hp1P0t3Ai13Q39fUY9RaV3YHiFw5AgTYFQiISO328Ao7wJpEcv9q2oYHGydd
FMwiMopNb0LLGLf1Q6gtcf+xJ2TkAKY3Z973TFvMGaDCP1bUvM10z/gjzYAf+PavMuefrP5ryY5D
FWxraX1jgzjWORkMQXkJJiXRZPtfweo0zBkwkNfJT+Mlf0CoB2aEoJShTIa3iHee7XohsiYza+57
f6OwdEEC6kFqm/N/NlEfeiSOo2Qvjz0iIeiN+BPUAtL9owvZDCoDMdCKTz/UqGrONesk9S2BNva0
9NATCT1szaPHyaUqfk08drbjtP1Dafd4DC2FRK84mEiKtQEYFO+jvACUtgA2Hxd/xsyYDsedgVx6
a28zet1AjrV4dG3lr30P/C4dlznzWVMUGJyvXzyx8REeJVCkeuXddvrfJVaMT5X6sSGD/mGEgeB7
ySqPkMDG9j/JKsbU+0rRkiwJ+GwA43QsDf2xIn4TFZqY3KE7H+To4aWkHB9iIEOplqjansc4l1U2
w3Ld3B6wYlPTW51owsvP1eaEcYudFRn8aUlwQ0A70nOtTnpwUcCx2tTNejCas3hxOQ9vtFQT9jND
T0ZBib264PwZS0UCRcCBVT6pkLQrj86JqVsl5bUX316FLtHultWUdwpP0dWVk01cztW7PzUDGX3E
E73ILPRmPRZejeUSEB3E/e3P7jLp1YtAqDX05OhVXPSvZtPFi+7hsSGVz8NTOZgt1kFFK5mV6CfJ
5IfDYFMjMu3OnAbn/vw9FnhURaOYJYxVaeDrXU+dJkPvl7DqwAyczx2CdfDIhyLee/J1BTzyfjYA
PFTiI2Yh73CV6TTt3QsMoJ4kxh+RFkyc3Xe+wyUDgwwyqdE+OMAVffCixS0+F2irYXTuS2/06E3M
Cr4G2lgMEfV1fXjHRFnCtKYybEw1bWlsJ+zMUkbE+MCV0Y1vIgqNj1gxM4ctJ9oFqbh9gn9Rn51W
fGnGHm5DOFFN843M1vSj8wj9+XJac7rv2b1bwVc77XqYbk+uKosoIm+f+Dqy5RVN7Fo5L7dk9MBQ
M1Mr1EeYUVFr4nGbfHaXCIoBI7ijsnwtyYqQTvFUQSliTxA1XFywpAoD1ad3u5zV/df95QbdQgGD
DfOgCqcdnit2Q8EBX0L2+VxSf+IE5tTXXoTapEtUE1EYtjUd6fvq99AXeDPKfWp1Yth8G0hqz4B4
MM0270d+I8S7PGTVa4Q8t4XhorULlbiD+KyU5C1ojbgpP/f30uwUjrrWN9FVcP80mnH2fbu5G5H4
jObCh3w1IgncOn95NWKdK+yo+jAIv3tpIYT5MymJOlRn5VyXjZ2A8BVpihO2La3/8Cx3ijG2HNUF
LajkN5WOc4FNwmyPuzbrQboNMR0UFRCPE0iQaMWkq5g0AJjd3CM4oVhvX/3+0wyxnUCxjNdDOyLX
M/A/tUMoVELpMd7J4Q69UPHO4Po4bEJq7+YxX9iFsgae27wS05W8PR8v20mS11kfNEolMPU15LUr
wGojXfjserK8aAwoaYw+bg5NmesTXwKQZCgOah+ex2erKlupju/t5/ARdI/MaB00c7xnjLfgvF5y
A7tBR43nje1o5B7XQNSLxEYqrP89bpGh7hioj0Y1CXVl6zv79UOjyJaEbp7xhJinU1x+eW2yektD
L+3Spp9A6is7VUH4XjYcMS0SLbnUEvlWOHEoPHsGJvVfFmxAq/F/YP50EDXf7yzo1miQl9buEa9E
BgScnQcTnRJbzdfPAG/UxE3X2qxpQLYDd6nD1LUR1gWsh7AXh/8d/cGo0yBCWriaNh4KZn/P1eyA
rX3p41fTzNGsFy0AvIXNJ3ceVHhTOVShRUhNg+TCnrrbL698I+0d5+elUAp0yoazP3deYO1OOJEq
JA1Pr8aKaE6Bbp+8jACuACFC/S1ApI0pKglifQe8MkKnNPUIg81p9ocgcyMXNHnw3SI7Y7LZp4wd
AQpTV94sp2ofB2j4CE6ipFMvD5hXmAnwLaE708JUjVTWl6SsSj1Be0pv0okzvqDGUKjcJ2nmBVwf
l3uDwwWCcSrI9cLHOcxIFNSO2pQXRCb0L5o1dgPH5+CdQpc0kRhFk/l8/qdOJ4Y4VfmTr6Wkb82l
P4cdmfkdB66ckf4VgTL/qrRZlsHL+CSofKkmcjdJGQbV5UWTU57LhYXe5NHGgxIPCWpBd160eh8S
3kgdlPuPSkyCiJxB4cgevS8UyCV8yx2HW5n26nYqOWM8b5iDasQ+2sMMPNec2BBHxQ7CaaXHToWI
9A7dgAaedv8NyPiF69rLSvMXnSzOyQg90GsWftZyqEDxAjLJKZA6gz7OhJJ2qj4x8WXKfbyQCCRl
hCqoThRPmntZxlEbqV4WYMfAYM1zg5Ql/CDWlIf0xc7/Ic9lPXRtmvrsXuknxeaZ74GNqG2ObJiT
sMyeRCW5Zea5KK+U42lnsK9vnvJVZA42Cd07OAPoR7do4EwJ92ZFIc/KrzO/puKi5WYvf40SufSZ
MiLivvThvgm9wzdOIOfGFuvtb7G3z8Uqifw4h/RgGDlBtdimfJMtzlTnsKxwokPW2W/FcIMinMkc
zuQ7anMcl1le5ZukYD75omWykWY9jASTqU1W3DqdubNf2k/LhM4xrzH7tMCxuuro/JrfK83XbKgs
xXPEFxhP1u3cj9ozm7oXcJbV1sqFYOT4yaQYMOvZ444/LybgoX7SL3a/EHyStibeHd8OiYF0I0dq
mz4vNi9RNiYmkKfGGQZTntFdUsltnx1vYVJ+5cY7qRxoYeSFQSa4StFzzEYJguewPUgZI4mOYh/8
Esh0JFv2xO78eAr8Pf+464S/RKEtreVbOmWTogqydKJ9s6kzKFfdCTxpCbULmlPPqLOeheS24rnx
JTwC51G8Qlk2xHjtW15mVTu7gtEETc/b/j+BjW8TCeDTDVrBoDZrzQdgULYOynPzPRtUbFBnM5LS
4wYiJZ6MhF5PEOuehPQX62/NzeHfTFUayphYYbfER4EFMy7Lcxf76XvxrvRpjGd4AOaUMYYgPP7B
ng0XNMDta+EB/hx5kz+Gh3/JJs7eu6q7wciIsqy2W4s1hlGg5o079xsT8DyIVuc98O7c4dQswUx+
fxFbD+EhPWlOCYrvkgAL88mVDnWq1kLlzGlFP8Fq6quu307nZckoXS/DgiczyVuNGfMvIBCff+HY
CnKMYRS00S1nwA6u7vsIqgd0GB5nlMAx+qt0H+dexigAeIhD95dNXEF8vwUpxJNeINc8SmUBboWs
qjw0l7h3rLp1s2SAEIj6IPCtvQmeIHUVIDHAlKc26Wv5Kgr4u8U9e7eU+BCTGkjoRSOzxZy69YHS
ygVk+LK2VFfzMRk6wwH2bdsmD8/NVdBW2cxosi5zx4lbxFxfhDIRyO39C82Wn6tP12Res/M/pEXW
daMSw9nVsRfzjtfz21oSj+6rykfkFBzuJ9WG17ORzEe0niGDvbnaVdZBp3PJxGaoHnz20ZjaHH27
svLKCLHTgXwXpnMO6Mvd7l5z5Q6SqfXpKuSPip3WGZfMEalLVAsFBYlULgurMXHABA7Tp8BnxzE4
7QzGEPrmvlwBBC1FoPpBkGLXs2qjU6hk5l+DDouGxeC0A8fOTfCmY4NsndCFhVrZLwgZ8sCcQShV
VyUHYaRzsaK9uWDBiAd5ThXL0lSW/uVHrF7d2PKTWHaI2+j761tc+WXWtbmLYQGQqa/U+2z6WVzS
yfI4GrlA6W5NNIPJtogwREzB0oaDsRW3t7+yvnZFGXaaGNxC9xlQayFnpFO1GFcsZsKcxlxrylYw
YJIuZGCYrSKINT4yeclEcSolhsPWWTD9GHW+mnsrR9ZvkS9mNePYg9NzR4/3L2DyLopqf1fUU6Xu
9gLdnx85RvjigCYNrpg8cSGbgYZT65Ch0KKlaf+LYVQbblYPskPHlM33rxVbvIy7banXiAk3w++u
pj4V25vbZ7zsqdEGpeIKYw3FK5bhuf642krJmCDQFV8axVHOGXBelPhdAzlovuNBG/EXleMHrSbU
447yx1ZFC6EBg/BkejF5//36wTRDZcste+AiOROp7YHK89UaJpkpKPZEdBGZEtQNRCFtMTPx19pB
+PrQYzg76rQDAs/VO5Ij2RvtYKU2tq+k68lc3hA4xOrdnfVzNNZaL0kla4BhERt4FHjSpJmpqQA5
8OChsopSp5MRFOvN9QVi6tRjY5o4px6x5hHbLNgURczjzjw9s3fuW32FGsQVCT24Ue+LY3qKgf56
mevoyj+qMudjw5UOLWIiG4qnelb3Z0sWbrspNTSapH7s0R1d0PwhVn0l7bMsxbek2dBLiGjfIUn2
BLC8GK1XjGHFgWH6lqksE0HEmlASiXcQKiPioNf5QkONwkPZdS+nBgS93wtllbYZKj580idrCETF
7GBG2M8ihF0JhG+sJBYIwMUxQx3+wG1If+Xmz5TRcZarIZLFg1o+WHTnEYrDOhDorIESfSE6/wop
wWweDoFGJlxrBSHG+5yXow60deZHmyrd4URGrPkxNYMRkl+pTDem/6xaJ4VEIqhpF2KGYsvsB/Vb
Qrj6vQ9iIEAuCjTRNXF5Upb74G8ZiEWwQzttvJxuZy2jQvPQvsgDNZ1jujTch5Hh+iGXFjbhmZnm
dG2oXDArww/6iLCJHA80/cIDv91OXlrWqajeaPG54NJoUbnznSyjjPbYZZsdagXlS0YbpQZTSmm3
nkJZEnpKN9xJxPTliz4e2B6unHWq41OC9Lqmjec5OdhPiqylmsYsyDltqlQ35b8US59s4MWznBvg
nJMa+WBDnFo5I3r+/3X7oSce4uFK3fSW7ip7SNISI3vcoHNvgejwiYj7NNIsQH3499TxCgzBG8UK
KYDWCRotlZe5m/JRx/a1uxlFoYejZSn5Ncw/5iia12iTo/YxTiehvBMW3qdEuqLYGTGwfrPKp7ge
orJqpT0LkIAx+HmPD3+PDZpW9CryZhZBkXVoEeEM1hdte8Jr9CnWkeuRuAezwky2PXOg57/y4fbK
ErLvNS8D/cR6fhyrnXao/KtYS/UE8MYyMydp8JnXQwXx+FNHhW1lEO7FqMWq/AtuhdfuY6J26gGk
utyGO0KtIVoIYQc/xZ30NMe21qUfpdPqDCoCsF1lDF0ejo2p8yaiJ4N3VlgbIVXPgUyjDnEiRF28
KhFYuOUjZEgQqIKrMJIVEBIux7p33XkofuHs2ENYTE29hGte/tRT+UP8QSQe0vpClJZ2fEvfBqBQ
aV/0Gz3K+WEfSWa+Yk+2iaW1yjbH6nyWlyJdSBgkxWo+DbW0kRa5ENm4+WdvLjvA4sSGXMYEu2qx
X7uXopHIlzUPaHouTOcYJbLWGuJ3QwWsz0w6V3Tboq2rq65mXSbpjIKT3eRCJguVjiOZjQntLO63
zinnnC7tJ4I8UKRyUmbjNAbzuGBPcpntWGKIXpPxokO2cJH+48cV6TwVr4IQgi87PkkPFupFSWaO
31HbzzWQsuiCN+O/HQ1XkDaZUCreEncfAlMr0uUYhPtwQ2ZrHKXsm9Pkegw6QERmp+kCuPk6I7Ou
ycm+dr67A7I0++XOz8CKjt7xADcdLuNAybVwRzjY3PFoqvTLJrDyPYdkDvlkIb4i9UZSrYj1Iiel
QnYChdPrBa0V068dwEqR6muXX9CE3bxhzUpYBvSuW/lJNZD/aDOrg4Hsj/2Vg5xNcCzcFIwavXzl
zPKvORtEiBrXNL541mHSEyd0Cza7dx2B/xxxhIgzjPWJZZLcUE4wosfOpC+h772c5LgNl/cW/1v4
Kzjg3vekV/B3nKsP6NqIU8zBuOSyouREWhsvtgjlkjaunmJ3i8nH3fS7vwK9TN+/TEo8ZDrGdBft
084GbrI7NQnNNRs9mdObauCmPmjsba+LgNpYBJI9WbjPcNiF00FNMVG+eEjy9AHHjlCcBLdrc0+c
fTx5S6b9sYfxzdR9hkTe1wg/55ARileNGg5klvZh5c0lLzhcEfbKaeYmEBdLOoYMWPXpR3C30gIE
X2nFWqMIMLkvDmfqgkAPpc852tF6SY4p9c0b4GNUz+8EE7JLjr+LUpWOqIPMO4Vx+ZWCuf/i8qRH
KTrcPdTVpqp5M1K3LhFIqdiZ/Gt9Y2diKQ2b7X2C4wMnWXXOoXWXTMiY8HAZ2hc8c23zItD+yJxB
qkyciLYnpVE/x49JiA/LDeNOsCdvOY1rck5fi4zvjpHnDX8j1bNvHXtnH0gQXiEsup8TC93VRdV4
2P9QKDQl3zuYEy5J2xsEbR75T8q1wnTCN3s6eT64yZgup+r4jq2Cv6pRHfKiB4V+fl0ErHt+ebxf
5QkyglIINX9r2J+LXdRskjQ1lkLXGYZlPk4v+dmHTELcIHM4YngMfg0sOdXrqJvL3K9zSff3inzk
CMCuNr1V6CNZBU9p3saQK4EbKYU0DkAsh66DVCqkBwMfymkX5R6DZeO3KoYyljALhX8OBa2A16ha
bkQSDUv8GRASdUqvqm61mKR3JxSJTEjsok9ehhTVe7B07xJqJ5WZSBRQjLa+GzU3ZdRlexP10y+t
dswaxNY1oaTZITu5D4o/8L3+lNOmRkdWTL8HkGUB0nwx0m7lxKZFLIe/+PstImAyMPlNtYpvlJfY
hZ7OPJUPcB3R/wZFLdgxMgtgGRqVA3ATYYApIJnzgqQc+n2eFq+IGXNIcZs0ah5ZqUghVFijX/PY
x0ypZVu2u/66nkuKDSsZ/5LD6lMbWyxFvQ9TBk5B8TGpNPVUu3PY6teftkMgM/4xN9/m7CdWGGE4
AwyYyIyONNTac7peKngDskt2Zc/B6qJdCpsufT0MwML1IEc2q2dd9tpq9Eg4+qzOJrCt+vyHQR/+
wbJ7TT3NzN56uW0896FaooZr2XTl14iqbru+xeAyisnA9yzaoRn/kLnr0sHY5Ma3ZjtEvZL2LDha
Wld++JIJDp8Ju6uHx6NYoCAlytuWvXuj8c5mZpUq4ngvITagQ4tb85jFTUteQ9rNwvDFKIGxxjuo
4WwEYmdVnAFdUEXXX/Oq/L8FJxPtZNgKUD0W3b1xhF794eUmtSbe1P+EvQ/HFScQGJu26ZslzsYU
naRwD74rYP6ACDIgLzzwqZv0N1aOyYenpTETD8jEvIQmiOTbwCQ6Zdl0DNi6Wmn0Cv6wlZLEKj+Z
Jd2TRSO7csGPhXi7VuqFLBZsmEi2mzhS/9ysr3Rtlb4g6ken63ao2eeYD2frgMFA7KuxeiiEPf1i
YjTDoq7m9jv2xdQmF7KA6hyL5NKzii4ki1WW2UyoebX3Z7XNkRGRWTyj+Nk7YO5GFOjWcLwzDbv/
dNOAoEv7D4icezqXOfR13oLia0tbKQisX3nrCoAgKqw1/WtujzagLY/jejiwlT5re/A7BSSZwx+K
71telr5z9ESVw/V6EwRGqwkYcpAiKCHrmiu3C4DWfj2Q9pQ2z55g9X+NRbGEF0DPrFfKCzPEgK/k
ThWudPhGvNCdL8PA7XlOrwTkNOKs55pZp47Sjat928n5O/1xb+u0nzg5PBYHdkk1+7FpvmaaFZoo
VxXlP36caI1sCHmhnsayQR7sSEROiQ8ovDFHoFCGcBCJ9WZY3+lS87u8+zTgburjfkd1SsEtEVkB
nnY2lQ5rHmPCLTlunXSEK9WGA+kLVKXrhlQ7CQbKAQMd2MDEPjEerAhrhICS7g94L9w66c9S+TB4
qP2ShH7aGlq21Ju5HEksdupSXQ5CIhq0RL/ghp96Wjr9Yx1jX6odvELuy6/Nny3PI/fPs9zPRZVP
z9oT4ZTittX6SPKAoIeq6TXWCXBqHB6qJsK+W2gM+XdFNW9YEMRMlDwSwk+PYC0Ot/klp7OeFzr7
siGkv9+HOeiXEFo12m/JgX/Ya1sQelZNx8s6HoaE8stFa77TMJC0Tc3kAT/gwocs7iUAmgiJ0JhV
6XpIrvtzlqv1T+OV+tkp7Fuz2/K5j7D6/os15ns5xpLrpG/sQZBM2l7aDvgizesf8Kgq2P4FUoK9
5yb0Kq70bUQ410AQa8MvzL5mPRAxM0tivtWaPLkFSLjUnP7VO/Eaf2NMXnDMgPJNCXmexm/V/Lob
HOsb8H8BBJpKcvT+HZNtSAwBq2NanAeHqWUmAjWyOZw2sqC3B3HOoYtoCZ4G7qHG2jqRykUnf3Y7
2pFui7zqa0Pm+Qd/+wPfD59TVRgzk5A+lWVXZbFIQJ/HORHBYPShN4Lhbu/DguFm9OCjOOttlEgi
ejSznlWLM3H9ACbKldOD8nUxPMrOrgPaSq3wc/kmwwyaFHQzkL0dRNwyspU7Vo8DVzRo/RiNye+3
Ae7Bx9v4Msv/Xgw8kGWPxaCT+fc7PhMuOr30C5B9U8EFGEEI1ph2TQfIOClJY7yMEEFOuAFLNTbl
WklzDge389A31hXnDOfx3peIPrQkeuNVL6tJrHbl4OX6MoRwq2Liulx1+R3bSG5s7z+MfQVoCZkq
UxwGPZYBo51zdsAMvnwUU/YvmgKOy3rf8IBp7i5T4aAauTbVyDS14xe7uXmr5y3hPG1vjydvBwpt
fG+k7Wg9kXikhlMmwhAfu+nFCA0J/vQDzqKnKu7Jb2wPQRm7cyPbhP1tnnAjKb8nCIpnzdqntNuw
J0VIJSo88Hm14jfj2KNsvB4TSRqmENa9/StXBuUrdNbraezAIyNRPeLHfBV1QN/sUHe/2GxOEivp
k6ujtvjtLdXiH0rd0iLWp6MU9jvxvabtmBAv4Zm3ebfJpvdom2MA1UxpNaNTw3YH6/JL2ozSJqqq
oiFG9/M74WXstDqiKO6Q1mYo/mWZKb8c7KhCja1XfksvCZ5sIyl50gQVgfQkcR56clxyWd/C8WhJ
E9RARZ8JW1qCaOrgr+4L8cGjzkRmnSENP6wEr2yTpNxdiJ8BlQ0rpnXIH1oU8oQD+GGozOmetOtJ
XPfPoYQeRLTkmRcSs55XZGn2nnjOSN3fnZJGjIvwSLarAiXKV5i4gVPxB6zTRT48rSASlfKdcL6K
EyM7Cr/AgRHWCK+pOgQvPM1GDIBnsM7BiLAEWqrNbHAKQ5/9LmzoL/UB4ZKiHCyaAsfmAfsuiRVy
FCMRj8VqNKGzKcn3ulzmW8ipztprjc4zvsF09DvlC1A8LKLfXDKRuf1hC0aRMhLGZid/6VkDrCjC
fIDBoYmoDLZc2cHCKEiqUCpOaO5dyJjvBmehLPJFuobD8skDRMLetR+bKcwpWqwmI6zSlROi3yxh
lrCTcgY+exrTxnOTLbh2tu9ndvt5jnNnl5tUJM3VcCZYXdX/dgTJGUrvaUgma/zjQ2uSVswt4QwC
cmBExv3R3xD+XGdnkVnQ3CFNpZeLR48AR0pkyXzK4Pa/6NtwlZ+0Pparyon0Mtq7wm5Ye+WOZ9kZ
wDEbJKSiX88o5GLy4PROmrmixPYUDnB4KjkZegBUYPrWrrXFW6/o81hgsiO1cW5b4IKdLnfbiVSH
HCFlR2M5Dun6r339sa509J3nL8eE+I2Bl/VCiU1rtnVg9MTctUNZbJJ58tzZAG85Etmzaz0GBEHu
pfdUAT+Uq+e3m6+Zddp5aXoyoQ5odDZl+cpmB+uH7eOsz3teG9H88BJFH27BCv/IAzun8rYDR6ti
FvN3PgWYq8kX0rW5pu2GNljhzjPeqz60zuchmF4znOgAN/n0aOKoiIgVXedBDPt78O7nXaGcRzcX
X9i5whMvQX08fKSp/WaSiKizAuf9A0S7yJf3oY65KRT3plctDmJWJVuI6wqqovtWG6BWLMshAwAK
xZTIuBH/lIntYLPBgJK/AVfzBPqYv+RKTwN8wKcQ5NiQomnc0foU0NdPms4vNr6sh+Pf8jxKTSV2
cX7b9Y0TmQuhUCIHuCrOXFTX/I3T/gRUA4VNWeilfXpszdjKeq0hM7+7fyluc1Pw4ywqnEWvt2W/
oiGOAxHS78QcdJsmQi/i/OiQOr8xDWvTElKNNvMnBfVJt04ZkWavaPWxnuGfAHw3kT1fo07+PTbO
JSio1vLQI1KTyu7MKpBFs8c8ddODPPxQboMVKCytDIZd8gG9gjWuMrUNUGZwUAdJPUAKt9fH7xpS
Ziwv71ab4S8JzKJWyh3DqjEEdvW+mJBiTD3sEoGwBZOlDscfQqY+fXvIf+qVgS/8mzwMo0T1XWVx
IDXIYZuYkWWWN3n3odn51U+CKcQzu4anEQnZdZ7587kQCByzqsg4zySjZAU9DBvkKJ3+UUfgNqvq
/Z94uc7nNk6tIz7+JBBrtSNkbfnuXQU96BhDBBknNmATXWWWnFiTQZTWMony/L5JfB5mRy26UmZ9
4Q7YN1yOxVmj1rL98vHU4mM1QeTO+zxcCDayp2rqmI/P1sAd4c+e7vDGbhE85HWogEhPFDkUg6az
kAv8zORskAKcQT01UkYIRKSW1HnCWAYYaMBE1Dgx5nrINg822tQX1YAwXrDul3MdmFF55shvl9UK
G1rL+nlBrnY0Wm+ZcVZd6ulBo813vwClnZxLRZDCVIXTZoBCJsvIsQVlSFcjUcyz2V/JqEOQArnU
0KwZNnXPLDah7JGiTANVKMtlMDF9u0XA971+jLMFzn4Ygv+Pa86bnKEwTQnJQSaEPTQ3/LV90kGa
FILUqi942+afTEXFsP/1HdmC2n4N/TU+1z9IBDw1dfupozQBrKxLqUkBD1XtdU6+gVYt/IM8PzrC
L6JeJz2WTAY2Z0JDRtDSupCp55SaVyCYNO4MrQxqn9B7zSLFNMIqvSrQpRUaYOE3PJ+vz8Zkjbp+
hCTuyqdBrLKs76fBDYdfpcEZ1xDqw0rJZGidOMLnkOaEN0c4oeVgkeLvYDTyR3gRa4WQgk8JkZc9
Yh/MN+DQzLO0RhBu70GXQ09xgfGuktoEZlOZcUXAXD5qNQrCqbsISiBllZdmvEXVIzA7cyZqHyQX
DLNLlQxMzA/BNIlsL0WR7Gmd7+Q1piKRsQ4V1qexT1yUZe7Y3OPYhONNFEx/edElFGqcWlnv6xb6
fFePl6s8IN+EEOZl24lx/rtrclHmMbnAJGphdane5xDSK5bTgts4sXA+cr0IKcyh17RWHyMUHXJH
icrFd98LhOZTLK7Ie6+6BRtwdBprXrrMlg34799ALYvWUiC2dpDOSp7FEoRREPqD6xdRcURvRT4J
CBR2thkcxwC0xX3zQDlOz1GLvtC5utGxaOZ2j993S248Rm8Ki2z/Ya2amuFYgLaDOZEqWfTaN5u6
xztJiIKSZByRyBSV+YjzV0CE1di8TvQiigbSfcVauL35YnjDnnYzlWIrATG/CiCcZ7ISU0FpnAe5
IlLK0pv4tWi6SqEu4pVJiyZDiDb5obzR9E2RpikISylI1vEzeyOHv3Bt18/azCbNkXxBqrEBvgZR
GTfgDoE2h9CcVvc2Aa5VLNmpvnsRImlTh61+qA1bs1RwcgLbvX5oxvBlg2hb6vsPwslepe7yuXxQ
IqyPb0eJPkTGSSa3sBTUQLwZXz+o7sRdDZ5W4Op+zIc+TO73lUb/O+xOg22RsomIHvawcxmFdPP7
MxY5BcAlkb5wQrp5iCviAy1KIrddVZVJN7jwT7qSS7fYlbdg9sBahNkWfcg9UM3JxLxt/mQoo/bs
Tfq3rYyaTdLtQD+B8hrCORPElrZflKKmVx+B4AbalWaXQy+F9ZZTKPtoEKSRUYIHB/HJgiNs5yEP
w3iwmTwMicUa+Cm9nVrtm0i6xnQSGNqXI4buUerh1GTDiIAoVWOEq+27QZyucmS7QVeNWJM6j2WE
MTNwrcc5eZkJpZlXweRzVShYVERJPBCKNNf6htM/xyVZAON1SKKxyZiLpEh1NOtfhztCjhD1jeHI
q9qOM9arFo6cRmvvMJbeRfxAwLBoN8ZrkRlNjCtimcPltiImaFEK4kiII7NN1hHwejGHnCOwG6qD
9/aunFhVa9d3z23X1HdCct15w3ka3numpOFmaMa4YKaMKjdCtBwgUEdj3zx0js8doJoftl+dtU/l
p4QvjFkc579aCgMeoQwj5xSyb23+N++FSrf0bhg3NYAdCYr7nPPLpy2/pVnGB5cLns1bvJ4ijz8V
nrVDJefLGwlKgk1O6PX6X5TUnmePjCS3MferPx2QmqPo6cCZCXy7IUwnnPJM/gQEnjNATvFqsbn5
U15CFmZr38GDfsMj1WpL4LOqKe+jcDov10rRNfD+RVS5HPpIOfGMapldaPNz3rt0l3W21LpU14FB
p9ovOmdzJLCGrUorLbXYc+zWASWw9fU5bLeXBuS2QGdMAKDLjpzR5FvDO3w6yY3DmjY8WQeiUm/D
agWl2115l+nR4WWh72pxi2g16fzVzp39ba/MZqOJT3TFx0qPdNfhcj7IGR1u9L7E+oGFo6dBZ+5m
gk2ILwGT3rEBHJksBWlVq8z8M5DpOTOn9528LyAI1ZcYot9QGQK8ibjeCtuhHObFRgwEWfQENQr4
G8QBr5vVOmCg2/eOLAJYB3LkmT5x4Yp6kgapJexitOSU1lbGvxFsQqFLvv0ql+iTxnmmG/M5StSX
MvRJCXFvMDl8k+YH1xUBnjVzYN54jCN5gCZcFGWkLeRPMmuuT0kWqkqW113Vw3BjPmtNo7PTMaXA
e6iJF2uQGccFCCof7bDzr62rHrHNeSMW8iz1P5/t50iZuROt0Jz+b6EFgO93qKAMUsFWoPulirGe
fhvLXMjwQgZg4uKjXM/0rIndgs2Fql4kL376Z6GrE9zxgtl1YqIV8EiTmktGl9MuTKd24vxX9U4T
TjQ3uIeJS3yDe4C7zQYF3w+iRd6gefEflb5RxUCi9UIz0jjl1qt1PzcAgwF6aksc8LvOgqHNPgaa
OhelBXexcecw7L2zfTUJwRDjk7N3yWnJIZQRqB7k6COr/tVavUea7Ev3M1R8hRjq58MWkf5ZcHCT
xy8N89izImPRomheWiz1U1brju8T3qiQ12vEfpfxTSOj4UiYNomUngwZmjm+7ra/Jc7ktxE9vr2L
3lnP0sjyBvn2beWxKlHqr7Yhf+yJz8okWgtb14ZCXKaWsDZbjSEcWBA8F5kbZTw+9I14ES3b4stE
eQThgmGm0obNXqqtFTYFzfXd2xyCN1IVZG2njQGT1QPCQ7zyzLjpA+eScNKkmVnpvNNPaNNYnKGm
yxw8k9sPcY1Er69kYmxC3omGbfobJ0fwA77h1LtvSZGXv26FFV73kJAI0p1mizuw7iLmoaqewH91
0JxJoeKCqsg2Bt94JSjE5ZvIhbdbmb5OuVVhtEYTwruq80LNpO062zDaAHsLYutUapFzOrr8Xk7J
jpMRX+fOJ//Fc6jnV0nu/1q/WB4lEIE5EwxRhDlO0XfBCaofPUEfFDHxZ4jYPNzj8/L4OVK7CWSP
ZIcPVz7ovHxT7zNhpMEAtOLdgEvnikVkqFgqxbJBD4+7Otjd+VKdoB6qCrCP13Y0+osyHQxNLPKv
geAQiOU1OYMILFekitpLTz3cw2cVMfGhjpG1rkqLATvJqfZaH4HqFv7kHnaP6MN3ESzacHRX2moK
wW3az2Peze+U3OH6tat5RkMozAYyR7Ht5vqfxEcaITpy/T0Nh4v2jer4XFwuXTFbHIirrvwnK2qG
qvZoQMB+e+TIsfrfHhaI6UPu695X2m918GmSg/U5zKkH43iguij+6ywRmKRzxaZTFe/QqpKtSF3V
WW7AtcOp9HqL+l1Xtscs/MjCPHpWYzuags2folvjKRC7yJqinqdgXMDssBMX9w9GT/UYw8ka7Q27
2mqNzUFLzyp1c/RLyV+iQWhXHPhk7MOaVpcu+6aayq589xYGcHPOWnQi5VXOHp69Qfy5LkLQvE4W
k7x8YDnbruird8lBYe2nxK55Kfw7DARoziehrrnsr4qwPddnihvQl6aMPLxTSys/CNBLpRN/+Osa
t1vPAvRmdKlVlPLYzGQUdtGTz2/HOngAWuiJfd9LbFDWL07pvptXMyTdYBwFq13VVsOh+hwKzPG6
vpvIRMSrBlAkKMc8EZa0w/bcnv5HFJQzXwUwoixYOyI5m3oM/qDotuc1+Acur2G/uPEQurzGHU5o
jjLHxTsh/8TdhFF0Up7Xo3QkUKz9XSnCO8W65REhIeWh5Seh9n/38VHLKo6VAaj8FFJ2V4eQFb2S
4cKGKW1MTKiXx9Jemkve/1Bzr1zBekxjQQcafL07j+FHa9s5rG91es3mwheejdpGEN86aHjrFPZY
ZkRlyNcjaIPlcZ1Yvq3CT3y/xseYDcygBX0wWIoFqr1J/WSnTw8aPw1NdM8B6m0+bE9SEa8Tr7Mi
85PiwRjSjW7e8n+m5eYNqgjOrWL+wKsFPqyA7/Nq2ovroqXw2E+hC9gzEsiD/BUGLWJ4sQDILulM
Curv2IcVkcQHiXGipnTJAIAWYoFuubO0c+dyAjSH+ZLt5TwZXmavFWq00iv6YTXQv9rlTEf7Y0d6
QVYHGKPlAvRI9WGuiMQ9mn++mQA/pFeKDrNNza6FePwCTPZrzJg/DJyL2Af7ASj/xCc7lxb7yzfR
pucqXbaquzt7eik1ezDgqBaeYyZJJT07xD6Fgc3uLVtCYlq0fcT4/8a32uWpEnEE5MLKKmd2t5K/
+fcnDrp6V6qkV/ODnKOF6Tpt+JhC5/g/jJKq8KkhLkzjN29c8Cv+fN+ieQmKqNAhjXW9CYCtuqPF
cWAx890R55Dk8pVgo1dLV47R4REpxUB4cvFgPL7lzUXscIAarx6OWz+GWxmAJynO6GBuHsoFxDhv
Uq/cie7W+3jsoUBriaJVsKnoJ7cLCANFYBsNiqzdEzF4TYlmWzlx56rJ06M7aDcT0PVPBBAMTdAm
b2/0UtWYlyoeyaIUys3mqJ6HhuSIoSpPcEEDQ6lXI0dU4hYE1pUqHSmMJamZLJtRmLjDZ2Tdl31p
BQVN/O+Lu+/YUYmkl37MDEsCYOqs13RqxNbRFJ2HxDU2qcos9maL/ZsGqSTwd/6NU/F1NjTvNPyv
kbI1yldfTQdYeU7T1hIUDxL1Y/zjScRVQeqlnDnzRgefzzMcG26DPZLE6wTDg8zOXuTQFHosBOY+
1Prm2POUY8DFHl5djY8Ls179oPBgUaCh735EdmvYmgBiNMJi08QWF2fgvRyUXo6O193WxaAuZeMt
QLmXhVefRl7siP0Bx6FAC3OuaatE8ZXDh16hpngkxiBkBi+KHK7FI5YNxwdAleGwHHQPAT3YKKPH
7ALjn4qi5REb3+TRPF7ptLNGh5sDoIjC4vsuZ75tUj2DHjObgj3+bxOOHpnRHrU62vwF0OkqCjNm
4N6hsGs0za5d+KQYY/3v+rBnxMIk3DV1T1YECFn83vJbhy80hrCXHKzMqU1SjHedVpWjBlsfok0X
3xeP9OwNcTRlkofmWkgGRTqb98JgoJzPlh5C3rugc7qM8CK1iQ9Y7GD2A60FLifhVd/ByqJ35qQl
pMT7QX47yE25xWFvdD2G5V9q9Hvttu92tP/tciBrkFe2h53MFPfIsxdewO6PQSj2bHm4Gs/d6Okr
FiMxFRaCVvxa0skeRa3pDbYTNJveA9vBzoXiFTqUoIM+OXemsYHQI02Cp9Shx5Ydi/n6q0QwNBWl
cRvYmonsNC6au5ixgIVlTvLhvjva0Nsk7q5bTElF2T0RXUmL9kbOEExIsSR/HVzR5DTx+YLS+wW+
ugqW1cGFt/eyGVK4bDMkh4R6YXSS944SHwQLPmTuH3bG2wvMTSI+1woMwhq1WdREP/mILWa3qSYM
FMNmp6Y92nl69FOKhJh8W6gNr6tvJI/pFxaVAfeip0y0YihZU1hYeO/aUEbs70y11ekYIzeP+9OM
WTgoR/Y5etKoasvqzhHdd7iZG2AcJ36viDAS99xR9gsxnpF2UXQY1ZRM5cKPMiVpM9y7spz2tv3M
UwIAwL86AgO9A5NBTLLbulFbMxPgIeQWLqDCoeBkCFRqPzra8aJ9SpW27hPQVPUfwv2HuzDPgcXC
ADWMGl4ViP9rdR1Uu2McW0PydE3mSTBG02ipIGcbJLXG2dR5Noc5mHtDNWt60GFrhL1Irwfj4aKe
aySN6FLWBuhPWTt2chZUhsdq9Qv1YW81DsCtqeoj0ad7AY9Jo954/HRtG3o94SwBDRv1X1SdT23B
axXLb5ZjyZoIDPuojPNFEosB9g30S6n1gsA032DgE4+KW+lVsrkvvSDBcASFgMh6HieS14l/Cpow
JNlbBIlnlu5msBNy59gHYg+WnYn2+64iYZxOIgBo+NjsOIKo9wtx6pzTNRjA/rZGgFsypDLNH2s1
X2xIlPKFDF3/c+Y8gazFinWTHjJUVKQ24hZRpvQC6c3TFpk0/oNyYxevI6W/MYBjanWp5BJpNO6a
bbXcVBt2AJfRUzN+cQ4+3iBFlQ5RcV0ILxv+BNDqGai8arYD9vScKd9LhOwcIDvXMCHY+gS0z1K9
RBowy0SP3mrdyeGoldnsuQIYOOFlQf//9RLen6l96vLwmsTZ2YRuiPEtfeRh2894a3yN5HDgHwTD
CQEngmslVFT/vyCJ7UcPpHkfGNeh20Il4fJKRSDBjIA89QIQu0B6L4zb1nlPyDz9GBx1OFDVT2VK
/cNZvyM9lUML4JiC+Jskywqn/RBeYRQB7VGAVkDV8rm7DCNwg3u2WlkzGz1ZXwNj/qRB4Z7nd9Cu
dRvnXTlEhcFaM+FZm2kH1H9xeAs25ewXqZWbaIRgLDI/YKYHl5voTY+tJU9/ycY+7YDRZJ5a9lCC
bKprCZ26Pkh92TbVIglMvUCoO+fEkWl4hG2IRth5bTKLmcpaEHfz6+Xj7CNJZJPyDaLI1XvvtpqV
Ovt0TOMhh2vcP1TBlvEPzlFCJHYUA0NmlbvICSF3OoQ4vMBBtwVrO1bGjEZl+lKgyY1sEkTspIs+
BrbvS5mUOQFV6sT8bu68fwkHJztvlmfipKcHf6cNN063217/BRms0YlyvhnVxbABV9g1tkueuvba
yq3LadDPCOml54ghi4c87xZW60crUNMVklEx5hODH3GkWWQyTXcVrpwVz0eJWxWRcw2CCNhaSmMm
uCduxBqGsaPhPzAkhAH/0jPJsOHinAswHyuxz5yPUxz1vmBnxE3LD8a9nV0M62pxdhOYluX2815k
K+aTQR9wO8IKoIhrR7MPLxaQ1qM6q3RZyQU8ff5C6nRPynGRV6EfX0veq82gqsPQ6ZABnrSU2QH3
yxyyMaGVUT3aSX2dK9eQSxHx1D/c1lM5/XtKvvv3cfs2b6/UaQywp4rbDGTuGiXQSGpanNr+PP8S
9WYoTpUFVWsSmU6UYMWixa4i3iDESEyV7wNgOYxAB8vnmiTiU+n7A05R8YZFC7xkDnnGsL+HDnX2
z7hqO3yPMXlkjYuDsigKf/XOcHRIfhjs2JdXxTaV4ozoa15vGdx02bn/KL/5qMWzHoN3yEqtXRsC
I63vpz8/UNgfsjqrBpQNGYgXf1r9qMXY6MPjnV8ZEqI0m4bu7KfLQZwr3OkZIm1mM6mrMwtxpMQA
gv2XcZT7G8JfqekqhEsKOEtRBQ9Dz75QnhqnICcxvnosqPH8/BHsUjTGm2bggQ48fPhkuuoWK39H
OcSWjTvdFaoLujCgEvFte+ZqgjDXqmjm4JyRvEcrJ0Ka/E6PyJ0CGH0fR52DXZ9wuXJoFoYvgkGt
YLLdWqCf1TcGbGIqGA2ngGvyN+72X4ZhusY0jNnW/Mn1L2CxqiWlm0lydih5L6BtSAk1TnSTqGqK
Mt3SNp/DFESTsRrbAiKbby7ojtS2UzlGib9LFWdk6Hz+pMxpLl9hX/w3fGVelbG/77s++dx3IDyy
TnSZ0NFLT4akypxYP4VtUQ+TlMfHCKC9rMYN5/eMMHL3i5fSn/6opH4X89UgefD/OKs7icVBGJ5z
80JFdvTSEOylYBcGgP2q3s1pG6x58uo2+qfMs44LTVkIDuCz2dPiyNVzDLPs5yb8HwenlRjOdXGm
Z7FgESKRwtL+UdWp1Qm/mubRS+f71TdpbKwn8FjFgtAJvtkqJJieoNAZY6IQPfJVbTgjyojS9o9V
3m0R9aUXAlpTt0ge2e6jAxbVWrV86pAV6rF0YsfWM4eshB9e/zmVfvCtTRhwhoxM1wzu3nOGpZ/F
elTgeGXGwLulRKy5Fo7Pr42zyFcSZRlpYW075RepOlVK/BOifqlwzVXiBmUoHPapON1X1eqCmQoP
iYamOAjX13/ll8LV7hv3AZJiYq++HUsDmz7h48HyAa+7l0U8D3MTlWeZuQzDVmIOJxXFQvI+BTtr
OPCKz2xUB3LQgNhNURasvZTVMyKbdyft51mKUcLxpTe3C2KavikxOS88ubHq+nQj/8dlo8CR01U2
Ytc8fhBZ+iI5AQyemlyi8uAzcxSjjXNGCirI9uPUNqM0CIJcg/EsFFL60eSK7faYpAAsYXfd17zg
vdTUCxunt5S9oiWjf73qjGAVriyIiD4j0oOw0t4KvhMKy4MLfeGtaefOkbaQiEI9zFxWwDZI87W7
q5RdQTZw489KDc0hzrFwhVYAfhaOfx1aKZAZ58JvUUsb1dxW95pauRTeQShXrODMj9SWp2E33BLE
C7AVGASnhNXDQBu2zpqzKow6FedDLIRUdkE9QZ2r6/O2picLCF6V5O1qNIOfzobdTY/KlqzDYkRY
496VPSFbxtAgRjdaxgNRAdk5zF0JRme+5BAKYuQsLhyJQ7DlcOMEBG9WfZVraOpwFHd4UNB7J0TL
ORMB6HZAHPCllkKdLxA61WDlXRkhPyrxD0gov8kT7JW3/gzolA5+Rlaxcza9g9wMKUKLALol5Mfu
96DyBYIDoGfKMzXIbicJTIslndhs8CKifMbWszbFGR/9eNJFwGme2qfWYgd6JfzZTOAoj/bfgWxg
CulWCFoQ0JGdInSRMNnk7QDgWAShI69zISMA+PlHhRgQO04PBnBMqvyibW4hnCMLdpoQfGB6rTi8
5zvmkXwvWMKtwQ689ZlrUNf1T7sH/BztUSxjXZYTTK+qRQBugEAusB01paRJsW9fmey3A5KAiSuz
Uoao/QxRbtGbdzS0Mkv79ugOPHnZTMjZGTffrl53tKjVhEcttd841rGjEGM2rrryPVq+4TUpfHEK
2VtI5AQWWXs0BRrP0AegtLJVEAGwfPb7wQjYWwongPTM4AZd+sEs4FPcxeni9CHCPZwoJaGjqiZA
Ic95aJhueklVGJkGOaKPHAYlSGyaeHF546c0bE55gZITYD2+HInYKQew3UASj+hcodKaOQUCirN9
D/Y+NNHAWlsHwcpWAtvvI2Uhk4EWrIRo9GBk37yO8sSutR8kacIRZhJ9OMIjfRL7g87+ZUVIg2Rg
/aAo3lKkcR/t/xlBdrJEmq86c+V47sgaNOVgpQwkt8Cy9iLlLx2ty4crvMj/u6fLBYkKMUs4A+A9
fpkIE6Ogg2ZdLjOYsRbJ6ocaT/Z1uPgKM8W64DwIkA9XLvfAAIQqw7Tgg/qbL68h1Xp+bYygdXhh
TegvudTu+YqxNAwI0xGvttGr0M8REqZKCkwC17yIKM8SObfjnnZNo6EH1a3MNtIgQTIxlNEEAydp
a3aJat3nP08Bje8bW9QxMCTIgkVr01J+mt9Be+fdxUFqe1rlNz4GMKdJpXzQaeGs57B1il+/fKb6
zZfKco7CdoJhWeB7W4N4hL+iIbEpHmspv8RkfFwXx4+y+NkxbckF+xVZ8teIdr5KiJFOXaBHB1vu
HoUFI9punCYZCFaoJ/axxF435kqBihX1KYOG8SlizJ6oTaubhG6ddLDUaUdtk+nQ8FkMbdKnvGy1
s16ROjAoZFKTIQLbILTzqSbPlnYHrsgb77bDZktXlZ4Nbfq0Q/xMcPwBRpF1wzsjBl6qsDgW02oU
EMBGakoG0/t+CSrvXLleEkKX+1F/GCzhgXJXFGnk9sAsn5p9ULaUwDdmoed/VtMgwCZdITd3ZnP4
VvldAWmR5H/yMBGJu2LfXEjZamu5pkmDQ/PFN7nBBd4gUxUEc1wpdfgrlJjAgw+W/PmPIr27xbIc
rWBZwbAElS9rjfFnX/Zh4gk3UHZDHRxvN8BAxB0fxt2SS3neW8rNPGHI+XGo94yEC6XD/GnWNPj4
HrAbMeioV4KlMcW16dhx2uLu+jH03YV1bPC7+N1wExByCIp6Qy0tGyJ+Fx8bsyw2KqlxuGNYTbYK
RxskwMo2AchQGQ90nhjd2VEYBmQDnTnavcauMsMKVkeBt5dhNN7u0twMMr8qfZLbd+k5Wv2dkULi
+//+EHNbZ6euJHoG9YoWjynFBjsVDK0uAWdvIN42fOBfV/ghZv+32NJPPSZY3ALxVusvXQtCSI9k
9bnKdhFM2KYYTnEbYuHkbqoYEkFbimoyDLphr2rqmSD4c+vEFAwvY+ArMqdhKcvUM1E3rTIELNEm
8YzjwsQuD2lusGwG+ovoyt/1WZOcHZUdHeUi1kHenoBgd/pdkYvBbmTyvupCeJbhhqVz85KJIDf8
d3hs0ruCTI1dT2wSfh/WR5QAksPywR3SyQU1AeBWH1seN+e92CCoqL3iMmj52LPvthzd/tmLoFww
qz2q6Mfg9jJYA2+f21KmPWrl8kPB5rkKaD8mcPlp1QDf9Ab9NEAiDuNZQXqu7lNU2FeHOcR5mEJr
PTGBdngJZ7je7e0RgiP2as9uqlRttpndYw4VSMJ1Ttil1904KDd0L3kC+uDvnLruj3enN/hsFgCt
squtIGvkPhLdpjCr4bjpNuEQ8UL/les6o2xa7jPJAyiKTkeUgFhQYthnAheUx1a/HcJQ2JLsnYet
wXr6rRWARTLtYNkAtEYFfu/cVPpkdBiTEU+0uO1JozyyjqL6KH/cfDaluQVXa4XRUVrPK2EX9/pH
UH1C2Ww+qXbcxSbyCxwSmUX1lwul7SQ6DqxNL1WcItZAbPZJOJsOqIvkzMScLUb4aR1dxlrv6jZN
JwEzDZHqp8inbOrK8DXqlBk5CzH/LyW4s2j46KQn7fJGWXfe8m/VbuMGIhuxsJ0KAqFvFHH88IHW
tiIk035sfiNsUi7K6brSv6ownBxRSYbr+mtOQ3shT8JT82eNZ5XtOcfb6N8TLIPrsAJcqyo3vV64
i8EMY0dCgokZaU6U6qQF5cuqRvzhsJLiKCVD6pF8Kt7IizlMVsbmhz9uXARl54IW5JOMedLErDzB
FRjMLw+3d+fFdpPQ/sStzZdd6M4GeRCzC+ImPV0xmjx23qARc5NH9bMpaKWDk0lXibwmCfu5yjMV
RKQXS+nGxdHTMVkUcPKpkLGZcbB8R4tFcn1j87s5b6cCZSgIFsPl59aXLru/nfkHXa+xNFwJQwBi
V1Pl5NfoXJ5jiLWEZKTfNZ/6s8unG2k9Z1TFQbGHIUm1gcmN2KDRLvbkCLoqbgjN/YiQuuLDCSxC
jpzw+UBVAzj0S8T6o5Yc/03gqlVg01Pg7HY0gdQOvQnvJuWvc1ndsENN1WsN0anvgx6OfA0DYXi4
bDXP1OtL060LiglH1gWYDGMww0aKt4hMuHmMDx8mQuayJBDmCcnBHW3b/y2eimC4S48tSS4A9zmA
S6LFyAqG5V6TJqv98K40NAxMM0qSLnl/33rzMdrEHnMA4brOhw5tQDGNhqyHinkbJ+wcSnYn5U64
fPr1Dbvc5i6BwMpcM6+3LdLsgZPbFYCA2DOAEEyVI4m5oTI/T/f9i0a7UR0wxHl44KkfBzG2I7EG
yLaM/3OHUYAtiurOFUQdffcXnJQwv01j9fia0LAf0ojJG5zwXwzYMrUZwaZAdbYlcIvAUwfovure
HX5WevH/+OHJDfIb9djVGfBGaNA3jWiS9VkjKQjcEphyZ5MOSe7fNbEBI8GgxGhjHTPoiYsnvNSu
KKqkGEVSJ1GgkNgO45UxcANij/HE4tX8ammY/q0nmC8nz6qUd+juc7dGXsHjToNMqmSlue1NYxzH
CDmLMZ3EuW/gNObHGDMAzqI61mg4DuzZ7NiALCPYPo5GghFUSMEMOjaGscZnVzal9RkxwdWx6B3S
FmfgeWwR2zGR5jsy08GWBLmkPoibeoEpMFotXceBPdw4NJ3Kyux735MmIdCnPIpu1sxbNyaW8QP5
dhthNEf3DjoEOlnDd7d1/GuJ2cv00R74xn4DLb+6hHUxJhlBIOv+3CUTLKobhSEissx+8li18lJP
IzsAP6I330Iz09u1dXKhmaBFX+6GjxrSV7XUo1vgDsO7wm2q766JQd5XT+6MYpwI1kBQ/rIlXrSh
RswLSzMPC1f3oX/eqd/bdT6zLA3LZz5naoM2PYon60jvvvIVZeO108u3DXjQYhTBkkofqPLM7Xbo
uovEMtYxSmm59MLJElqRB9sW3BJoBkln946jQRIjB87cvsgokTTddeJgDg5Fq5ieodVSCM44022v
vQPx1PIegLhDKdGCezKsKPdxEFswiYEHy9EIMPGsednzLQO1AJ8q4oCjHNIGcU6kglGSlPCDRtaN
3ydnNTvhGs/j2kwHPbb+axFVQAxtPHB+10ryoBCZYaoAMlg9Xc1nAjrtG7fKhmyDmlk/4yayu3tL
W/JIaoOec+p1oQiKjG//Go7LAuEkLVXsEDIDf8+UPbbL6Z9WmDGw+5glUwOkCMYwMKESx8Is7PkE
nlnDsuGyTKJ+8llfIKEVZzv5jIQb7IkQ8dgmOqund+ZQqokpH/wU7A1DUgAE7uoztzzd5WcR1pL2
pHWoKyo1JtVRL/6gELzYuxOVXvkx3B8IBGW5LTctBR9jXEXd0++bGnG5hdx1mnzB62PbZekrY2tz
AuT/AyQQUwEqkKEQgRlgS5JNoeQea2ZesEpgoj31oRw1RwgmDW9TGc7h5rbfRcK0bZwEZW7FVtrl
8BTuiRUqai855pNEzlrbZS3HvqBJCZa7cAavxWeq5FkE5xk6L/U5aLVTFW+RTa8rg060yoe1n/nG
01rqgC3qfYqv08EmMdpD6nOxI9esfAgqCldOSJ6Tz3aEHGFJl4aRG0HippC7zJ+31i2ArL3G1y7L
3JjmE9b2D4jM6CzeHt5nKZpDym6FcNrSnKs3meeNLUQpoN5xGPuDs4lYe+wXkI4RYBSUKaeRV+JG
YhLayhUHjZ5vmEE0mV1/42oCbIeElWNYTKilAVmupm9+NYCvdD96zVK2OfBb4NgLoemcaVUSrrt4
0ypUxqzQPdGyKUrW5VKAhS9L1M/P0hdHuvjx8ni3SyFm09AVs84+9vDxzL/DGjjc1y0l6jwJX18E
I0nR5kePySR2myvGmvqSF6pQSbKigPzg7+/4lz6Ow1eLbBIZFv5OHINRKLz9bX9eegdAsfAb3j1h
UPzH+sg9fwaOFYXbrt8cLZjLq05/nmT1gFMZxUyoexvcWiP5g1/lIWqkozKrtnBw/r8Odt8FwlYL
0t3CknIq/nzoqGNj2W2bfLHchqv6WvC3LrUqL8eF4d96PT+jHMSOeyTP6Y6FKLEZQy18cz8raPD+
WtKh7QmY4o4zwH5d1FMvjs3UjlS/sfr2EfqizHFDbLI8KEmz9x2ydqumJFLzu8Fj+e+pgNZbqG3K
a3h5l3IRfYVDNeq9LNn0yZhBwP18ZLYov109t4HIZOEfMKtXNPH8lVQG1WlZe1ZqciHk2FiVMNzm
OnwO7SMQx/sTccVpIdxKUIaLGXxkr7RVsb5IHt0RsiGsYIHaYZ/8O+fS26XCTNQNm9lBRYcwYIVt
TjjmTdn7oH73ngtOzFDLQEJLq1d/OwmREB4mrfHjl6rzhe8HnNtluL7Dc5+iBi/93NFtUDdzQE2o
d+6aUJNfKJrvRuBdBLcygBeUBHjnCDD0cmHEKXX4e8ef4dRRCkKJaQH7m2EOLNKHV2ggvCuLBm6A
wi/hJqfYIhFpTSEzL8GdVDQ/9N/JCfwVS+ugIAUlG4L035RrBxyZq+7EVCfkuAQTAw2dpbGyCur1
wBlwwOz9AVQqn/NKnBYrO9SKeJkZwlQjioaJHM+lFxt/A3dMRksp8wCln7nSFnruKbbct4ojN3Qv
y9iAR9Aahf6EMnEwkrAJ4fwvAotKoX3nzOH14QB2tAkfQk+jyzBqCPiyP7NOZ/Ha86qd7QPw9NUS
d/18OY9daR61UErXUolduhrhXOyKS8y9U+WTMUY+Kh+c5+MJzLQcX4fc2rR3lFTyrrTjXWHfxvQk
JzWGL5z42S97jQWWgAO4pLQWFfAEdlEQzSjPGmUUBbRDAK06UNmirVMcha/+74vRQfmXZwgfEBCZ
cJem0sE4jke/gdpcxaxA2I854eR3Ae7Ge+nrSC5Lfp8ezr1oLTnOdhq3OCmRMXGZRz9Lupj1GZv4
NT6yerLFg5IYnzJVK+bQvGnOnOnSnwr15p3Akzv9ExHNgo4UtG4+kvfmI2C2I/Qr82gEnWSLBb2I
5+rvRmnPwL3AHkynOKWlc2hN3YP59ZtJEaOx+ODY3HowXWs7BDJLkGS5pgzRVCzgPGV5EhcVwsZB
bcJ5Tf0Gjisn4ab1DLCJG9vv7T40YTsgGRJBWSIb9cBgv/ygMaURm93HvOBnqFL/WDD/eByq0nHW
OJK5xP6shUwNQWN+PMZk1TJP8OxTaFzVgGnhrXY2YmV/SB+xH6RbOSrc/mjzb+Zx8OpXzLPmqEEY
VjNiSX7v+PVCT1Lrgz60cnwcIK/t+er6/vzRz5XLhzSLjVkcsO/EZEIz05Yw/eBPKeCgCx3f2xr/
qHY3WzUtvfAsLXDFWjHuV6+qrOCD43dIRlwJkAriW0fTXim5+K2F7VNtq73hSasrgh4D68yZheX5
mx+7a8aVQc/gnoDnY7TU4ztyila2ybKeSOPf741nWWaD2O7vh+PP9FGT/LnZRAQpmaRnoNWkECFp
5N4eLmKW2raRuWB0hBsSjPu25SI/gQEOn/pPFYLeIcnvoOoBa7hB3TqUuu3kRYN7HlPE4tkFwFJ1
bBMM/o0jfLz7R19OdxR9m1eZJtEyroG1SEcHBB+oIB8xza99K3j9wD7gySNdpY27PdCtrzSBcfXs
tAewBIj6B08JKAMDnR6VfzefUXPepjTUgcwFD4W8u0vQ1k5vWlbi8lJQye8TJ40yBSQVdJS676uA
C86KTi1LKY/z4CiblN0eTqbwopqUJaVCpU5P9w3bAhdOdFa/fDAk/mt3g1NBcUdeOH0uo1WUaLDO
IsweDc53mgVHXGKBGd2tVpBnneK84ZcoP85DNeNnP8np+msuDpWqL9jlkw4ol5Z4XoQBGfj7Hdfw
eUNEtT98VLkWD9IsT4X4QS8yWAj0mkX+g2q0k1eqgLZs+1Z/EvbCYMcni3D/o4zvFTCNeDNeb6b2
PRri0+GRTutj+VJPQcwtToUI6cuzanVK3j+kEOPPASh6Sy8lY0D2y1TOVjMOlvGGen9Cv9NZgZKt
NCjKlJUddzx5HzYx/DRiHq/sxnuFdXQWQxghDXGDTSR7RlfUrkxUiUQnQ26K7Og5QcXfq+sawWF6
WsYPwyOAEY/7QWjKb8Ia17opoONatz4AXiUp3CmEdaAHVixw7l8Pv4ZCoEbYbPOkTd3eEVlrn/f7
NvXU6NEG2QuGZtGACKboCgCMXyeCqn8+aXniHcAiKwcbwno5lX2rQBXEmqzN9YidJK4uRxDWkyo5
PobyDYcMgGJOsQ6rxvOOR89RBDMtusud0BaXO/Io1epnHRkPhM9rMNxY+Fi/4VqI36okmDFvINmV
MMfcjVwF1TNI+kBz5BNizH6lD6xvJrhfTt4zafWnNvqicTOHcu5l0PxPWTObKQHxwthQj9umKy+c
abZaX1Zoa/uxeCTBgPgsN4j3XoadKrvI2pymiPZp0Wcr69CkK2v618eT1Xaf3OfIvx0OCnmmkphk
zcuetUr1z3torlvqCxWxrEJo0rzOexdZa/TJdbMdikRNkoA3HoZ2ZTHiQhRj3j54d7jRZhpYFlW7
PFi+iW9kUTyC9Ddsepdn2ygxGKaEthcPcAo5lALhdYzSAVfgPmyit1UXPcynv5CrHbINr2pkJljH
Nd/MaEnhf0gX5baUy2KZVPnt386JFvAivAXxOCP/eeTnq73cfB9+CWhuSrevgx572/6OwgDvu4/A
dixk7Ws6wNx8YRzLG/9u/wl2ieI2GB+7foYzzuHFdmlv+CSE9TPERkgFkIs0YizHhILFWDwkf1RW
JuQDhoqJ1Iqsupt1ATLnz6cjCczXtOgh/pyARvJtNlgvCQdBXfoaZRaYk0L3Bb4DLWC/4t8UfWzW
TngigurfwElisddLuueXJCjzG5OfMLFYmitsfDB0EM66mt1Fg/whhzVwY0XIGVJE3pq3cwlwIhY+
peqlP9YbsI0zdZvQGLTxbyJscF3CHdyJyh4mlyRUtjf3WWFlmlbpOFUlvIh9YAMC2pV+m4fg+ZOH
1k+7OtqwBtBnxstrEBD2mCar7zzpqPsF3NmfGwVUINlUbOnfpwa5NlNjEYhX9far3qO1C5afQZPr
tEJ+jpLiL1pT348oNz3GJoReSyp4ctyQ99/xdpaIpjazEE/wY6Eu5zrYf5HcGutd7TkCGQBCcf8o
T1/V0TPPBAu36cJg3LeQDMIgxUudzH3vOtXxvrYUEC+ubjN4HNB3/pBKftWJv/hN5CJ3qZDQynqL
KYMJlRAj1XrkMmF27kQRfqGDcRTlql2uiLhfZResj98cf5/VqQ3NuPbcmmVrOLfTdE4EI2ddQMA1
V3S9bTo542bob9SqzlLceMWvmID5C9DFWZe3G8IcHvkcI/5c5psOtnPRhItPIRgwYMhpxIGj+Nmg
KpYNij7gKn8WyOtywNnXB93iUZxYDPx8HlPmfqQGf/YnvMDpmtRENFRH2MPWrbyWKI6b+815Zl3W
xTYJqz9HYKWpEEdn10JFVebr53IJS57gP3qiS7S+31HtlofucGlRsvl/xUJ5wReVU+RDnve1Wumn
Bs+EwUF+wzfD1hB9YSnj3iIrDV0z1KQER9+HmkjxZsQAAt+AVkUfj9Ckn3MFWToFBWVpH+6SimW+
/391hh+VCVTPHj/qMckAtItvopNPy4buU0XUJZO8YXg+XXkw9e1YiySNtDHqqwjPmsC81SRBzSEE
BXjGR/hvQwAb/8poP5uh3Ln71gV8667Sp9Dv6LWyu+1+6EQuSZ3YhKVvpyTw6H4fQsT75o4/ud7u
Fe9TS6hXJuEoxd3QhHbstYIEJ0xU1QbHPK27VS2Jvfqma8qjuI7+Gwe60+B9jvZgnSjXBH8YIATJ
OBsRQi/gHQb5nDL1vHe4L5HpoLj2x1Hj53KtSQGg1mISn3AwoidhLAwjSQqkQPAdQF6gajqXGGsn
YvZI596MwvfFqU4+wKEKZy6Xp0wSU3cmxtrCuRyqtJKunI6gamk8OWXDWgeHA1dX7Bd/tOPtA6J8
14S5oVKiGdHtR6ISq1gch6xI5+4nlJfpUIc8BqZjW3ungilAa71duudpIVrwRkD0L22Ra4JJsRLn
b0BFcqzIhox4nX/teJt1T/9ifpSOBeVSxIZfHPHa+7PGxy+KVtiZQfr5AHqWFGJfqlCjueabft85
ETYLzoBzuXq8hL7RqQJ5SFLBLSwKa8xw2iNkhED7yVvY4UniGAMqUvCHRabgs7XH+4R8sH5hh8rv
M+70YXaSdzq8BancrNRWONQIxxpyUXX4lJiY1YcZwXrU1f3sDcKNybsV+3a4mXrgoIDOoi6FUU2v
vF2MLWsMQoBJiVFCJgG34MAQ/qyJkaJ9lERgoBgY5zpvcIOKXwhmMX6FJmDHBU9u5Upqdk8hI4nA
qEskXlOp8qOnYjKvnKyIWAPGkbP3CcEQJJoMSEaMfGEMKTJaxJIt7p3O2mjdK4i+aG8kCkgYJaTt
G6ndjx8LAvOERNrV4mwxn2edt4JSdUAaShCsR8sShp0BfER9BWbCY4ysv+oHlexySQ9NL9tBb2wF
r0rEjRvuRC9eE7l9sUDw/js/CBpM7yfThhV9nBqqe/9jgVR7aMIe7lGK7T8q4czUDkPkfhjh+Wxa
/ulzEh6J2Pm0ViSYyCYGDbfhxfdiP6d1dZe01hmY8JzGRkjfHK2DA88xD1MxjHpyHBbWQ4d1u2o3
l0uz5x50rh1u5bi3rLfBkX5cDhSbemnztIg3rjmyI7rBqH6XN9NOmmGD66QT4lJEQv5OWEhGXv8Z
I5p5fQU3O3WsCcTm/bn9Qw7STtCm1Gnv5IhkWTpeUHIMWSRWjYh1Mlg7u7k7xlUYHEBoHngz8isd
kV1k1nQwRrha0dlv6J3Qd1GdDqHB/QUdrhpHx3X6qDQneX6LVNbrtdtE5wNrK/TWfTEaoP5oqQJ1
kE0jx/SunCWRrnzI1wtAJqBa96vwefuVnZo6JVujlVYxd/okW14Kp3fXeMkZqO3P6Fvz01WjKutc
ZMiVZIPJdMsarp12qGB7Kfo14XzByZElbAEX6Dam+NAZDytH8wCUPrrBFHeuXz/lZjgMSI60WS0Q
+crnHR9Ejh++u3LYIm7Wz7jb64zahNUE9eJekPwLmqUVD+PVaSo9T/IuA4qSM5IC9SfFuMNieF2B
Xo+tg+SXfzdb01IiKKzbYRXPlrN45467fgJc30b27DSLylOW58Ov5cDnnMyGshLJHBQT8g1zcpPD
rlG+ERRGGCZ6G0o85Ga5VhdGf+q64jASzRyq9MhAcbo5B6LzhgLp+Cs1WROxTRnJ0wkTBysUjAvD
5FjQFzP9m7XFgUyWIbW25AH1jTMX/CER8H8JNbO//MJEFvDxrt2JO/x7riXTAjOlLDVH7XuPTTsZ
Z4SzFWgKixvjhm2sKU9AfsA4inMC3T6RfoCGZv2epbqHlHU38ff9wFGNVG7ibjQ+4nxLHeIKRU57
0/wAlJBU1f1BL0I4ceDHZj/hWMTsaasRyunFMwaVToHT1zJj0dg1XjE8cKhH5KSWX4dgRqAyf8MS
i+V1jY8E8VMMdTnmIyajxR5Yn1yJEU+WQ+aWSABwT8Dnlkfao7BgL5ZiG9hboOZqxQHtTj5VIis6
0OQ5Kp5ddksmGaSu7nkDuiXmCwbomM7c9vGNaXifkbT32i3jsoxcIW7QoKNks0IVTT976ZusQGoH
e+tm5/+OIu3yXW4PhMc6lBQT+PlnQUm283Rh3tyXT3EXgiH6q6Gq1GXaaJQ3HoD19lVDgrvh+/oS
waltqhu2pCgvDAnAHYc2kyosLDNtbVgzZ0yoz8ZKhunS/htnNVmhrzRYp4jAqeJRjTP86J63ZcwE
C2CsC/Re/IXDFnN8i4IFnr3gwxFzejEdgNxkBoOZsCpue2g2UpyIhWQTQITtOB5shvcwQwST/f16
jVumTorkVJkGUMYTgy4zH32GKGreuFhh7TBFBQfbi7ODhDZ0GzB7UHdcv08POgbZWg1BAm+VALHM
40bYszEOAueKd9r7W4Sz+WkTmrlC45yIpR4n5Ki6rZpte0b0WzQbg3rQFxmrzCQskWz/8UAlyW0j
OCmjnehzi/cJva88/LVS1xmT3GEVBQnCR8E65K1GhuY3bzhZ1B5qy9sgakkh0Aq6hYmr1Sf0RsKU
K8jprEWEV3tHFfHZhnkhPPNhwh8kuqRk0B6eAq2nK7+zqEC3SSkBmMlseDpRjyC4PcQvgBPR/Z3v
e4KX2EyW2jS4LwvQKsjA5UcOORHP3O1AWECObqBvMVy4QFldsnYAfx44qWlBuAMEMv3tOKqTHtIf
1eDNnn4f7QHKHx43yn5x91dm7k8gr/OPvWK5FM/NfyIRKSTdBzpnC43QPrxgzXdmdC/o+S7Q+PcL
Lx50ixqb/Ru7OIO0+qR/3+ZzclBEIXQuP4KquMuX/LnEOGG8qg8c/bpM/Wu51/zAtX19Yen6pcK7
p5xe8cmzzZuJuTV/gQIA6pMjxYfa3fbc9wTfe+AtSMV4zuRdC9wZeoPtpRLFoGAhxaY2GDHiPtOM
H3FdIVL8WhtdX+dW6B8FGNxdkJTxZ6RYFlAMhJXG6VIcgghdQ0c5ewBKtq3w0jjMWPWtPh85FW8J
hsNjDWsMWhRXY0sTnwYiLUVK4dNOZVmHacePRtLNOyRq38HN5nHzrQEaiMPUvD3nsp5akWwNjNsc
NeiJMld29xtEfJkyQgd8sp9sD26q0DxWQUXE5GwbsyojzgYwwjB4C8qOzuE/xyXdg5vqDtQz1N2w
z553iuO4+mHLUhKa4INXQnek3T+8PzVd0FQgWlDEkzmKK4GxMIu90gQ+WWd+r3NZo9q+M5Eq4wuw
8EClTZB4ppA83G2EJdCa0acZUShsj8/qCTN4WzmU/S5H5G7/1jUv+mL2UQonb3jg3JQQE/5y1fGd
rySjayoQYBf+XPUdBTfu/ICWVSxQdIEol6USXmzxA6EqIjuHxulJn2sKO/UVczn79PwnbDdnhRdX
v/3U6XHPsIiZ2QE1BHVJ6xMIeVipa3ChHtJ2A02ygOUpOFhrF2ZDvP9v16USrCnPiIpiPJ5urAbK
rghrO21FXtw3Wy48YeqAt4B73TGReLzF0OacSBk8JeRb7aPKXfj1gPaOOlmASTrJH8jUbSblyaUz
9/7T8NjwMFFIs/2a9yN+krGu8W5WnMwTaRaaMHIc7/d8niPrHkohOT5wwxvr21QdR5fwinlyblgz
yIQIpUPuCbSCzIlnn4uVY2XCypwgLG2Fgy8qQzNLGpUHDJMVbR1toi8KBx6hziIX3ISmvKXdyHry
SzhaglxCoQd9KrCndQyrfHwOnnp4q2fk14yXnhWqoV3OLzxTCF5baq1cg4MBPxRtZH36hcU3ufGe
V/UugBoTUAnttZj7AfI94LgUkpbCPtIywBq23Ae3azkM58kiGWGn7cQOdRDRHgzy/BMHzeB7poqA
KE7CV6DzDj+JvNDzpIJdckIHEVT2fVMoXSNwjA/L1hZKxeJSebmTExpGhF5654V3KCCrfSU9G7H8
N4aCCsi4U9dAS6hwEXpiAqXxxLl1sooX4sYQ19iOWZUmtiG0RVZoe43cCCM5qjmacT7aG5fkMIoT
nSIyxPSz+ooU1dyjnn6gKQEdgDK2z8yjeAkfgoprLe9lBuyVilXj0FDhtJIe9qFcOq99zjN43xrm
KTAK6UUH6yMHp7Dj79g6BBEr6xjksKhKoQoQSx/gLcS/SK+vpGA4xILEkKbtB51Vj/ozpbAOte8F
6mJeDAKnvYJDS6l7ik2i+n87t6dAnG/ESaAgPaN+UqNghE01N20Hn8sozGPK8EbV8Vda+WQq//VA
oQVb7qJsxZS1Wq/PrbpzLiE1cSVUKXuGH7CF3128K13JydIXgI9E5gJKWLVGcPYHTky9D42B3Uiw
XOGkr1t+EgyZZIS9ZerkotqEUlQ78ihOeboXA8RrbC+o0UhKaZKw4M8m0/qEre0vjPOoV9CRboG4
RUK1Yyg07CYgF5iO8SKvD7GaJFR2SFOV0Kh9kTdm31pY4HuavzY+mM6sRv2Vu+qqR2kQrRHW+I//
iXu5AAEJvniZDE0X6/6G5akQIDOeh+Lm2pZ6HWMwUntHq1tvlUaQadNKlLFn5ipkNPnxUegZMJGq
rUdHdJTkTEz5u36n43kvb7J9MKwBYooRX6hnP9vcTxgWyB0ZPFzYkFoXDa/LTDn8/s//y96fCojx
PNOZS2R1sBPN0b3/hFL//RH9AXGgeQ3lARD01yD/haZ09ACr7+EaZVxoWi8k9V9QiMFpN/UWJEYq
92QZ15XwJcPORDU7cQVp9eutZDek5sbDw42IuOkq3z7jJGAh1XW19/M27I9NUA+zj0eXfWrYH69s
KiGgCgttPHAzRv32O4dbLTdx4G53D6gjpThivi5r/gKCc91ZmOOirASxcjGK+PC6MRr5HUOVREDp
xeZnY3++CcAZoVGOdhz8WVrI7T5/vK/eKpGzqH8j+ElJX8LtCjtxAj4SuVQlJE7pC3McFXSp7KbB
Wox3y6BNixa1Ox//kbj7CT+ZNu1ZLAqaHBMLgMuOJwXOpwKPqzW+PBuOxpnJxaBZJHxFFwkn0hN7
P0WuqRmIosyzeV3/+o2tFwO4UtU3AX039hYHpC1vXIYDBcUkkTfbHFotu+zGR/h5Ml5bfEAVIEuK
dBJgI0gvdysYVYV16XTuXlJKXoDWj/dMt8+89le595j40tzjZfK4b96WQwiBTg/KwuCetvqBSsse
flR+pNybZQNSiNpxv+i+soO3MeyNFT9jWLo82eDKSmQ2Bg5Rkjjfv6XQaUvVFyF3/R1C5eiZLmhU
n1IARPvXmSTibrF7ev7opSGbZmboHQKIKUpyy8VIMqkT1QpKo3Hlrp4XsHAR58Z4dBYDPDoMKFV0
5OepO30fe6vr5wgpXIPxz3p5dPOsomWOF8s5uMb7CRXfkgc74ttgZGWzJ71UFHFO5l984D8B0VQa
LPrQzisV1LoCITD3BH9WW3SUVwz22Xah2L0MRKHMgH37e6IWzRfcBlX9msRGroSlCIUBmz414J8S
MAS4kUBc7sNTOZOIXB7C5QCK3BMZ+jI5XdQHcVii3hmm7dN1zAGgMWe21Jx6Lm1hbLFSH4MrhQTB
K9vGuMhJro1kD8WRwlLKbQ613j86oTEvDufVbofzxDJ0auY9fRdK2Ammqd4tFOXgsybdTFfjyzLn
9jrok0wnpvBjqhZmwRDAKbsoDDs4RmOlsU2XrSC9DEe6doRtPWXOzY3UFPlWGS2s8HSUXURMqodq
ltgCaR9Owb7RiKU6VC7/Z6ogVuVNv9jNZhakTZaTO7IeTqleca06CLI6EGt6htVncqqqzz4LwVo1
Xu7r5WxLd7ISWoTI8+v0ilp//6IFpoSkxO8QndGS7Zp4zaRQfVV5b4fM+WRRiYDMkihedf5V/3s3
NrdKSaB7/hwsEruGLGHCki8pS8d8KsBuxo8AgtsyuHO4vj+BaLCUPmSPxLKVUf/gE9JS+NqVeY0Y
mzJA/2aY2qJ0eHqWYCGW2ZG5/QOYdrPkFIU3luKg70y9Pxucxii2Jn106VLkE++yBoMw0XJyOE4g
Je07NQ+JWU8CAeCoWb070bQlBjk3PNjOPbaSLTXkoDzN/lh7H23eVTWN+e8DM+ohxpmINdmQmQhJ
5afrvD8pkF0NQ/XepXvdqbqIxd4KlqpovxnbVp9gZ5JTPjXU+sANKJYgU1XBv+477HUepcympUhR
l5xWOT6GmqfUFiO/sV64/fNnYpBbDtpnQFnTx/QLLUfKwdVJo2NaxOzLKJYSezd0MN71rhbWF64q
FZ6u9ljDhy3sbeBGxjBWdqenfTeZ2MKeLruVHnGuhPrA55p8p1ifvEtNl71LhuczDFmJl5VxdXHX
gWtA+ju2nbs92Y0v5ug+kaSHB8SgM5JpraR+6NrsyVg1BbvfRwLqe1W3PqeePzwUtq+r66KRPiJ+
16j3+O6D2C/DcuK4xxvBBRKXjL6JhzCeERhvLNIhTuTCZy2FjS2BQtGBNjj1Egzk/p6rP9TODiVO
f7sFR6O64DPyxPMxCunBDgKGlkw44vTg7R5nRchtMtCLZ5teFpmG1cOC0/t3O1QJkhxmv4Kt0ItP
rfRfth0TCwFHaSF6PyODufMqP1GWDSRPWLeSUC4OfBn8S4SFbFSOUu+9At8rYG996UT05R1j22Qb
TLZRBXrG03wEPpsfJ1qbanBMYhDWcKm/bjdcQw8O7L+d1+mF8nPW4epJsDwN7HRjFg9HlVXAKwLc
hAgEzBqqJ2bLGd9ob0W5whSsQUZJxPEjvImcgXeksT34nu5CAu6uKV1QPbSndJORMwjPRuIqzrvW
Uc8ITc+0NQkPS9vEAZfUlvZxaBinJPBO10fJnpeTIhXgBYjMPDmB0e0pj0rV5ueasnzTFPGrsdYa
yZcZ3ff8DZOkeiL2RlWowX+cg3SsXTZj574mfrpVWEn4z+moNWjErEPISmEHGEysSxftzQiS//Ix
w/zubH+P5Be53ridu+MwWjiZNtZ4wDJEsRVPtId1taZNdgo07rAtESnV5l5zT993vMztvkgOzT8+
+XLsz8in5v07XviKPSus4/erNGq5E5KU0JdDlpsGsxoIrcMKMlyjPB6pitTcnM3X87M4sOVmm1+2
kdGZQ5e/mkJ0N68s1OEjP0VcQoPloXiPiWhMuHIB1FW4f6pvSsDtLHuvrRrxqxR+I/9wXNKfIZIL
X3LD5C0HwUh8X6l+otIl4WS7aYENlt/xrjKsPqDSDlQ2Jiv6UpvD+fGqgwHczoTqxg0HooGLiNZ0
1qthvWyip+Hd+LDRfOG9S37L6ku8W6vQH1UtymqKZZARkl5/d5ZExxpKJT7GMJuIsahuqIfuvtmU
GILAeookG5hLAGUkJUwKgIO1OKsvz36tsGw85Ev/z3JVDI6NMACCvPFMVxlz1co7jdoFdnUro3V+
Uf0jKBHXlQG7bubfqk/H0s5Bwi4g8f1nrGPCZeqawtAp5+MjiVB0XIiHo2em3Mcpy9ePUYjcDaou
q0V/4lGZbQPvVlpikcmhQiDiO87zlx+X6pzCurv8CIC2w2U2uhJ81Ds2zzwoJBpP6qCOZkUnoLnj
iuW/NhjmjotANM6kKQV6IXzTLvnla1UEKD4OwVM3gTkK50AQQlZSTIFMSt+8KTIbOnWb38CrdeFv
GgA4tqaDlQBWkgCtjyloBNMDpAsDhTeUIZQzv3R1ZFEKGy0HSMPE1Ehda7nGibM3EN4B2AINg9ed
VRF1wQ7wL66hcT0isGFKmafMRFjhi8RJwV8ZJw0EzfkxqyHiAGMmJt7wxEumzCA6yiN6GKf2+9xj
r3C4hPqE0dMxgkh1jTgpSbtFVZLXLhV/82uA3y3/6YoccUK+22WReIROI0DlirPUb5uKVIHnU+du
eT+hQeDh+CQ4uBpdssUU4xAr53SjNIWG5ety7TrB0ndsbCxiWgWLtQT+AOaoxjJ3nw3UuTTmU6PE
zU3fUqbnW0JC5Ac6yhrfSbdg6bGIrWjHS8/etnvrGGLj6dQgGxXNRba8La4bxCxEDfB3YWftZwsA
YxeSX9O1xe00QS3G6NjNQm3fLp2b/Ln24GXDpY1JrO1aayWnE19tnxITLt7qXlLXB2mnPdv4HxMc
ZMo9KlDgAnao1PIMwNPunG8Ba8Ee9f4zO+eVODJx6YkPNdp04rJtcIIk+YMnw8n6ns8x1jCcnJ7I
K0YRcoEN5Mrfkw39nuTUEGbmDs1HPyb4w97N9p8+7J2FJLeEtDFcP+yEqfz+2HrLt5zT/cIT7d8Y
Gsy0Y8Ttb/a+e0f2tjemyPi/NPyV/7r4vFAev76EESizzo0ZDfhgiL3VPk6CEJLa3GgOxt8kS6pC
tmrWKblclTi86FDVjj9/FumfL/YB0tosL+JGUKChGHCErTZv/r4CZ24M9w/YFq2dYcMn3L9sjT9X
s8uJN3Dwe2/Vk14R8CpslHP/d/5OMOUyim5s7eQ4h8tm6eZ3/MQFPYiIZ4IDMm+0MbJz7xGF/dhs
vHqf7RFZS92ZHn7FknHPh1A/9jUrrkcccvMj93pP1YoKOytJQy27M2UGzXgwLxbhO8SgRCln2Iee
o9rE9z/wjFaFaE5Q0FYtpUwHjnGTsIcrZCHtT/TTHwhFg5UIp/yxbcp7NDvjWApnK9FvHLzqwqQ/
q7PJ70iyleR45NpOX36HGxq5Je6nRAKC7qoYLAJTdYWfVtGu+moeo/oddDG1nH5N8TfLtp1tiLUG
NsFoMfxpdbWfCUk/csh/zkTMDR3rHo04u06djmEDeC1To3zW19y8zo92XTPIh3lpbrZBwspWFMaW
xZ9azKpyyvvS9i7nX07bCMyhi9Mr5Z9pjKNqVQEBoTDHvJjjyffg0fEQ2CfL8ARiUv8q9yqet7Ui
oLdIEW64L0fS0xiJoJARaSwDLCv2pIesfpfv7d2QKyOT9hSTwmvv3Fkmt8k2ai/IC/xMeWqNQ1/7
xlYn/pE7WdqVApGETXGaJ/i0X6MQNilM6b0cVV/rxRHo4VLBInVMEhYJmAvyHck6ZASzcAPyKqXe
kxbvpv9lRRvqv+CUcq0yQips7nNrAbzgP7P7tsJCPVCWj2O54Jq63dIt9jQVmfyTLmZIXTxyXxnU
BKfFcyI8v6n1weMTUv93gPQp3n/q37V9U9XTHFT97Hso/m6z75cdK8AA99LWkOk+422b11GlIPRr
y/V6dEpmSqkcDMKtwwXrXncNTPfBSqo9Z+qkPQS83SXpWz5k4oV6fb7lFaghR71B89YH1q1q5Kiz
bPXJbHyK767m2nRXiyzACv5AgNiBGh0hM75NNRGnC0j55E7UumX6VlMJr/GUsrl9nTXasEmcELi7
EKWFueg8W7POHvzY9g+70FJ5iMssD16x2roEEQ9yR6uQ5XpqcNQH55MpkkqTrko2YLjDADV1oiXt
8xz4QeAbvbOHFQAHElLEmNnbN7qcCzVND9UnvBuHvCttLSc/mwzkoaR3sIya4Oc+boH48F7rnPUL
wc9RLP2/knBys233XMGHCnPfbknlPx9nZSovcnEMog9aXU6GWES0WM1E7oJdP+bfZ2L1pkxEMo34
N43wHHBA3M8QgJrt7I3ar/Rpd6x/wgjPbDhbpDONLB5VzkrTUPQEcQWzZcxHPM0LKIrF789oXzMu
RRvqzPWDJIzsNv/IesUDTnFagP5yGeSZ2LqDUgw3LOH3QPVshJ026a6JFWJPvow31dwO7LwnYG5Z
ZSQnWV4ODfQgzw1oWWfKtyRl6lgeohaXHyyt8UMtWopAb5C2iWWH4AFrRc17gj3pEIN7lJzKDaCt
/IYTFR+ujvsbAUsu1FEbmOOsgBK33d3kIStJoDpLRw+cbNvAP8P25mTBLmMgOQQDMoqHcv+Yvatd
15vW116xTqJwW/d6jZHseWtZhIoCc44sWabyM5y2EYgnbQdM+Sg8aHj2NTZ+YlJj3h029hPqDS8r
7EgMQj0J9JOB0Z4Lg66w8agR3AZ87xW2UDFSo7tj3LuuBQ3fivHKlRySoP5vp1DEboyzxCraf0PJ
m18OawAUDHfGlFq9XocL+ki0GET8yemAmp37XaDv22p3D8jxNFsm1E1kmfO/SSht5KnX4OECTdM5
TWBS3qDLPlydi6WX4u/xI220T71sHJHGEnqjSp3nrXXoYnBwdcwiOCIYsAavCaMSvYry8PGMdwXC
dFxIAEWJVV7zCy6YS3pbyex16J9Pc9cxnfVzH22Q2IuSqt4UcIPyN6s+VuknMbWxxUGqIibpX46/
Li19kT/xc2W8HWuATCPBDXQpgX1qfH1G0v0JG65dAh/7JUYCVyZefoKdRuehfPLXNjMsNzJLH0AZ
SgMbfJMJUtUALCqqvKVUcl8SyYFuitVtAUnAdczqXK9KdFXpt6MCIP7JOgRm9hN0o8F7hhFhMAuY
GYVOSbE/p45bLL1euRVhIj8U0kcUeFaohVHkz07sUDf11E0Tr92nKpi5zOQ/jSrJC4MtEE6tqE4o
PkVLCMZ31Mitzyay2fiVtOs9l0MM+OvlBXrjVDrb0pma5H/kvX926DRHNHLyUGy91YditiEDGuYR
gfuAR+SjFwzwnzAy9v33DSdWuYlKhuGEnM2H6lKi7YDcbiFLfWT2vGd8xB3xgIBp/l62w9eUuUAW
p2Qv4vPrP3xTasYUWcwrI7GzGmglxuwkRNRb9zECsWqWkJBMY6axe8vN8hKYawEy9R7G/f6p8AH1
qPJu8eSamlpoI8ajZp3ubrwhIDuk+PMOlU2gGtzdtfBjq79D2K2T1HqDd1xoPzzadgRxIcfFXqSy
fS5hah83+IB/zme6BfTw+a2w8E/Tv2bWhMdXmpRkxIp1OUYCJ0I86kH41uvuzu/B3KQW3QLa2i13
yJlamvdi0+EjH2IvA5dyR9pBo7GAN96zM89xPEUQ2gxy/6x4epoC9MCccn0diP5noBfHBglw1qrN
6FnUaEQWZipEYVqGidUJY9RB8bAvL1Ml0zZwf+ergHhO8OR/0VkpheKYSzRd6a1xMNGPxI3mG6e9
I0+RUH0EW1PbE5s6L6M3H09NEeHpS6lMP80u+8qryLynR181lvnHoYiskhPnSI7kav2mnf6sFcpS
73uFb2l7avGwRZavMKFQH2C+c3YopnZTpE2lLjG7D2jb1UdWUKAgvKrePpzxs7QMbeGXeTXD7nKA
XYPHWxuYXi+/09BdDHXzk9QeQ0c1P/TXrr2cZcnNVq60QvFqpcjb416iLwiR5sq+2/uLslckpOQn
A0EpO3CFK8NjS9RscdS9SMHu8KlTV9F6/08JkyNDpL+F60/ODPbFBL8nkd2/BAWV2hZWnpwQlSKx
Mjw9ULQiWW7pKnf5ERDeBQO1d+LeL48mcC65NugohG2UZsQYSPTIU1XjTvDQvEXUJqwyrwIbiPMn
VzJiT6N+V8CaGSJJ6IiuRqc+e6CD9YV16iWz/5Ri9xX6rgMAdRr3C31gUEbsxGbA3d0lMW4NHRwv
2sWv3iOQN8oYR9t36gPVN1E9PE/85XpJBPbtQYAE3zxxINQen50sxe7tD6lZq5eVOStVTsWqMWkX
QGuvhp8+bwUvIQA9f3LelaGwhpsn+yO2sbYEpV0WEkPqUfe7oH6GHETi0qdaZeg6Cfbl6oSRlkqU
m5gFQf9C49u5Rm88B+O7BPgGDYAguH4R5BTrH02GQZ5OUEOaIfAehWhTLDKTty4OdF5SVlqUZrXd
QAMhccuggihgXhxJSd7TlGIN6OMAX0DzLp1s5q7GlWf/l5KVcOTqWvyYFjhU2UKvZVQ7vbsL2fgL
OHc8jRaiMQH9KByOXY8o9CURWWibGVMSm6s5SYMYMyp939GIn75Mox9TM/Kf7hreVR8JtT1yPP9S
rjxUvRaM6TQ/Q5G2h3ZnDVlMObXecLJUnv0aYtePZXwP2D6kO/oLXa7rDHIWhLVsEOTmDg1LF2eI
ePWsQP40lSKijFwJWL0C/r8+qtzipgJ2bWqBSyZ4zOQyFFztDj2dZ0PP91ah19iY3bte/RfFz/Fz
WLYNN1CLGQ8CUdnPMKuAshOhQ92YceDK/u5JoDWCGpb+Y0yozUeU5PzPJ9RCplaEvOBXP11vWv2Z
Dz4ooeyNCyXb7Q/8MmdB3oKSCTxsLC0MeFJo2w+u/2+WD8/KcY6BJV25j9uYmelYtOuDntw8zmg2
LqS/M6UbltmbLeSs671tonFyJUxSuXrIvu9LWofw5z0ji7sJmNqOgVUamUpeFSwJGn0UAVozb3AV
CmJEeh2Qpn0T4GCYA5EFt2uDlnxzAYCrDZZ//TQ9vm7k8FIU1HWYKQFOzqACyCUW2cpbd3f6/5/F
lxuFFMlVYBPQKZm/DlGG9/8oHyU/jvwijOaA6vPEu/VRd/815jE0AZgM9k2bLghycn/1ByfU3gCG
BCb0a+rJ5+BwHeiVTjpbqhzcWi10vt5KYy/q00QrB220VtVhB03FeK/2GCr+iPAAGP8tJj6g1J89
JF4ucGzF3Yju6gwAE5BUO+X+XMeFmjcyQq3xA9SraLf+9EbIlP6SjikU8AU3s5aAmGbU1ksk4Dsl
667FVn+ghgMeiYpA3XVSOymmkDreQ3F4ICtL6TFh+m6nnVwH3vqO1zatujVStWnEkviJs/Utkqec
K6WzglHO8zKfBlJP+5U4ofO7QHF0zuNwX8bH8pXGu0yu10g8uuHh3Oymf6X1d6Y5Y36SNo56aVy4
qUNpTuXLmYuj3uHUcP0423belRPhnj4uHD7N3CuB+G0JGMQmekjScqAlesNFMgzZ1IVPHiV/LSS+
negU9RDZn6lTBNX/E/zkiBdQtw4xEui2jSxLyVgBNs1+wkrZJwDxhCdx/PMwmnt9UMhDUzeTqtQD
cCxEN7rKz28r94QPh16O5t59RmAfvk1ZlQny9/Y0SHBPYy7JxTdGnu1UWisC+9QfPZCo5gxsVLa6
SzwAEZCdqrnCuCWSZkHvnmLa3moNXn7PHGPmEL/UlOWefDbPhbdejQF8DV2wi7kWu23J5ikIDuh+
RvGKRlrm6gpoz+HF5YvyENGjcOIkni7/eobESkU4PVSb5B8F1JgOMPiPxyvArRt9YpIxIu+lidwx
dPrJkCHW/lIStBGl9/SfTOY2C9tYtXnroRzagoVk2T9UjrhoAG/TuRnvvdt9ResKv/Cc9H+Y+8jm
3s9te5HMPMErm3sn8JLDsBPVwJiqqpJ4iL/+/aexlmrU1ZR444zP4kKi0p/9BIioaPOc0Swb3Oei
tMEOFXPzPgtXGoMX9Nc5QBuwBrQAbVlIVrUmb8BP56UbUj8CAya+1vVf0aVjfolQJ+6MdT34GXzf
FFldchuN0IXiopUzRTCzLWJvvaEYOjzecAvwuUpPoFgygIBcOxspYJbegb4VQzE6BdIsLw3MLoPU
WEqm4tMMC8p779QMCGnQufk/lr9jQQtYlN5b07AIhBOaeEitWHiR5v5kirdFuIEzH3Dma1Xaubko
V8sKNn/4y7pLXjwlpX5GqcvGuSHGu7IJzkBxubvIFXqDh0gQsdorLmRXAsKpkEr7o2/6cL2gbGNE
1o1OFv1kXDf86yYCUVDwczWcWI5qVPT7Ir6YyDm1omDUC0Zl2SdLmZowjlFfpGm65LZMwrzjOpZC
o0phL6xJy21ADinjAbDnrHpilEVCIsj8WkpnBhhAiJrW59pdaP8ho45VHapWwNnVX9KloNTGEyFl
+AphX8LrYnJN8fa+t28r0iJHsyKIHLVo9cHSjFb2xqIJl4TSt24oaiDXD+uzNSH6cXm4CiVUoyw7
UOLgPcFSXQ70p1D7Ajw3WvCzPslR1n0UYSh+KCHb3iPgXkPey7tLtL5PivhV/Wn7seQQ6o2h1TqD
FNQURYKtPCWkCjuwzVlQbUq9fc/Z8W16mqqS9HgiE6b1Gx3m7g6RRHXa5A0X4USRSL4AzK3WvGQ/
DBDyVKNMokV0Ksw9Jeckdx8HofduSN4nsZH89c+JlWXmhVEHdJYIGM0aNy00FFlazrh7NmizlgYp
S2+dGvkcRRGNmwE+mFwSOAS7NJi/1NOb6ZSCtCTu1daCTXCTZHy5tSieGyd5knMt/bg9uejyqajx
0urjLHRb9C/pvOSFXdwNCx73/H2cTJkl7ulL/eshcJi4TYUs73+zs2AmGf9vODYHepARJRdyjvsj
NS4L0HkaGJRsxd5Ku99RXOAdusyaSG5yHa5tuBcVuCUENTZHXa2jZEiocND8INyd0BQegRGABByw
FuocUCMhGMZLC8Z+NEc6rnxrYAQTOBGs7U1Akn4LX88RU+zaQ9uu1HSnh2Kvbcfae6SxWEoGO64M
SB1Q8+zSMm2FhGtBnIE91eSdPKJH6T2xnVYTrLmTliface5Lo8ydjHlenhFI8StIad4tTXPPa/jh
onUJE1nYKVCmrHCrUn1QL+AlK/wE6xzkBYUob9nLKPwAhEakxOyW5CI3ikKxh7wH2PU4+AAOn1tv
2miTRZ9uHHiJ7x3emizqxva2jfNcRVMRSoWgawo5++0QycKgVI1wCOG+J+bPu0rH781+joy1P+wB
VspzTAn0VHFB8nEbImjaA9wslaYTnVT5SFS75G8kO5751eEOTl3FmjVdR7aWqRH7t+00wqDBUtI1
HESv5UGFXZsE8cIIVX/FSxS1JKMzzCpj2daSRimQ6FSeOzbkJOv6bOQ26e7tfScR0FwvzYGsjOo2
nayR6TeSl1Xg/9HbReog/3/eiZDTK/u0gDNLc4adyHr0AkYa0pPP3cxhoixLeKHKoqJibY4z517W
lJFS8s/3gw15s55DOFzAsK+8z0epE4sF/mpNv3evOPnFjJsTAlMxbMh3TZWYaUoG+5JyeKpsa2mz
+dbh/z5zpC77RtGfoBzbvilAomBIK4qwdpysIuFak0/r19JcS0GgOS7Xlm9N9G++UH/B6YpehL+C
mCjWwRsCVhFAxbJrQB05NreZ8YSHwQybrRwpcdEAtEEXRYAG8Ccodj/HrnkjvjJ9QHxwhk8j2Tzh
2y79f6YcjbYeBtbF52cE0Xpt8yFUfY+GMmm1Z99VEK2RVXD42JZo5Q7VGKH0tNDPzUrbROER/p6j
5+KVEMNkR/F7+DUTsNGezD1Najs2YLaGXUmLld5hwbJPZIAZR9ft9dz3eXz8YE1C3a/BBictJ/Xq
QMuR/f70ZfwB4ozrW+g7xSlqDWPiZ/OgRK9RUAG1yWDoPMY1Dv08NsZKyUltJj1z/H72ly3mk/2j
kxVXsxMm3FcAeBP/qsazRMBlLIMRQl9Nw2byASlvu9NbD++xSCQOe58XgKqfhY6xIDDeoQDcIjIq
NY1CVLqikDw+aSnpjYZHbBJo8KVUw83o6z5CriZzJfyufJuObkYx1LVcFqrh/3tsS8xPW1fzROfP
g4aL/Lj8irg/07Qez+lGtMIbpHhmlLpEBur6HI+IoKLrxVrtSvFsX5Y//ia4B+OfYb/wlcxRY704
hB0RZqFkYA6rrUgU4lodR1l0xElPDES5JLgAaEJtbkMAWLo4Wm+tTlWc0NJ/dWsw0rn2ZsUEufLt
Vde6GbW9umgaihokipgUq6vxK0eBzd5Ar/OY3/XMjXQzEUH9rzNHMgtG/wpMYms/VfAxcULzjFbR
q/Yx49bWJ12v5GpM+zlExdOPicNGBmwaSMrujipE/zoSVF1ZqXAnGl05gPNNwFUAtT8P4UqbAqNp
Xebs8g1mMZ6s0xy4l1sMr39R1y9po3+SjOSdE2zVB+JTvkvgVtFXk54KqJRrgHF8aSIzBODjkqvG
YZFv8TbnmJjwhBIjNLb2yrKK10A1QoyYBAafA+l2Vq/Tkqa5hz0r5/1c31IPUMQrlWzkLbOOetQ1
ITdrfzZSK7M/UKmEkfgEadiI729M/DeyIeotLrJTjGMPXII9PMVDN3fxRTlvF6gqSGuw6CZR42ns
vSl1UQ7V+IQfMEQHQbk5tK52b++Hh1J2yGr0vJIpYinP/nxaoo6OULhlH7WsIgC5+llff9Mrf9QM
dWdck3+2Fy8gWeFFo5ltRBP4iDOxZJAQubH9XKz0qURFFcx4jrKU8Mjg2iWOu2oRtQ26kb0fbL9p
3/dV2Cyh+0HSynZRmWuPlQx3lsEaqzd3+wzJtqeKuOSFyThgcf8HoAo6cq9duktxjoXDeclEMaG/
74Se2J5iQX9NtArGFY4/rfXhBQo1DpmuVgc6MtR7Q4vrDjNJWPVahq1d+BpwwOvwA4O6jBXMOSSv
rRkDzckq/PqQEahw3rNycT6/CKgTwKGT1kEkyk79rizz7JZFMe2ZmG10VU7i7/FqNDDB4XW1Rh04
EZ4bkHVR3/UpHEGI2USR2zUSg26ihiRUbAyOflI7dAI5Gcang9I0k3CYUM/6BiCZMHQyQ4KEPY89
OarboCrtbq+HhelFuVGJ8O4Nzh85JmFZB/zOGqtPukDWHnHGuro+tYqs10hy6DaqP1An7h0Jbslt
NmnxdFxbFj9f6G/0z1Aj1xdC8+ZBdlbFfwtXTtvr/qxyMfzjdWZ587gRjHuRqdD/V2ddwNwdIPUg
bMS4oAEVN8E1+yEEfYxU495fTFobrAJ5v5NBVDo6Rd+lUBuwWsIE/efTU9yuypYCAqcwAL3biDr7
9jcN1lsWfmFYpAcOc4BS8/WVI6/sqAVldla/Y9BCUVKQn7z9oDuGpbRA7OVEEeTswMLQB1zjjbK3
+DNW86wbYjgqKh3uide/j6UX6CvZMbH6UtyYtKPuR1yNumnR3Iz+sZ3B+fdDU5ytlzpI2NnacelY
3gQObjH1gwbP4gVuW7vw+WQY+unV4S+ShaxiBeIQ57DiRG78RHRq+uCtGUSKbVTGj4W33FOaI09M
qZu02fOeBuxgIpnLIr8X+Hvx0hE3vyEfKkMtfu32dDt0XHVOPHTzjlZiAGrMk4HCp8UrtSaCqDeY
zZUUhqmlxmRsWKH9o6EB0qijA4LxFHSbxUkRQbN5fwWRtBMOcNdExxpHpx1OwgtUZSNdHm8nvWuM
QBTUs2b5yBkwfbUNE+qGbdVigpiBACOsVpLp6xbKfvqMtm5TUKFOr8O8ck5Cpf508daSlJV/Z/1s
4T5OlgpCBMqYPdbPoh0wztyQfWYikk1aU/LEB4tBxE3WTH+npLKWdFrqEC+Ofi+os/dUY1T0Oa64
Qdp/Feoye3VzP9jxsU/DpqB2UQzMEAZsL60iKazm4Ys60Fa/ETMVFBHGdc+KVxCHhjw5yB+YDd8E
NAVktaoPkzILTxS9P/NcKw/mE2dFGpqDCebp56HBOViiRBTb3sin3JtD3/2ZNqx411MDLd2HPe9Y
2Cg5FP2FJd3xEX5w3JZT9Dqi2RoTiWkUsUaDmb2encrfxaXuFyUa3g+M8Hz6CuoihX3PSrtheeEV
aBGrI7c7dYWFrAZ3e6S49C+CE0DBECCwHC9qCChzdGdgd1qktPpI+CYhU4SOInzhjIMH8lRWEm5W
JGScFN89r1QB+5Xi9Z1DN66Olr9PaS5bVFvrwSxUFdYzeCDOCWkX7W0FPs8IEEBD8zJi6RI3+tDc
fRaqRGtUshFFxKWXI/LbuCTg+N5SiuIX0u9Yvj3W/Ahj3GgGcjE/MiVLePMbFSnWZlckj9+1ngkn
zvcDQ0YCRPQOdO9tUdCFzscHPksgVuw0uiD+JZfUTO58qX6dBFUsRq92WrGvQbVfL4InJHWGKoU2
Lf9hMO1zx32FCni7GVjgBKC1L6u0R1zseWpccwDLxWzQPhQYE5Z9Jsv7/0XcniPizY3ZIWcapFhP
0awNrIIV1b/f9pk2KOB2/KGSA9XQi/rn2WJe99QBeKEzNgEMo1pW9H8QDQD3oR5UH10bC8EP4Vvk
6kmI2HqcLxkk66DRecaZr2B3376sBli4/PsBSzoQbcjtx2SBP3c74RFjN8Tb2EHYzW+JBo7vj6EG
YF3KbBnOz4G1CWhD8WYJml33PAz1GQDz62TysX1JMSNUz3eMTTxMPSazUyjqpHk7E/rq2KUu4hx8
V0p1gvfeQ0S0zUdkmRthFtLZUsEhCeRWPJEPSO+y7z9vC5U3bzrkThMxXEHhrWCn1+/6V+er6dXV
TCZeOZVvdHk8MbBYVEsFUcDC61yVZ3OPS9lY8qkiE3mpNk+O4dv84NLyUWJyveASJWcMlfAeI4h+
Rjgud/JQLxEmfNh0P5h9ybP1Cw2uvzz6qHlhL0EabbtTwHuqMzmSsl80FhEZizYQCqzXo2ueSxMY
IWi5fDasJoLIIczNNWF8j/K+NAyzF0AQC2jQ6TwTjTYKsSHLXwPpBQVIjZrM94HrvIhUqaY9RTWv
ZrJU9Axlw4nVvldH+edUJ6mJbTjQDBjUF5l7FRWJ3bMD+mXxCTZnetSPTVA3WA+TDZVWhXEaqu/Z
oUWVn8ze8PgbTB/TsEUrJzR6NYka3I3HJQ0JqOalgVj9iny9r0j4IuwOTA4p6eYsrHJQqjoSZqPX
X18nUqIWUy86wHiGrodZJObwltw90ttoocBShEK9XFPn8+WHr5mjfyHaonfiwYCyNrYPsM/ISiSF
IB+mZG0sk++fDZ2bG6r9f3WFRe+dDo0rSlgZAernMByIQ30u5gCyIZR8NCfzY71iw45UnOoE1ziD
wGuSt5hhZAKkftiNqsH6ROQSZ8HW4EhJMR+4rzQOBFSAcbVgDosFSOzTDrdJ4bwoBC5Mod8VY1xm
O/5Hv1brMFyuacwzWXId8QmkaBFJC4+pWqW9dc3eYFAzJr7a7GCDZPJ2tLPew5ITAfVJdLwOM9in
er1dnnDDjwitJhsE4p6wphs+bvIsvM0EM1USMA0J3lMlnJhJNPrIpMjR6QNvlwfq2+AIm1J0Eu2y
FCH53zaL0cHISwuy2jEE0RsJF79edv8qnot9bMzTs3Gu/SDrODst7g7YWqLqr6ABvUQ2itGy8gfn
nP/xvzYOmtJTVVQbbilfA/J6MfLFGWjXjEu5KgsBdFL61wmz/JMbYYjYPlc+M7sC0yK+dB48K5FH
UlCUty/eYWh+hjAMF2Kv5ZDPiDD7XNxoODSxxGwkDDrMCT3YYOBlc+YpirSMWhVLlxhOxHcR4rUg
qUY0xRN3auzAEKXEK/I3hx0Xj92DqdGBzTHS7DwbNKIYAezG8Kwaa1ag4gfsMkoezJvnK0/z2LdL
N0T3Wo/yncZXGZNFhPi7NUlM2kTaSFIyc/ntqoAO/sgsUJOpvbwhYEVn8ufgvks+HyuexqG77yG1
mY60jejxxxyasDuLhMnD2EgvxF4TGevs8yWcrPDly/cFEtOu/j8pIkvrS+h2bcp1iHVdXoUtFcpQ
UQ3Lt6yucb6hACEAlB+ajcWa32AKSZqDlpIPAUk9Bw7Szp8Xole2ZFUeHdAgaM2vKvxSz+X/Dlyc
IyYQihedrMi272RG+ELFVMlerP6hwQK6mDoOGyB9mbkz7BKBaMnkRao6hTR1P1WclFswVDmKD8Zp
0wHz+6LTmCPmc9vuq+X9D5V5Lu4HLx8hlzrOTuIHrL7jAtY4ofrx0P0svuexspO6NKW1UAWL3oNc
MgZBHQCTV8EBYlDjrCoY33yXVxSbGcselwCE8uMGBYtp2hQMPgtp8IVoqLxaMEL+7hBcpcY/ftuR
Srwxn89dukuTEqRwu40qiyY/tq3WmrOiMLjGHJc5IjG+tZVJkS9txA2WmtPUvuvpuqV9S65Dyu9U
Vr0phZYc0ytRmkzBexqYfKO1fdOYleBhtcLyfYxwZwXt5uLZh5x75Je6VaazU0DC1lAy7TPY5uN+
Uc+gqvGB1ajtkH9j8UtGMsx711hbcIINsIyMf5DseRVq8zpPXNfk6CzqXX1e0plCP92eROAlZET1
dOC/zPPiQBGSmsqBJUzIXFhuAujUyCxWb3D2Gl5Z+5AOJQPZGWjvdZbmWH8x0OT3pYGBpnxCRHPS
c02qY3s3OjziaJFSEFHt3e1akp7HWDc38U7k3jWakuaMyXRu0w+SXEbI19TE4FVnjiQXzFC7qXdA
dX6h/f9M4ktDcI3WTRfbmy2RZDksBkvHMvDOAtSYcsEeS4ghCZBCe0WhdXLJWv/Rx/HnWDtceYYJ
BEtvl2d6B5yxSiyqC7ophXSZV4W8jVK878ChRbjnXi62KWbnXK4tA723QbTabOgWd4RcB180qXbg
zmUmG6xwq/QFQLLmPUtdPUmhaHGQNTja8jKWvopIO4tMg0SjU47BRBn/RfMtQdMfQAlOBhg8KPR+
+2NEa4Myy/F8GSkVyDucOomAdNvIKfa8DXowrsTepC64HhTO04Gy4I79B2oXEw0hYmtqhJfJz/zH
4eob8wo52IAJec3b/g9r5ojcuL4btZwaJmpVOKhTPiiF4oWW0YUukxdAevTHxRvbmXUXsb/GPRhq
8GQdCP86fd1Qw2ijUKlfqxA0Dd2tzROUyOsTVfNNSWZuQk3BVdMpcRnJwwSgIpsHXJceeOnicvXF
twYHLh2G8JTmao4z83vCRoaJEX4aDfz29CC8L61HjBTO6VCi8H9bkiigP6I6jiRBkLLiGphllpsh
6mUTr3lkxSDAjnB/Sqen+sFJ+E5nEjYO8BCC3vquvoMl7yhdyt/OoNEr+Cz7b8MAPB72erRgP+h7
Ai2dNVj3gh77X0YLmBEw1Ju9TScRkyQtMXvzsMVS6aznzA8+oDlp/TaWwBtDAIdZLRjlbmTXQyCN
yq/Q7TkX6PY/DNmFZfnqvm4Tzq1fYTtEe3RdkoV4xrewk1/c+ylKRZ5mgA3flS+NE1JH/tYBiADd
5ubISf+dnOz+YDfHzITUpItrAdarANg8VMcgfHlh7bIqcdOXRkrcE/QeL/qzJZr+Q/9kJPcawAe8
+H5HngoPkDwVrYph6s11OTkmrANchV9EpwMUbGaCI3FrSglOosJKpRg+ogH4Ewauo4MbQqSbBWni
UCKPUgdXXggMExzrOMBNlnyp3DadmRT9SVo/t4BOVW8lE6hjWpNFK/m3ExCjeS/RorpC+48p5Zk7
zM+CArq4WXrYuO3GSsFqmTZGF2XelBJwAUWcm8YDV0UJ/ebuMHnk7BTrJs1KVk2h2KhMF5EqGebv
veAN3nAmBQS1VlgM0nFqB8CxVrecfZiOucT9S17S/5WY/axFcBzia9Ez9Jfca9cGu6+XwWKR0n9R
baEEL1q1schNShnjO/xhu1Kpuyk36yDkWr2ILjNQKQpnTE8VbHURmreBlJhzaUzwKu8OPibc8gf/
jxdbLunmDIFQSLIRv+SB6Ch4NqqFXZP7yDImWUoTaAXYo/7h47IqLWm3kwgjBwxzwtgQPg4DJJdM
MkTDiP92HInQCkSZKqkKJuPOjeSx3tsBe78EVO+dVQdrhJzF5hEKO7ep8w3CJvfFFqGPn0c+lmEl
IWyMS2bLiFA5HHPrRKvHn01paZ/jThalc8aOLlQuaMSVZhUKpq7e2P1uCMLio9678OoV/96AnIpC
zTfVV0mWOlhDJSG/FA+axTXvRdDUjLObQNdl2LoEnlfwaGY2l0zCn3RnKleDIfTFZ4Sjpw0nLvSt
XjZsC0cszzR/BBWQGcwhcGcXBDkP9Aa2rBaRszt6jGkPjzOuyqs3ZE0L9e2KVk19owwwWsrwrf/F
jSv9kCZMFb5ll+xwSQ73EJkN/7NIKApgNujPweuTPR/CDjXR8XnBUJQVY4lG/NpU9mJRxVg7qFjg
3+nSmg5R3/l0K8iQeygg0evxceaxvrOCBA7Ma9icWp3fUXXLBq2BMoMzhCqggbhPgI3/S5ZDz0qb
KygxmnkVkkneIn5QbBBWBJKyOgtEa1AK7hzlz527ThUKOErE7yAHDWBV+7dgafP+J06Xwcx9fn6z
eAgw7yGCME6KDgtRJpifCSe4hm78vwvmbIhHNQ7YyJgCPni4MWueZ5aSyp5IBVGu3cqaCTg3cGJF
+haZF9to4CZqpoYHdjymV01QO9pXXJAb+oVjRVAj7C4WCl5iOhOqYkKqDrYJkRl12+Za9pO2ZIvz
EFu99InpbB1StA80hjJXv8zNzGepzH9ghv5uJSiLo5gIKsCnbtMe8X1b5ia66N5kltWMjrSHl1EV
l7TRv416AJIgDXD/MnB7t+Vgl3cqdK6CmnBXKAmC3UY7z/SvGec46vYVowwDnx8CdYEyGujDITmT
wMIfsswai6QCB1wNXx3mqkiPbufRUvJqrGR7fAzpnOGJ2v2BCqS31LIEu9WuW8df52RBU9eGdQ0o
ChrArqGjaPVkF6U92pGZIik2UxslSqr1F0McolYAfqG0LJnA8s7k3+TZAbQt9so2SRirr95GMKOb
3bChHqKJbaOV2OHbi8PuDDl4A8eJQ3jP5IOmdXYhb3BXKwjzU49lz7Map6Q9pEHsPb24GItG7KzE
yv3vhonGq/0DAKbJu5gYjgXnG8v7+B0paih4usWYdLzCJK4PODuNZEw9KZlj/4oEvreFEtLjNJxO
lmrmqPQsPv6hoFn8nb4X9VvOQBYyh8zmAcsv5+GWJw9fUhnEjSzrYnXQaoJEDRun85jZGXLqvcRr
5Dx3c6xg197Pe6+FOjJAWJ6i8oeFLv7HNVQsZyxRzUIB+OylxHsuaxPA1/cVVHTL+1qXdtaol45t
FJytwtMyJqR/PMvtNpmwI6VL65jhu9nbCtwyjyiFSzYAmaZN/fTOZPG3Rwb0/lP0THcH8BvDtj6I
tLPaMFXaBKmg9t4r/XHCGDJBkC/G/0Fsm2ggVB3Uttxi/jGyoN5Ld+Yo1mUwfPASvazvpYNi74SY
FUOiBnekwgO7IcmBNn6lNLGDHP+wTtwVgsUlK8Yw3sfTD6BVpLejoOfAByH4JBP6jUzveNoDGGBo
pKgdbdKQg3EReW1/Oe7dVYbB5J120WEr7N/X1Yc2haYirIvM+b8ETqz8wDmPsTq1LsMKiAxg3K0g
O3cwJCzXTdxSoJssHNl9D5kFKlWFYzA2nbIXU0kTHaE1+G7WXe1ucwPP4ZvV5yocakz2RWx6OoK5
EEf4S/T++O+bGxRfqkSlNCz4jSAkAx4bhRPua3wfoEwuWPELm3XIar/g9v+mk+Ny1gqOGiRUiBgL
kwtE/Mpbk4BxGHONyBgShGpfiVoL0bKdgQpVDgsyWk2N36N3CmYvaxZpU8T5nrlsnGgYMVztr5qw
QNoU4cYsH2EoQckVPGZiiPcgq2+Oq4O1X16U6v303w2ONC5H7SKpcTORRjKwtXRRB88/JjpU8eyH
ct7t9/MVbpshF5ekuZKNEaq1DfzxWeYUmsv0omaGjrhAYyyX05Z+f+cJtgB4IyD37bgwXlTM35H4
COcap7+g6rFuCbsbk3T5HTPWBTDmIp/qIoXgFBg7psonuWkyWAwqaJEWNz3Q2hGhIJD4d9Nqq2+a
LW3T2hSbTPDsLPQbRg2C2v/weLIfiu7QBpcB4WWCUhSmegf0/wjqdMUoa0YlYxKB0t4AsepIRWJC
PpTp4I/cqVLY3MeCRhNcilXJxHA2N5DsFiL0B/+9RtwAOzmAGiQOrt6j8CEnh+uezxihPOoWYp9+
elVOh5tBNxH6u/FuVyYNA8BuzqAnB7KZwUEfThLkD5Dh4MDozhj+yGRKdGvNppRcRDTHeGWSmXxB
s0lcaxLuUiDOF0w4lFoAaqGQe5CtaYYpmWV49Ivj8ZegMURZynf/VJHIMH1fXkO9X6fT4UHmcGxO
AvXBPcE0nwW8QWeqdMBgfsykFaXdw+zpJC0WqS8zGrz321bhM3VpmiSabq9J8b3UOAQze6PSevfT
IjRj6T6klkDmTdjwmHednrWaX9nVo3XuPd9mJRLd8KQwtK/2UETXAr+fX0c9lyO8ofSeaWpAjs0R
CJU+oGD5LkywNak1o7xtHW6J+0W22Yg6ftI2Twgj/1qhdZ74GdpD0FYj5IoI+15xu2OFIXkdgMfz
FhxQHckvHdrgKiyrwlqh4MdYArk6YVN3sfV4+W0D9XoIgtRcUcWEcg/x8lwCcI5eXDaBhScv+REB
V8t4rCQQRCTy1A29PRk4UsRccRtM1ZtwsjG7b4L/AqsIAI1SuhIB3WzeP3nlz38yTyTc5udWesaH
x9t+4U3JxnEszAibF3Na2QsTTFBrfKTOV3qG8vPmcc1Rl9dg/2RdmOF/D7Pz2p7mLlnU3CfVxi5r
nzei6K9bc1pD8MrOf5FHgDs/4ZgFX0P/Or4uFx/KsSyBvnfWzRkkrtCLQxXOyI6UxrEep18iQh03
ENlGl+LmX1Sx++S9PGDm2j2PjlUbgwjdT/X+1NQ1dBI022HyUdUzkYulx8z9Z4SIinu2N5eIHC3p
aH9Y7Crdf07tNVfoH4KZCNls5PRdcGiSJMLrWVOWFwfZH8hMa0czjrUnQAUaxb4/D7yCRFR5tfGl
LKgw25+VL8JJlw5cTqyQl1ZR6hf8B7OzuZI7V9J8unKBNJA3Ib7z97UuZ2chw9k7LEOA6Qky3mDA
tUsoPLIfez+xDoRCm6SMF6lLkJenjba2KeoIHvKvsdslhaf4xQxOtIZORw1QfSvwZX3s6wQLo4C1
JFs3Ja3JGkj1rO3rwUpKCt3UsR13/4EEADCRkTxCILG+dvvanNkANL5m5QKQg7KJfaBpaB9t5X8k
Fmv29wHvzFU8cnkmbTt59Fm74u32jFnnyC7pc9kx1o/p5dmWM4nFLRd2b4EV4Yagw8QU4t++2qjT
hx2+Hc5XwO+vr1i/R4a2U6xyX/8RA3GIrrz8OR467j5FXGgnjj4W3tCsHeCBzpaaVsMEFQyRx7Gn
TTAa1i6PmhcXo7az63tG1SplOo+TAhAev6HB2iW/in8Sr778diFQYRUVXGZUJqVXWAIxcvg2iARn
IfPErO+SWrz0IVPGjSC/AwIkNHvT9Um8YDsylq98WHUCcfSjYSqrkUxtFO6HyVoEf2zldQAFr1kF
jPgNjEfELgiVo1l1U7iue0eYpw9maydDizkIp4G+oqDLlzr+O9wN1vehV8+MaX5C9nREJ0ZXObda
/TKyP9Q+UnFH6uuPZdGZe5MhU9i22mCJzsRzVDwtfdZ2NEinfs7HEpIyv2mRpq6z5M+4qSaSA2JK
I40ogbCz/9QOjSG5hBAZIV2piCsVFYbh2Zw2v0SiAbNUI8SuP4YkMph6FrbBZDOJH4Z5VXM/danX
YcbnwRxHF43nHdV8SfP5M/lSDMJYLW/huYcZPdYIEwl9w3KeXNukv685yJbH/MP5lVqRcwA6dEHT
rKH6iGqm9tmZKsnFhot6L/thcmXuPg0HpWf2b4Ffh1VltjHmAqzQi4KfpB5P5CVmJjY0YSl0xd6I
/rlVRNJAMmAjWuarVj7/9Gkxs/d7peW9JdVGNG1IVZ1EtxYnKwh/umuqiiwy5gseltVsnfbEo1wY
jTok00wsfVYAWA/KkoAMGT1NsJkwrxl47U9Ll4272Peca5l5QyT25qFIywZ0gg4Xxd0gszUUoTmA
31inAPE8T2p65ALYAzMWRvv9TRIcy7NpmgK9Y/CSIJbCISHzkKb2NLUxEg2hjiILoSD3w1tOz+o7
MH9jMp+sH//Tu/tOAV/RRG6z+pe9yDaAaPk3Y0Nn+TnVNLB+Y6jXwh4VXrBhnFS43hMo6i6xb8H6
tdzeN8RChlf4sW82U2LsM2WoA44gdj125oZlujTllRO16aAZ9eFeHiKRVH6BE7+DPKZpc3l1I8mu
0BK7RqOK0FTQgA2vaLHVqePGCppBRxseCGoUv4V6GCdwarNRKhLTnFVth0GbbbA5/tFmkVrsr8sK
YqeYZk59yZJOMPD+JsoKryhswjY9yZinN78lAljGF9KIVUowilP2gK6byjVuOTo1lpBL99M/zKUC
/HjIiSrCq220Dfh2/VnrOiILE+gutMk8GYsZKeVMCsxTwEc7szNLnSUGBMOc6WpbeFMsXKsXWfzF
lh4IFaTBE+NeXMJRlwFJi5mvyrbGeMX3QplM0Tfj7Tvq1FbM3GqCp3cejNxegKb8hqmxUvwRW4X2
O08yt+bp3t9TMP8/DFDNrwymdr33xlLGV17zo45lpcvq5H1OeqLYTZWsl0/avlvDOBO/EvkM+sz+
W4f5tDeJVS5b7J6fWziuj/YbbCXCZUWGJ4AqCCowWmDTaTJ5IrsHB1KnFXquu6Y66/CqeSUx5mxr
pcRmxIOW2XQYJOtGSWRAl5m3/mFOpgHzOyq7+iG0tmi+GX3QdihPdIROWYo9HWY7S6MPF1jCuMLb
5BAJME39p7cfs43EyQMh76B/MT7enF8LqjBmwF1qX2iQ41PiejXrOAFP9na3qsCXB5hfibte8qdP
FcY1TAqCh3gxrgeYDacmveNX+8VISkidp5nnrPCM9DttKJdkSRELcNf7/WqQ9dgMNF2uSSd0ZYjO
euxIsBBQ/8AHitQ3wEK+8Z7bjGhPW7UJyMMio7lllEIwHsjlu8iOHwPUhnGAbR1pxNYr1uQ50kkc
2E2aqwn83GZKC+JhQAaxunLZ8jemr07ymQemorPVRtycfPaZNOFcvjkpRD9ClP3WqVpWwbO3qy3k
vI39DmqMgBeG6lUWWPTa7a7qBPSF8+uWno62dMSlkP0DmICxfr1E5xmbuOUmiNwpYNGuDJOkCCSF
rn4yrmB9yWmXB++tI40fMFifQ7n2LP9u7WIY5c8m/eVt93Pefzczvdxdbz4QC+XsY5S2jnn4BdWe
tcilvcEtjfCwsYps+Am+kHyiCbLBbycdjlRyxsnrpwrZsXMfijtrqHmuSeMh5eMSMX9UrSPCBfah
SYgd3wBvikpwVNb4voFUEuuwYKaSOA15RbH+Jngr5iCQge9+hjEJ4BOu5GpJrj108VIwOTXTU0z8
rUpXZYINqbX4ef0SfUriyjBF9+5mcHCXeLzvCXbB95ru8x//PAjF2cJevOWSR9bM4/TqoL/suF5d
Q0b6wJAYFI8zeEJJqWI5K8bD6k0pAY9dXLYk72H9hitAGaQsy0n40IYaeoPmQxL2bFmUOuG4VvDp
DjGAQ3VHQ4w9IsFW4ddoEWWA8DPPMeqqajKvnqOXvOMTe86/oTLTQGxWgIzV/tnkMr1QDLz/uWN4
W8gor8OM2/b6zXUJN7wB6eFiooroa8KgujCowhd1j3yCHyip7m+4mMFIdOXdawy3otZY5M+qgkqC
CXaiIj6jSgDa8crM5aM3WMCif1dvjLEmKQN2NRBQ7qao3pkAykUN/g/fqYG7T0OcadNStJ8ql/uP
Z0Ru1b+eMjRjIw395dBYGbf9seSz1XJGkSUIAf63Kc+/F4k9gBXH58HZ5tUl3Xy9EAFykmB25V04
jWN1C2DUsyhfIistjJdPVcSgpdnWJbITQeBpJL3blDXf/GaK+8w8z9Mo1VsKGnnQO7bZgJmea0Nv
XdW3wOLCtrcdX4GmPBT+C0C2APm4ZT9vmaj+7R/8gJwe/YZLwQNDCIFAwpqCal6NuWI+9iLTFWLI
MKHg+ocaVu7fKjl9eV9wvZuzino2/uGulPY/c/z1lUUiHrVhargOYLY+nfgTirTbMC4E3e7yaxqk
YyVadSm/LOWaF1DdSY5i/JzqlWuIQ4mcov15SY73NDDbFErigqDpL9BwFGyRkgiPEt6wP+qmvdgO
33Rzt07S+LP5ubk1dHGOHJoUm+aii48xZco85doCMB6jCldZNfrMvPQ5GBlShIEMe6tvWDo3Ncdu
E8SnMt6GURECZh+owqBzb8Cdlkk7MR4uyEzSxITzs+7uo/wlg3HOgO3gLsT8nMIyMBv0+GWQ4gIG
f0WbvmbLvireP6UFn5VGIlRxMo296PhGtLbLgw/prBJLXUO66g1uzFo2awp6B0DcZsGW6oIRI3dx
uvqd5pRecNq8ggcbLQ6P4bPmXLhfHufUX2GSBTMzGY8RIdYdCJPyzpoxmqHeh4wv3xqfDLM7ATrP
9kCcCGH9nQJ92YjfsnUPbg2SCGDvIubXKzuVjtZSRdyEj/bLLKlIYQHbB0yp9puUZJkj0CCQ8HKr
nQ7tM/Hl2BcCm1xqwwLQd8Zot5449F80DNHlBYjIUSABEQ1RO2Y5i2QRB/4CTLMApb+4xlDMiDT2
jFDTOT3T6d1v/u2U6wg4jCx9tHIg9MmDO6GTv9Z5ll/wdILijxqwUUWwJKib8BJVVPnoxEEbicd/
l8WCT3YjZEY281/Awx/S7TZfblvEZeVh8XSrzbi8l73gTqk0jt4FA0VBNAMxnwTcg2kWIl/KLD8q
iR9CB3zm67GFZjz90XA2xjcr62xuZgXygaq5Yc+VNG5XS+FQk4+31QRmLBuueSWMvxpu5R4RMEUE
oPRKuFrf8OcHofzAx1PBC080guAJTbomS/LVah93o2h5UGdGP/QLI6G/z5uCBc7+yRUTNqwNS4t8
FD5FWFS924KcbieHe84zGGG3LBrSjdQjF6kHTmrY32eZdO8usdDuyIG3zqS3YyMIcuhmfzVtLid8
xGX/p2v6KW8FaFh+78jzvHNTZ37f6mIdaRn10htOndwcfpOjtzfOAmqCGh0hDp5NJEWAioCfW4zc
YQn8MSoY24CA7jgPcjk6XVzYVrUjuNTSKp8yEWDnMdKHWCV7ox7OGOeqNs/yW8gSgEJ1xMVoE7pL
XSbcgEGdFaJqY9AJ+NSATN+ID4gDpogAfi1/TY0Icj3q/RZVnU6phKoFo016aJYufXt7fDzU8tb5
iprL1PlnwkgZRjBbo2RMSc6w5AXKcQoC0ufguVYkF8va0zQgccUbFwTMLiTwJ51VLFOQf9Lfd5Sw
shA7eZewORP1wGIRDyNXpuQd/J+UWJxD56jV+RZaew/aNOVnm6WtUwhdXY6XuW51JR/4I5WOuI0t
C5U0/YGJGI4msHlpVk2gt5XW8YPFeE1GOR7SIdOndjWEr44I+jdOUyya/PH0hNEHK3fYDxSyRpMV
NdMa9Yvf42XiaoH3Ehc9URC7h0pU7q60/JHDDC8Qp6B6UpyAHAQczDKbdhBMjYP3j+tCjcAFlklL
7X1Nh893V90JswiWwcP6QD3+ZqnDIxv6d4I3lEuJXc/fsm5/QyBMRjFnuJMrHPc0NlIMz18cJ6Dk
V2UNWhlYFKFdynZEgXHdDuyVpurjqZgyyrEsKfw31u1Q0XZQPSoSs12NGGOT+Qm4c6Gx+gMnMKGn
pnbSDLkbjchrzO22h+gQ6DN0yEh1CA8Isi/fUCuEwnBuKxxI9Qst5e0qeCXPizz4rrasPQvlq6Vp
toOVg+/m2jP0/XT97FqUlO7ZeHoRFXofXgYj2+MvNHSdAhJiYYH4w3WIDSMveRxYSJzWQqGAxUN/
IB3z75Pxa8jqsD9V8kXwTXpx1S/wJ0ocxh2ZlBNdTdrix1pliP3p9U76cc1bHYyJecdN1/8ODhwc
c1cF+LUfZ78cq2heEoJP+IUdE0NLmhzmq3a8IwvnpzfZ8u0OFV5hmzWQoxAvvPMoOg0YM/lwhj0Y
rFN7/IETCe4YN8JDyrSm8N8dsrciLk2CSSwl5OTMCw8u0UBPU8sEednT13sfKKKmRztVH7bvwf4B
btz50TelcOM8Hnc6SYI+rUZynrZGz7C4dFMGLAfycNaQPb5BTtga7cbomi3jlUF6wqf5o86YJK5c
PaIIuROQlIU4DH78JFXMGQ/+LMKaaXHZoyGT/2qcjBc9KfBc3lvd8onyKWpCxzacRpI5UMNV54ij
8lSkq3Ot/ndeASsypYPy7hh9RLvvYxGNzD4a1vVtQLtejYp2x6K0I7Cwx/jWvfGhmg5bCSQGa7vD
6JaOhe8Sxb7K7nI+v4c2H2aaMX5L/liKJRfEowshPrkOaFeQ6NlrfJzBq7G2Ra+6MyA+/zYzjoUX
05Xam+/3mjbQrxskGZ7MzcQbY92McqbiK+sqiKP2Y8R+Q4cQbWrJNI5mHOQ9OZZ2831jukxZPHxS
QMV249SnOEu91E3dLuSHBcmO+1qceJmJVvYw9vuStpkDPHsE+Tm1AWgtFOUrO+QIFtfDqtA5lMPb
KV2V+9uss/mfsuQPEtITqbhsWktLkLha+EIVJisq8sKq+ppMg527R1Qv33xwUD7JxnzL7vYXRhYR
5bNtd86dKFONIWpHNWrhCoMuyEaTUtEEVQ/MlwokUT3ce81SWUPbovvPy2d2bx3x7PIGxNzUzsSF
oR9G4KHOh/+wxBBS8R8onsV9rhCW59AC6XzhCPCxk8gYLWYW57Z2qM28HNRwuwiiRrmQ4dQa22Bf
UGnTLM+uBQku7YZKx2eEkdw6bNNzbKI6daOgyUBAS3Xvlf6KAJssEmywm7f6Qn1n9C45AMOFSvhD
HTkzIj8uea5JuKDyZzh1F4v3zy10487vYV5pQN/W++41Hx9F+vP21fJUvLSk8o4bc4IoEUsxuSdH
gNgbodR0dSkZwhtj1BmfQu4sGuaNJAC/w/BK/CR+mgFpYfexuQ76affmCLrYaeZ8Gpg1z13rPlNX
RVluzsNA/N0tl2Rxbs4Tj+0o60eYyOcpr1+yQFD+5w34BoetfC6+/GxRRXm2Lz156n/s9L0Sd9YF
Vu3tNq/NH187Ki1ved2TTyJ9l4exzfRCB0EvsIuRZ8LgNCOB+AzWgH/PIcHcwOXZVxduvNCQvz1o
18FHEJpI/MLASir3KHXASKU+osYANns5ezaxLCw+/RQh0Y+f4B6E1wPeabUAnN2Zwa3coeRarJb/
m6ICL38QgmmGg4Fm7PpHMubbPCwziqxISHXWFGCH98CI9nIaRdA2B3jzZ+5M6Yn/Ntm4M6CI61kJ
uWs1tWRAteu9zUEyUy66AYDMspvkrpTHFA6C+BtAy8o8ELCdkN0T34jfDKsypPAk7cP/cd4hRX/U
mMmsAjML2zPQW2zyToPZXfEscLcnJB1zm/dQekvpEksltOngnOUZ1v99RnCNq9TlVYJ3vgiLzWAG
lAlkAt8yR3b06Vvd8Is+IIbePuVwxGjYGMuW6qFG/akS1gUeEzm1Vb/IwAa4478/vqHmodZGQ3Dk
SRIYpCxzmbihrHIr+2x2nFgzH0eopuUWVOg82tIBlMCgdtz+065uE/pWGqy5VDY6uOtAZKpOSFC3
LRRdMERi2lrr0N7/znv7H9KUAF4cAP9o5T/hKamP7XiaWddc1MhgchjOnksaD9IcdQh02YJZ+ME/
VPvi8m6hC3SJdNat7Ugs68DZl4Dwk5BJHXAp9Gj+yHqfh5F6mwB5kpoTkY28b99bvEZkogFiKGPO
jIlyLUcsKHBhQXY3U5KGQE6DxBiSfRohuXcIEQdeTqi95LpRi8ZrEAZz8KF/JldZmFoqeM435Suc
cpJQiYyU5q297B//Q9rTcip+g0o4BCNI1gX6GsAJg1/RL79WyRJp6y+2B0PGKQ7RfTQYsyTB0RGo
hsCYsMrSLM51/hk4LZALW7uWGjC+ix/z+NgoiI4BDKJa7ePdUwVMS53TFfgZniUOSUtUYjLrIYG/
L0vl5IIuV0D5iKwQQMpdMtVLrQrInQ52/Gwecsh4WOPrQkIXg5RsjCE8L36Qc/CiS2p2WYJ6HG1P
OppcAu44uK9QCXSvm8zClj0KV4MIAVpZSD8Zsc0jKwjYHRvrOFCqt4XM7TJrM8K+bfUGNYjXoKzd
maTlIRZIfG5OUWiJIVCEBOR+t18B7QcL/ajkljzfH2emH6GQOIBohrt51gLYESA4XCOsKdjIRWct
vCfAu3NgPZUFm/GQoxL3NPZVTlFqdpk1GT3YmWMGuoKXH3x9gDGUMK0nQPFqPTfV1ppMtKj3nlgK
7xxhXyc0jY7dD5supEUcL7su+dTYd43/fhoWkOQXqWwrlEa5Of4XZBnHAWW91gCzgWMBwwZzM0Xs
tcolIZnxz4Mid0KrShcn0QxPVC53tW5WN2CQsRZhzDjLDN81LAwhJ0YFPvxwM8zu78KDxzEFLVKJ
YtOh30EjRGRktJLpKwbTZaDO4kcPZCo+bvXbxqSKPSVTzsf7yG6jo9exlIueqvGNdVPAknwyYFKT
R6BWplHYAaMQ65IICjPP1KX03S7MzTQEhw+G7XUwpJDX3y8Num+INW/wFwixhG9l62FBrLGhI6ce
F61uES8k4PolIVIWqonIyco5vWN3mYY1znhGAQ/WWOnefnQxcY1imuwYtTuqMGiZMZAjoPT0/4b1
Iq5x9H6s71WepUXLrch2WjakSaRI0OWygUjGdiO528MEwuKYSqDUYlywv49wxAI3Q7cdeYWYwH9k
1VD1AKOdj/c3a+L52o09MbF5+4+DRVep/j2otqhF0kt7qvmzOGWgCPN1yPyoFdoC9rPcOh7vI2Y5
A1vSfo2tzTvJdOswnBVR9CetfhJHJKaYYmqhb5Asf6nbtebO1Ajs6SIAQAnZweshupzwP9dlyuIl
Qj/tQxAmFnglN6R9azMlq5lf9PmbbNN12QEAWQ+iglndr18WcnQyB/W/fqylg5juxrr6zlZgkiVe
agJqsk3ccKSRAVNaKv9NSZjGmdniONxyqSXPX6OqKzmG5PHHbLyRjTiPugK5ccBqUz4UyZ4KfeJi
G5cAI5jUxtoNhv/GqV0OhprCQglB9DF74od1kMrFTUN5w2rtKtWlxHChBe5JQuDsQXHCPIN6mEYg
GCYt4LAHzsnTj1Zmo/Uwp+/tXh/19Hye2sjdbgUA1JFMpwjhPSipnMcktmQ5kVc2qfQy8xOIOO9u
/3SY2tzd1iBID5Q3F216U7y3vnp8RuV/pf4Am9D0b54yubUfBvXI9DF2CKGWomseLBZaLl9aiu0G
tzGyam6PCcCsVvV3xreQkp8vJMkvVx5rw6PWmHUnsKLOyRmkw7Oky0TAHmRcZaYkVhiUIRA4BSwE
RgBR2PAVS3jAXqY77/ZGuBQKE88jZPxa1j67Q60vA9T10KA4LDCSW7GnGz3HT6qTHsouEnQ9rJMs
XIwwvlx9pa6iKLxPm0gJrzF5MIS4fUXr9eiqwKAmCD51T/uL8Hdxeq2CzXbgql7Mmw31PK9prHAX
+TwO3CoQ3spd2UtJ2lHfzBqnjo8gFhN3B/MrtrXt+CCmiJo8j6OrPWERPRxtl92L9Zh63hIWx1B1
s4dm/B84Jwb54ab/CFP+xmHVRquc3v3gLPNV8E3VQEbCXTI4wE1sMIpMdStdUNs98otmLI5M8KP5
78+kuwElzEdzwaEF6wqkpRcYcT1iOItsb42ysTTbFiPx/1XOxLhPxFwr3P7x8hlc/Bb5pBJRa1//
7IUuoGOMdbveKG2HFizvqBjZJmfVJRMu58awAoq66PuNbRjtY8diCuNoaFQZRWwXqNmTyOKTJrvL
fctXShC7+jLND2/mVB1qoBt8/McLobUrrCV+mPqHKCpXlrQguItcs315RlgPxcEaMIMFhHVO+sfM
kL5esVNzGZnN26u9tfpUcgiseLNLpZeXPHOwuLsQjZvtls1Nj+VYpzv7HHPPZTL6t2Co6PtqXN+6
K8svubiinokgwCw4Rza+mJnQcTy7VsCHN1k9Q0XyDE9Hdr5hbKKOdf2HQRqdyZgDcq1CgdkBG5+V
YEYkAK830lUFHNhCF0UJnCzAqYP2eVposByTr5dR7czsKF4z4Y60B5jK9KepwpgGho1P+yujY5mT
/6fSD8RZKD9p04qBp4XAEZs2QTtO0W/XvHHhBHGeVdxewgQaQ9AgmOylkJxqHjJjD60U6VbTKrYk
lqddCfmacaHVrEsW8mhrgGXYY6sTncPaAxiv9gS8/BaSRQ0oy6w49nXRUWaXBAxx7yis6qkLEB62
WV7DnBU84nJyg/ZYwFZSzGfh1p3Ja/YxX5CLrg9Xtj0OZbYLrJMD3Sq26Ez3OdYtIRox24u5qPFX
90tRArs0I+tJAf4w2GZ20i1Epdy0b1M16TaVznh3UDq3xyPC2bZASb9LT+L8oyvRVk7exzET0RHM
i7RJMi5Ycwxjx5d58W0qI6VD7RSLkLcHep8hk6hY6NzzYUYVKfEKiLBFDNScYfqFGDnfSqYEkigH
0t/o6pvhWgK+MvQMlcAIz+SykLUe0GZQLjvmV2/Nw2DBl0HSiguzmLyDfDrg6PH/YWgORHI8G55o
dQNpdiRNToU8Zm+FAEFuoD17UZmcLsRlUNk5UsVAGmnoWpc+qB0ISd+yiJ0U3Wqv4oAeVeFe1m1G
ZRhkoSPV46LsjW/dHjMwrpHnepvSr2G/aocbw+nHQMy9S2wM/iEaeHDfByjblZTh2DSIHQH1E2fy
5SR+z2POR88qcOSQYI2W9lumPM83t/ZWL12MUgcah0DZ3SrVACUhYST01j2/M6zOcNyy39g+vRjl
UK9O6icrPo7dHdvybzQEeUq7uKGx3b6zU07UhONxvOpkTm2PqOUlip8kXbBomMGce/b/a1NropVN
ourq0uI/1d8wE2CXgpWSKPLCQmu1K4h9VndK2aulHzRShhNvGZjSDO199gojxVmcP8ceaP27HrFw
mXlYoPtw5kskOQa9fQLA4EsdddBdiN97CoMCTMwXrrp5woe177KTyyNOUZxBb+ZKOkpUvgzqu6P9
LDreR4PXUhqw1wIRvtGPUNrI6u+5sigg/nY6XyBCgNRK8/TpNpuZuXceUVddJeFRAypVUD3LfIj9
FSsYXRQMsh/bZ35miU7xrOEcVuSc3EC4iX+/yzzmb7anAXk9V2cx2pB4sWfrsnSh9W/lgldTSWGd
iG32hfPfUjhFIuILmywMNVxYh+MK0tPmnoha86IlHH4jCEXbbt1Vr74y7FTTzZZ0G6KE61H7J0SO
z2iJcULrqRZms3I1YIvZ2L40FwRR8UyTI3l0eGjtcQxeOFDCaXtWgHpw/A+Su/3ilX4o2q04K1LE
vEED5aDRBP+SvTx+6n+lyhOz6VsiJmEdcrjwkR+/NLnYxaeXVfzgNl8rEVLe7EhkKc1cEZOOPi8i
RgwmV4BaHlWsZHOgnzUyPxG+Vfnrf3mzO2KmIwy+un7rfqIwkH2m6yVxmU8AHS+W65ZvgSWollCp
zwy3vByB6Fm2NIiiNOLeY/cuCeY2fenAp1rUYQZjEgWUWBKL9l3AZk5eSLaqOyU9cgPtkSnJU16w
v43KuQUqjPEbNurleUv8ESqECLoq2FZpGzfm2VJjpl72s+1AFe6dsekknq6jr7J5wHygWP5rSO1y
kSOYuVuTrjarXQMkbKWTry+LHdPxAERzTBmhIMXdxIozmgueAaPx70AvhOK/VFBP3SY5NcUWQLfZ
EX1GY9XR4ZdZm9NKsulvxr68P/z2gWGklTUuSpnT5A/n9rR3TbYXQQZupxRh8oGMKldIAdeGHS1y
32kux+w5SGICiFiqHLEb7gl+3tL/v25AGzFrv6bpqM3msWp+3gsEjnttLnGasnnZnYWuuBx/u9Bn
BRAVX+kmMIOrrmuOsQBDFwCAByVcJezUYDVLL6fMfJDsTQt3kekE2rlBzS6yXJgqxEcaFB4Ntzac
kdGJPqM2UVLKiV8+w3DzUf3FHOdixyGoIW9YLjd1vHJlX7FbupUIhzYc5pgtr62InqcYh6ecwd8U
W3RV7mskhrvjLv9D4oHQHCZwwnVoRnUIeJETOt5yJ/3UyUPywrhODIsfmIowyT6idcnAruc57Hnk
BVIwAmC7YshkXy4AhclND2R9F1rB4wqcOZpcQEPri8lb2aXuqoYuwh37TFnb8iGexfty0Ghq/I+M
lATZB2zdJVrTruutg7TaKI89YIZUbNVmJ9ZozO6deP0Kwb8APbzF81/ZSgBFkD689nvvifjlX3Xv
qGYvDEjQyjrqbUdL0MUT+t4fjqMiGlMYoWvYhj7/7t93A7dbSvdyM+9I601Vtcg6dUi3QX4CCcuR
OB98Y7ThGiQS++Mzu1kCDe1strdkizW/QHXMsBU8/cofxJTP1JPo/QSjnmuel6UcZdwLRsyU5ROA
BCODhO9SVb/YSm3uGphWxJvcNwGrFlSIevTVLgZuvSf31trubgP75roWPJRIjOuPLISB1Nq9F/TD
DHR9uY4hKbbuKe0LrMNH5SncWj09j8jCZWC9D5tE4jjQwvmATt3bswunS2ZNMmo0WGnzPcbVbqEl
rMPk2UqR9xgRQnjTVR6AXqCIENNh+2+otymd5LrOfIXd88vHyDgGPmaEv9R0R3+ebOiJePC24Vhg
qt+heh/A8hNLkJ0YlMUEvv0FtoJdSCxKa9T2C4MYlQupI2MlzrKtzeiRLtR6UxfUxKSzRatcHkiZ
z16tGApilu/CbVRci1KY8KVuj0OXd5vDnHFzuJCxqBeDr8Sp/YcVVIMCOVMtojrSPJdhFXxubCu4
lPwQFiJ7LtJauSU8oE2a6rWLlb0ZXWHt2sOEjZI5whVC3h9OIjtSCLk6sTFyu4iyX39re5ARD4qy
oEoQqqswh6ZcR68JtET4mQnBD08jpsTrQqqk5atoPe1rMC529HUkS3WPESc1Jh23AqP4nxzVSHHp
QbTwBJsw/7URpyADRkndjf9JcEXMWv+USBE0Zt9xNPuWCw3ZT4s+LpO8mIoN/w6rW7CzhJs7AgUg
1AVwFN7J40tHtWATFIGnMxO3bJX1gksz+R7Z8kGQX/mf5bV/7RJL0szcBXDhwn/RJBQXimXLxBNs
BX0bc2kYF93MqkFvvjPIKUv5XYZ3DWQDF85DKL8nRrHnQQJXzSP5tej5EN+W/fzmZfm6f81xgVt1
L1q3CUrYkJgbd/9Zsigb3Man1nIccSWN+tVHPVSnI5r6ZG0qW8KQsdiZjBf7fBmUVYvUwcRDbIdm
ksttO4R2yK4trwIXZhjj9L1H9YMYHWH6wl4sVJF6Xf9NqBsIyDFdhM9zjn0MmeTwlFKA3MC9AqoF
Aw1w7rnl6kXmNBiWa4KKv0hMysgDD28wj2sDKiFrL6MQvMfAFtheweHugWETzzhAxEEfIcJ5WHgz
HHqLJSAUfe2wLkl59QPtYjnJaHRnbYUJvV/21GmeiHWdjzCenQdMfmRQi4qanH7I/UmEfuapovwy
US4pKmXgRp78fa4LHWeCR1At3alnL4kmgP4JySicI9e5Mb3TZrQ/5OujzlAcCOk8dLSJejjaMdQy
9QQ10ryLAuKbpqZ2S61adCv1yoNq4xgd5JngbfNiACJbcwOFM5UCrYRY37ep+Pb2RdVomwT8jzLP
8yNgnKKsfEb03a5Ztge73hE7aM9rfzHywq+Y1lKTqA6GBZYRG669AYaWHQmBJIhWEu7ls5Fjxkge
y2sN5mWfsizQigFpxOVou7MN2eCH+FHLSYarLMhV6elCEc2ATB188ire9YdqKeG5x+flvtZRevo6
tU0cWw4ioWzgni1N/dOsjMStXMhZdgr7Gf4y3nqLugiYdL1qBHpHkiPjC9P0PbqQRIBP1pegVpqu
EmQpd8vnYKF0C/ol4tMDenlWQoLazkc/c/MGsL6HuuY2PaeS2p89avqCEzNj36swXqFBAxV2Ajkc
FAMF8vX5JNA7A8AfVz0AfJm61I5yovgI6urfppy7HWky3xdZzGhPWjO9ZtZAdp23Nob76BX4Adqw
yUMUJ8rsdbaSpjEJUH8bXjKRNsNb6un9HPiO/lUsEOJn19nNmIOFCUM7l0iZYByGT1zaUsHEwwnP
ok1yJcf8wjIqHdJ61HAsHJUPdjmBHj//SbXg4ajWmeqbueZTaNb3H7zX2mWKqrZ6hRg+SOKyVaOc
2MR9EOQQqGYf6cwvdNwCb3XGwDpCDeFhcKxZ5DjsOBXIxIvOJMepQ72MMypH/bWhsKoA3v4Axxwp
uhluXafZArJwX5Dy4dmSSDKPaa8+j45XsfRvN4Ek3ujC15qQGtpJd7Hpopj5XAMsdfhMpKm5nG6/
xyVHfA7tqIFnyt01LD3Azjrq5sqWQfizfSAn0c5x0d2hmFC5JDlTTr4TV8/6QpVH6XY3/f2rwc+k
5HQSluhx9cC8Al0obJ+WA0KVfPdCt1CnSwy30gICyxA1+KRr7ngFx/KnNQcvqhExgkYA5ey7IZHJ
DnCv91UENnTiGEW+1JSK+S6ggg8WDaOQV/nAMLezwCGUHJFEAOih/g/0bVuqyAG2D+Gt0FtmSh6w
8nRFeDKHsy69Eg5IpA1Glse+ps4gbQMSuN+RJau84ghmYboAJ+bvT7bVb3Q90gpUKyn2eEJj+5kp
YIgiZ2k2lVasCUb2C9GAwR8r1DKTFuHV5TJJgeBDZ9j94PimDRlnvvrm0d4KrksbnV0+SNwCx0Z3
AjJ3SSu5YxcGMhLeQztPzZtNPuKw/HSc27yb65KlJszFQMYyG/Uq10lZqFDbjrPzCOUqi4mMhMOH
OgLntK3uwVEVccQDsR+Tx+FDnZuO5jGzVhmJebZ3i5PpBkjRj/FdbcuvKM8xSr6okwFiZ3OHrfX3
Em4i4MGzlwjdYHGv+ktI1lOyVO0mL3Raf3bupP+16crYu+JVyGy9kacsLvaB0mTuCphk2jNxUTx7
zIG2cJQek5utasK0jzNXZPRQoDdoo54Jjp5k7BinAWYuAT0dis1sf/+sFeMHCeAI1lEsARpbiX3o
LDTwQtxMUGW/MCSxUHDywYwhzVa62eRSFYwRESuX8lMmJ3/z/E/W8MpHkC/+3QPLLZVWF/jgN3I5
Rpg/458SSouwhtADqaTpez+rGJga1UTq+K2l9PVZ65FfGj4b7VgsAR+yrfC6HflGriqwrB2mwhbu
VVqdL8ZwXFcAT/8OuFQBkWVG8/NMFxUKhhdNhQbNw+jctHe2lNbeEoAUxJIw9d08M8ZCy9wpYNRa
BFJMBT1QMjJN0DFU72OqZtYnCvt5dC2rXaRAd01Wy3bKGvKjV6nDHERWi8gGveKpuTWKv9XsRpLy
vBgbQvzeWsY8k8USRBKE72OcWqy/ycJfPl/2tzUUU2yVPMLbCj3xbmc31jQMCDQ11bd7a9wGly9f
mV5TWmG2imVPzq3pqpCtrq7eCmtlHK26kJpjvD0ZcOv3V90fPYYo87gZDoWK8JeGqobWM5h2tDMC
tGA5dalLsRiq5j1xFAxnFoQsgonvYmbOLh4rqJekKR+q07aYi3tHE6wwiCdcT+aPEM49Dcxe/GdP
4xuqRIQcSHP0bK7TxMBomFOEpSECONMgX0Fzb0UrsQ2lmVDMcoKkW/hVPpsY11Vx6EQpWBsZk6x7
JlV5Ral8guZZGlzsEm1f3u8X2d0aYANdBivlv2nYybLj1Lhd/Zh3U+xeQSiN2owmgfS+UO4aVkHC
YfqL8uqaFt/wLYjc01ZjbnInP6KaSf3QASy2jfwrJRoKhakkMlBfHepBeQtvtO7S2iNTj/LijX0g
m64piasPPgDPvTE0FXN4BsLdtLaCN7PJBGBzunTXPG4bs53ghdGV+EuyOxfLO3uS8o/2FCdlGQDl
dhMuYn4Cjc8iHgcdUq10Wv3a7/iBLQ0M2ZGOgM6hoHmDSNRh4QpLeFr65cLN8l+8CcXpfpGjLGh7
mWcz+oZfCnzkhSRufmBHLK58Xfp0EkSee/yTV02aBGgDPg2V4pGckRh/YUP8i21JeVersjEc6B+p
eEBiwGGxd1M8w2CWp2FXsji+/xK5LfTz8Q82JnUN1dfddWZlrr+2LJ6c7EhmLJ0hPCXZ4fDBmQa2
o0Wm7aBp5avDR+onpFFYZdmVKaoUAvsn9NoRo4u+GDGjQJgqN/y2NDHHyLlySR745a9NMzpNNFuF
aYUpo5k8EmB1IB085mXdERhIOzH2RqMupTGg6Cd5kZuvVylfwapyFW9anZxX/i0WGjiwMsW+nT4A
8ma4yYxo2QEebLQoD7VzJbLwqyV+v2cOu8jByiU24PB946yFDD7Is0KgBVH0I94BDrWpC4qFJ1HQ
PLc+DhFHJC/Htz73hq5QgDpI48nNS6k/amWOJgXvFjZPxLUMk3UqWu+O4s3a3I3IDif9j/We0Bq7
5pIFrwQVIHn7J2/7ix51a+LiRSPiJ6ABapTl93y6L2EENsfTsf4qKdgOPMQZBs3Fa4VdUm/T1/Zm
8ChNjXR6wCpVC4sKxqIR4RFpQ2iTN5lIfDGDLH87a5FH7XVQWdaOKGXb7Nxj9fp49bCdAA1WbqFj
7YW9FXC67rqd5t5F40T2JbEgV0o+bLkiqjttX1i/IelLIBKI1iupezpV/IqIuXYtXGoaCi27qaEn
SrOyuqVGqmv0rch+5jS5LPbxhPU7MELT3KN6+Tss57D4A75KjWP5p2LntMa4HtDpzWaZUW7Atz31
Oid4ireiDylxFa1c9KLNYPAz6kDMQKkrozaAJArKXYsrzAZGgaikQncyRp8s5f7nU/usYG2gk9Km
NfMCviZYWrSddlHeNvadD78TE4vLQJTOXz3elNk9K/JsDkCXmSK9bkh6W90xT0jJeXQwitI5hpYV
KKiAXvo2rZnvohJWAN5u8srBeK+VXJ0DPUYUIJsfuTkmRlJlmDog2/CB/GtMBK/JLC1SedUvRU81
TOfg4BDk6bQ3pf6KKiOmG1tkVcLwPpoYHk4fw9S7DXp/V0TdMb2yHDF2eLCnSXHhUz8L1UhdFmlp
eNePIbePvpW2yY9mP+Z7z6w+i7RvUREAXCDcDxX9J53oh6sRyRi9n1Sr2ZDrVoNLq41Up2ctaBJv
oqmtwwmERWQxQfq0hvw+udshzN/UjmXwEgPUCNbufgKPBCsKhxOPMbZwhHBYvyPHT3SkpL5MtuUp
RoXHiZyxABF8lhEYN1JnKUR/eyaETsrNrkJIjEAvO+tYZeMozkvLJN4XI4OkEdoFw/CoaSU13oLB
hFBO/J8G94PyxXpk/UmpvqUJYNEzXu88RWMCWirVMQlKfdPXnQGAXCf4TtyAeOxW2DcTYk7Cjtef
BOmVPEpCMEBJv2UAG955Gy/nd7tcABnEZFcRR58n34S+fxwwoA7Gg+MWkMUO+KhlpGcHAbOC20XU
faoAunEESOaIhqgiWsyl1DkPEm8F0/WYPQiBp0vA0/ByeI9b5LfxYdPi5iKE/8jcT62fGuOMDZGv
02yK4dXtcn2xSTGsNCG6JhyyltTWQbX/Y/nIf/Hi565Dd5ax4dvWb4Yf7jgROm7FKXvtr84t56eF
/j0ITx5wcmUO9xgPYKYdzIJG4mBWfQQTUjlOndF2670n4QrC6naFSIpwM1YQwJ17gqWFeVrur59e
RZ6AJSl8WKmAL/IAhF1sFIGQHsmY9aGVlXuuiywiHjKdxgFs/noTVia7dYbCe++ux8+NkeYK/6VE
B3GGQvHFfOP06FKavP7MRiQsrZ+/1TL4l13MnJTHxVjXYTuHzUSdujSZ3pPfBpLBLRKpf6gEreRM
fmpnpr0cNIdHxuqPN4xOMkJT3rcNfNJdfsuIBCPW/smKcKawAdf7ijUkcvrNQi116hv3n84eXwKr
6iHAKLm289zwJE7khjVpm91/5JpQxJlWZbBUh8bvfTBakoSCUAQZay64/DsjafagtSx64MA2jzPU
eqSDdPYG5gmd3Dx1uuxcBUdAS5Muf/YvSv77F5noTJ+EzfEMXjjE6WEG1WIRcU5QfFDIaqe+RDMd
xkpP4FAs2KS3SS0nzlXyEeMUGWYDJg1+7AuQ5s5BqFI0DvnkEYQPL7iiLj/C5ZcbfrJBtudOBYIX
ZWkJcfED9Tu4FDmQmmYCS6vMvgT3IkPU0PcUspjdEJR2ofpj13DBv2Yl/pNP/gAs+ss7LVNz6O8K
NEspBQjJPCXjbna2/RW/ezDGxbZonJi/V+dmnGnq3m6fX6tLRGS0CZNPFb7Jdjlpvm5RPgoI1eDi
ap7m18rL9azgDEavBJpaAT8GIXLKcIrHQCNf/sZBLF9TIyCQIclpUWDQlak+Nq8/NWAZeMSckkwD
8xu3YzeV2yrtrfWpMRIrXoZ9mxt2gRYGTVXjQ5UcWTdYTk5fW4F9Wiu7aDead2SGePfE56814fyH
oE3uCVpcZBSDmgW1wnJ6mwIk5CzEHomnAwdQz2ZpBqExwMsdmgCHUfXw4bgDMKdAOP5+KV/dopZa
BqtUF8o4LnGU2K/bBH19BnIKVFJ3rpEsNvR38PvkNh9un8ahgtu19p1Uq9Znbof6xQPrHjpp5GVq
KxtZ7s7Gwef8a0fwbuJq5rDbp8eGdqnlPQMQYYY0x7B53OJR0NxzzzkuG15qR09L3qNSE4vTt8Qw
X3LvMbxFjs1pm1v+AE0pnh8uEA45N9mc3oDEHGMmTf3VIrqq8oXFaM8O+bq+LRwHKN+YnlNcRxSt
PXaDUI6tQN2TcjrExZhYn93TpfnSiBIgHGjr6pO0by0QXiSPSBh2vWCF/pc8LQCrcaGOi6a/y2k7
9oA62CaP99th/RfMxQr1M5a5GOIH3WVcbjH1Wvh/ExoFo1zanBt3C1P5KWAntj6qKcIk4W4l65HH
feTgLCAhgRjubop1vqOCEerM9NiOW5KTAA0tpMjG7ja1IHHqDcYjYQ7+I+qnMwk27ZfWU9tYfJn6
V9CHx6Eo0ku6hJPYHXcOSw0ue5tTx9+eqU3FXt4t2/X6Xrl/yXsEMCeVV6cZH8FTotaz+GsKnd4h
JoXZ+yz4xS0m9112vDu855onXvvHjD7TG1VezCXtrjxJSL84O9EA+YzFeVYnt0iOD6s1Uqmzr8k0
ctoWNzHf7tcsk3f4uHFdtZNxjDSlskK2qJaFvgXdZEj8KvwrouTjGTDNieojMT4AMaVdDmsMlTiL
95Qku74O8cfD8DVqiVPMN/xhe/JvR5W3u/BPSLyoYcylEquolpzaelPit9WyxFaBLTgeXVXI05SS
ag9s6h9DInTnDocjyq6N2cWfkmLEvXh/o/QqscV189glnCHQBJw9KlguiHd2pneDB0ZhlupGS69Y
mLA7IolzvqT2WdFm23mBPx/zfo/KlfG0nI0soouCwh1cdkMpRArrDafR0d12PkHKJ0iaRgu597qd
ZDdt+9JiEOmWp8bDLThieMh+9zNudFnQ5dhdtwdvcSyWbuxSqQuUoE7n0pEoVhFlvWg+82KQTqJ7
IxRzityCii3g67h9+vmNgv6uWmRtfXsiyLiJ/6yd9HEChxCsN++kLqI5GmXU0dGBkoswXWPRurf7
d1Mv941fGeDFqQ3PeY/qN8F5fsrm5IPDJGimm7ic83e80ie8l64/jX+c++BQI+9sWJpthrL1gOir
aXwFI2Z27xopcbjL0F03Oze/EUTOc8fl7UcAtASHGFi6m538wIXRN1pV4X8QCSST+JW7DU6M3P2M
a0fECkK9OOzg/fnGhEHF74r40hcCrf+oeQd63fziNqE4Q1P+OpfnlCkpaje82ltO835mnuwFrWS/
hiBgK4dI+ip8YY3OtfaA+qygbv7H1nz7gTAXjdoU9kV2zJlI4T3OAh5jbCfetxsQNB5b25QbgFDu
zwaPBGEGEkkzEvOl1UXIj9u5wS/iyK04+IrmnffC9QEB7fue06+sh+I41H3HDCKLNlPgmNJ2FITs
2vBkIZ72jGqO3sZCaprCJZB6kq6TzknzkvjCL+4G/l5Qb8yHPuAbJZEVgkm2Mk6R3SfE1lqgvRCy
PMHyV7xLsKwpmpbrj9gIjn+Y9qLhbE1Jc3rlVLc1KEDcqr25DeFwhoDoMJdLvtLfYjR3w9K2gliD
NebNI9GrsDR/bM9jvX1DKzDMq8+W5KYlUQoAe278p3lErR81Wsr+7KBV2OG1DV3rDxxuIdOcXCJ/
IfxsU24Eow9oo9FcGlBXWbZJdvWnoz5/m5NHh/PGIgMLS5rSA0uuUG5nqraDdt8/nPNYzlr2ZwoF
2zQ0jiRe8KNXASiAKCJ3n6QFegJ5ZR/Kt3M3QGmgi1vEHBC6g6BJ4wdLO1lZBlJBvHKF38OzZp7V
52fW8i+wqDHS8O7FX4ZGTMnLZWbCzhkALo0TpuRBSC8HSH8KcSzoW6xrpOEI8RXW8XIrtuTQB/Vb
Y/sgHQ3qvM/RAYgaWm6egHoWy2nXPx6u/Np46Z7zyypf3G9+8tyvP0spUiEMVZs3cyV7zO752olC
lZl+h295sOsC03unOXZ585iaV8KlpUc256pCdfjGxUUgicYpYwCzDDS15LMuDSg1Yh3Kb7dal2oD
KjZsq5BhdRDcmlHp+Jft+5vMwkvzBHsWLOq70bhk0Dd7Jc1r2b3DtoRIvNedi8fwr2P/R5NEGGMo
XCw3jjci5Fv/NBz4WPWzRiTMcEtEsl8hZ+rgs4ATSBlI+2HKD++FdQqr3ZKcX9kdQhmZkD4DyGvE
bG7wtDgmPm6EJT58qyyulFaR5oVjhMkqo6sJ4v4Z8t+XmkDhixaXelk7bMUUNp8I6yi9g0mkRgGv
DTJiixh/mpPsdlRyD7RV5swAL7Vx5vcqHacrDbAQoDY8QQTvurmvg170UrCFtOXreyvYNQw3D7nK
AX6VyQC/EI6EaCa2N0JChuTrfRVkN/p9a1e5YbfKkNF3fO/CtfMYT/vn4jPADiQt+L7xuxFPPkID
8uOcjcDzziRbsMFIznKZMZJF3jmGhLbODmYkUcrBEpo8tloWweDShktMyheF/4VRZUpMiUjqVZhl
rr0hRcU1sJFdqhNzagN+j3IUxBVTHSJEVv0QeL4clCpMVElZll0UelxZjNz6K2p/oj8XnjYX5caj
LxtC/WlgRseZty64LaR/imQhirl2KzpHYvXX4dqwDS1SqwEHv35AJYLpfbkk+Y1hkUJ92f9ShkLT
ktoy5iLU3a9d6scnSTjvH7/oXeTSGRQeO7EX5WurGK6XmTkuvGY0Ry1ylKkzofpDziCzH9Y8Wh5s
LdMRZDrVsQLpXOoieAcLpGBy0kBp1k4VPN6xxJn5L5cVhgo6EcEZWzslK8p+DTEzyn45ukTMOsJb
cTS7I8VBZPmq0JA5KIaECD7Vt3rJHlISYFQqPHWnx/W2JipIjsxn88uQYQo9wsLMNVznggZjIXN5
Y/Ftrboc+N/DAXc65lAxqIPvy2JPaLcqAbJj7Y0qoE1lq+dERmeXBqTKKv204X63Eo3a0eDtH5IA
pwUtDsjPtAOU0CDfyD07aSWUZuIPPoxnbJAPh5nVjqwLiVt2y5zHoWq+k081SBBBDzA9gfoM/b8O
1gJRLYxjIisKrcAGPhktnRRf+bLL5K1Wa7MDVTuGr9T/rMs1ZzLnyjLAWdLK+W7zWqMFwrFkDEt9
jOI9K6z/GWFmPYrnJH3CbGJdO4RBHwT/Kuqw1iYIKIKc1N7HOEUcYr3nnlpgkJcGzBUy3hoKhSfv
Y8FqpTkZ9jC9CqncTj0+Xt2hdXG5DZTqsM4YRdndL3StemrKU5zJ9PcVStSd0D4WSf7X0vEMjIn2
vsktDqWquCVD3Cfwzld2ydIu+ZIF4HzWkI1OwEtd+xlFUwa+i1YCdP71KSxwHoMxQ/5NcLMn7l1g
JUIa4btyydQJjrFuPym6lAhQPJM+RJ4MR5J17T7PVSOKwCQNr90iba8fKtHJjyczRymK38AAdMWe
6JZ7bEm/FbD1Yh9gC570C8U+4/MS6vPj3HW2mhjGQYY1GNNzvVVOw1aTyW0d/z2EvxbjcNaNUvdB
FoBRhw4jlaUDMwU0Y7zQCIu1wWfobO008qPqofD5EeEtBu8ewa4Cqwn3v1SQaq1yGfodFUO+/YG3
mtljgURnnKw2mk+ZPpe6/T+mCb/uo0DWu6ocm/wGHF4pdBSH7vKFmSSPtAZxugFGrR6hKDBj1NSU
q58aN3sq1KHXJaGnnKe+sTEz6b8acbf4V/XX0QTvxBqaxYO+U2bLNxDkjDe0JTylA1DsjxrdLEZU
cNEpnhbNaNglJoYZzRXhhBLXrK5f3YZVuSEk5Gaaq5VCcrjb0j8qA7VKMUKb81uLhHZAuLVscWkS
Qbduvcf+0O9X31omiR1RPz3ByCn4Ni6bBsM/HPrXaJGe1ktQ7ftrAr+ihSOPDQ9rj32exnhQldoh
ozdYa3zdYPdPlnC7arJk97+JpvMXQR9VhH4UDCVki/As99E1RxUeMKvnzyfd512gRosYGRXSk3n1
xfuy/M127mCIBzhjikH6Cw3O+IceLMFyUAUylYw5fHF4Z13TaDgvmBWzGltLWRZScEwLEhLvYUyQ
VkNFURkp3EIBlbmuaV4f+72e9XqPh8UgLB2L6Euu1u+NY/+C6q2j4438W4ysIyD879E9R7jb8qAn
EXSKrfMXXi3lcTq2LD5P6AafYDJNInuwwCcOJ1IZJ0GHhcnrotM04UsGd4WG6UiUNNLsP6GFbyFt
1po60VdJIHB99YWS6ptKVM/xjZFBuCXfX89rjETgYsUz3eF9uE908NiVY2YLNMnNm+wPcSmc0BEU
3owkEg1RVgDOzme4kbl9KCX/miB1opCfHkJKElsV241cUpwzD4cpInRdxXiiWXnHWs06X6eYrTF1
VApcKGSU9jKRfP/azgqsPYCq03Ym7yaazfU5lvb0irqr408OOBoLhbLPjMMI/88aokovA2HhT8L5
cElzF5KNPZFSNa/ulPNM78zf10QShMnXjR8/M6dHJcMKNiQW9wZV+2dmbiYV8jspbwYE6ib3t6NE
bd3K/HiYuEYkAXlEqPPyupzXlv+hqrmj07mk/aTzLgZDAfAXFZDP7F1uuCtcKgaY2cb9MQGsVmSA
iyKYYY4ZgsaHoEVZzQCPffEG4H7My/BoZX/z4ft8KC9rvH9NW7ygBTLQ95Y5/TnVHeKdKDOSmriX
pxIHnulULNfDLYMRLDpVQwC4UoR3RFN3mCK++FzdM9NDLFn7+ZMUr9u6WASA14p0BCbafeWMES2c
IY0Mfh/MDW//8AcuHZ83agYHWOHuD8HhIVuEH9SGvPT1/lyFJkmN6f4irU1AKVinn/eExTFy1CcG
nkD3atpPeV7ggvw4OUOkbYb2RNTIO4m/YpC6aPLr2lf7XOazYSIbBvM+QY0A3eMGszJMzYks5R+a
hhI7znbYnV6G8CV1hda2vOOFt6JVndIzU05kK0RDjM8LFYRBL3syIbfp/VBNttI8GJSg6n49df4O
49pmPDUjmFr0LLRTymfPu6pLDFQrRF9QZc+R4QaLtsu+XOWpVd3m/G0VR4xXxhAHr/H8iYmTSa8H
IvjAk4fP3LQEvqe9dDNPQ4uQ9mTHf1AIwoGGB9CMcoWPpRr1W1FIjSvn3tj3V4jrSi8camY0psJw
86+LmPZZxlmSP7rQFjXFB78ABq5RiN9AJWNm9s8P7HD5013nJXL4nqp9H33ugV4vcaS46UxgC7zr
GQxGRJMEUg+ONNy8NLiFWFoxHwoWNyM/ERbqw0HN/MNO1JFX1ghMQYxBen2a9U20bBfs15XaDKxR
qq4m4v7TaQCCroMmLxBGRzjVLQgjgOCyDN7b1A/yEfaX8IRGggypUp535fNPmb0e3dIh1tKF0bjC
T8cYBrDd7lrKiNwMZpLBfPqGcrmR4tXI3FGQ55S9/SgRLw6eTaVAFIrHhtU8MjR+mS6bwXGRfKch
UfPBMOdLPo4IMiwePhAbzh0JnW5P8hxnclcfwbyaOGgmWYWRX2UXmVRSAXLgqf5Fg+uDzkQv4GzL
K5EMRWWmyH3RA2XY/WM2sw3XAb5Vxd+tTe9QB0S1Spf7i2EkYTYm8bjFt+UWyx/OZq3U/umuwKWQ
dqwuKOimcVP6y6Bw16NMqISqsT7xygkj8MU/T+Kyyy967POInNy8jN3+kiRNTG35vWqf69z7NI79
Y7S307NCsIiIXV2ocgtVpFFRyd17Q1mA1XPLuxH6onCY8El2+9QlVGNIl/RbcVR0aPbYLMIwtCWd
dJkeswsNUgw0JlAG+UmPiYJxlNhlHE2fWZ5L15BYNUOm83KEOg0z0fcuLAzBJYHny/lRoFaiDOcy
iiJ6voCICyQADePO2+8TRAXYYlmt3Me7JDG16+WSmZEDF9aMUN4f4G9P2nB81NBgW1otM0Zd5wX4
EtL20QK4jG3zrrcxg++sXTbtOz8H/Go06VrG5CI/0wuY4ZHfIBAieKXIyCAXXEMGbZwxu1Ps8TIf
3v1aHM+vU8nE/mKDS0QgjZY2RvGpvkXW/6Itqg7OvZ4rL7oSVKIoJNoJnm6QPz2EzRK6gWot40bZ
KeACej5/Lwcvtu/zPxwBAVUdaUgenMiWktPAUPvNiM5SBmOHvVOiHr/+/zn1EcOQvF+ka1t2CYYt
nq0s6zku+Cef1iTD54/EtGfkLLW215bpMQaeXdB8vVJciDY8vkEVb2PMoCHoc6YOiumsO5hk4VIW
W528A4b4fMD4W0s1gRDg6LQoQBicnsYP1FFesb3w0vpcv1FWCEgruhi5fvL5Z5lI4xJbx1XJ+sJQ
YxvEq9XV3SU8e1S3vhRFx4vwKawhyU2YFvyq3nMgPJwmHT3LWoq4BMYblEp3P08LkWnsobfkO3CJ
Y5K9wNQfpmQQOg+hyQm4m5Yxsn5o7wxpCT9yTHsawUbEbT1GRsf9NsdWFChAXPhtDNNuila0dusA
n9MJnDuiujZGcUXDqwvqOghG6w3ZbcSGDXDCH8UR8W1noL8mQ6Tp1dOTXc1bltuIfkPx2iOl7eCB
A3BTvP6j2hsoG53tf1xCddZ4hZWdIRfJhv09JSmgH7ziKMVcHYT96n+VxHbLSHEMzA5XzeHxDFU8
b9H1wlaBtCSN3VdwxuUFZoyMMIUklKh9pO6EKWLunCUJK8uVedmvZo6Ftp1REOHRhRFaTza4Y1tC
9WAxxO94kesVe613JFgLPR7kTd+C0qDcf3q6c1xsxI8XJFQWxstSMXBjWEfxjQbc+N+ruzNMhNKt
DswXh747LbFeZRCdUaha+nNeY6fQjh/An29EB301jxqUCfOV6hBrjFjy6nXgZCWSKvmfVDoM1IjQ
hzEwCQeEroqazso4GR2RjBP4Yn+R0fmXoyMV1IiNB3LiRI7u2nal7XBtqS8MtQ9n97X2rL5caPXS
ytfZQNYuqoCmI9i4jfHhU4MCgOR996DPUmnjRxEv/dIuK+A0yxEDLAVVM/HqzSB2kqND+NXxbWko
E52C5ToEI/zkKvjDX3LAlArIdCtFoYl095U7ykMMYe4V/FJUxcdivLj1CmDAZEVx4Ttm45Jfc3ow
qr66NzxjLkLdjPhpPGmSsVyVwMIsxcpXbVbZyfZBckcvzyfw+CVzGZqLn5tBe1SVZ26CTKGXtLL3
+inHpHj7f3OMmBzwPWzibpLIkMAlXdGO94OvToh3DuSAiB74asAKRndT5eSrbqb7/XsD6Y99gCTp
5kJC2A2qZD7Bw5mAVfOCciQNGhbKNKiV6amGD8MzTgx0DtckCf3quhWWVsrB+F85l4+yrivkjdZa
wYU2yp7wXZeMehOoYvToT/N4ZtBA/YFk6m2Xvg/bYlOfDORlZqLfAA0GOl3/vdV1GbJvj4vKZMIE
C9EnaE8A1sgyCdSsL8WNtRZE0YpU4vlgHa2vsZTZSXQuXGwKpNbLANkvim/n/SQXbiX17W3gcLv6
LC7K1M56HJQmfIXpDNqQv0J8iml5AIqan2Ux/TN/h+HZC6ST/Q3B0tVdhU7oZK2czLp7fy1uLfqR
Fl2m+1wVRL98NJu58T/zXBiux6R7rSz8s/l6+0udMg3J4dvBQIa95F6eYS5zeb3qYkDWLn/k9erk
PnBsDlyIsKUtFI3IprP2b7ksfAgadQFiVNQiDz3F1Pdrm8rOg9SLXq0Ny8bNRjf32Xs683eIJP0n
q+Dvh/NxNTPUSgrzx/vZpebTRC0kzx38z00InB0nSg4VV+katvWkHPBOd28lQqybOCfgBuYH1nD0
1QYOs06LLDjMOzf8y6BnobuBr5++zLfQ1GIV6rjziabNO7FJ7E7+giqFySZ3iGuZ1FFVISIOvqck
263tuVcJwwW+jpFkjeCRc4dlM0O6rx7yn2Q80xWIj9tFU1cbl/ZQvAX3idYrAig1yImOUmgIGrn5
+wpzgtyz9SVXyNqA8AQoyseL8Yuj7oot63hS3yLub8k9D4k2SdN+/8arRN27SOvyP3IoTmNnJDuE
YUFJmmm0ILF+COZHk/t2t+pzJeVPC1ZYNMW08iK27AOgOO7sxOMFYFUb8qcRNaa2KqWzbsoxQO9i
y8T4JPzcwm5WPmBN7/aezjivEgSG8DhqV+8JAIrTQkzpKgOyNIBPufzO6LXAwmIqnNFy87wMbxP/
dTxGw/YKUncbS/ag55MEiM4sV2V3InCZ8iYQwtN6dXaFT/3r0q4ub/9OzMDZHAxaEcilCkxcEXxp
xrkXPiVSoxUNJ95c0U6Kgo+o8xy5D6N6xsw/a7GCg0bSBvyAY7ecK6CW558A6O7uA3PcDrjTx6lU
mT/oat+oUwonuMq56HSggvi8LWcS8nv76gQfsTiYkT5w7WtxKN1FohfwP0umyV0EZnLS/3GAy0H8
qT7cM5PXuqr1um9s4h24YJ+mjUUF+WsSGt1ROwqxVoX9nLWfaTPuB9AYqh5PMonH53IaPKlcw8jf
Vx+GnGzB8yQLH6Pm9WunqNUh7az5FQWYp/CS3rm8YaI12eS5vFCbq/U3N3VHao3xSiGc4bnEXpRZ
DVhO7FGdyDReAE+Tf9w7rrKJ3OLAfJHjAMzxu9YMvlyheDwQqxjvuP6FHlJI5pzf/SaonK45pn5G
8uzPZiW0jw7OkotU0FsUctpQTInGgdtYdU0eDEKxmmdAgMII5on75ep/4DSFCTyjIGqzbnmKzwoP
MXts6/9dmdE88TLJ4VRiO4qP+hvEgtTIYUmHCn5ZEgJUIgyITSLyV1qWjTiEQ2puCLrUEdc4uakE
Wy7sGxAEPpz8djdLphEbNLumB3MzYG0VhbBtXbADSl4ieeDZ872RYgGqK4qpSmucJx/+inAyZ4+C
LtxUmDeFmGAMGiPMgfmDM3AfP9VBGZnOnvmOAsWhtGqqikbCnOSigEbg8r5E8ruMvMXYx+jUR5sB
XVvIScsZKC9ErNEA8kevNicwWkUs113y1q3w8wxlDr0S8pIgS4MhGPsn71d9pUZ6lVIQqIGMYlKk
2vEP/kjpTvILI6RV7JsRJ6Gah7aZFZbxo5lf0VghiaoXjXYfJpe+f4VDw9Q8t0RJVTHMdmmeeXYu
tf0znX/KBo3j8rRc/6ZCYGGcQUVZz42QgAvlLy3qbInuU6Oz5++KScCrR6mmjMZRnmMpwe/I8CIs
3Ql/WtzGWM6r1ZJYX07BWESw2vbThuUNkHeR6hPxm7amRGd2vSKNjVewq+RrQGHPPB0DItwKQHhT
wSzKhk/06+K+o5graJM9Ac2miZI1I40zCe3uC1TZKyfLruqMA38ocIzG8BXplxwwhHgQADhrgJZF
kL5higPBCSJvj9Q60FE3zbYVZU2WAmD6bhfiWDpW0jwyXbl/4V6voWONkiRH4dRN5b4pF2YaCsj7
AoUJ5/BzS78wIIbi5/ZHaUNNraYwOfKFEAlMfqzctAjHeqri0qdI8WxYngfxexMAk+koNecL/qAH
/wHRuOux8g8QsJFvwvKyPzYQGNPpCaKU/+fB2PpaQ7SZJNwJWOxnp5I94T3/7XhEH58pcUBWLyJr
L0CwywO1lnMCcw7gwBiMyBPn8VnfMxRaH7fugNgUXwbZtGGMmB5vewPdDR4SA1+hOlXMrIGqOykV
Gwibe15M7AEer0UpbsDP1h0OuU48KsbXZsDAkbucFC4AYReG20HwXqv6CP/fmXhxe0bDbbF0IggC
B2ffhUBQfiHeW8J7Onh1lJwMN4MgHLMRDZbrWv25rI9RnS4OopjW4kLhYWotWfG34ZvRtx4AHRVn
9JjQdMrRnDAIPthHad1CLec2aUVNy7MxZpDyoXmakcbdbdTNjC1GZNlYhcdvcRF3B811C8U6f0wk
ECmKalIPrieEDTWwsaTnqQJhpyea1KjhWmaSo/rluzVZzDzqJmx83cxtbwfRjHKfGN7DWRzoeQTR
5ZP/rl8HkPmTPsUftqvZL1uSWesjV6c8D2X8u8SqBiHSBbx1Npli3cS4+/XBZgtNMQ/JwRxs0sPX
V6lD6ubj+7gYCUx1X+cx/vHCdaRuD9CRmW7v+wAlwxSFHwmE83qyGXE2FSMNOtc6Nk4CGr7NX8qD
DgHPTD3tqrt8ZO/rACjpV1noToj4DKktMaANfMfWvEDpNt2O2JmOOceE74iiajbd8RKgkLaowpbX
BUj44ebuhpAtWCVuWPf3cGtuubn5joyLGoBxWXReCX2qW5MAH4grG5/CjaPRGtyx8Cm6oINhuX9e
gcnPXALiAEkwKC8ZCJH11v7Zdusb9gxEhJ4UD8sjS7pFCCJN2+OADt4S7mpmHYF393H8/UCGAzGI
BolO/KMZlWySinIq9i/FnUNWYCmIO44qOfHZVdPRjDlEu798JVd33jAjbpcHaqpGbIzVH+M0tgMx
OvpSMNJbj1L27i74jOfoPuojhZR41hNhgzl5DdnYpQhr70vV4Q78TH/5olzXyOO7g+JoMF0wBQoJ
9l+kK90Xmvz4Itk9gRvgvmTZ1rQ4piONB8tHJCgJuNnnDq+6SpG41fduT0poNs/co7cYlu1KClrq
bOELyjp6GIPt2H4ocG+cty+5darGtQhoInYyINpt8Tdbv38NQcLuM3Uog8WxT57/EQ2Mtcs4GKQ9
fzb04oKAYhhive6YQm7ZyjEKpwdIkLIoGRhNqWTIoyUu4yCpNokYszAT0MRsRQF11Si3Eve5B8C3
WpYx9HXMiYlvex1svuc+aOcRKjcqhn5zk5f3G8wehg4Sk7eSDTnAYcFqKzeERNxRdlhp4QzMtgL7
mPzd4jRcus0JnM+tjqQcR8oy5sDo75E4B0cvYb9WbvdeC89H83rs1urHL+dSjK3AswHxqt5adglF
CcpNrl8s8McxjoRhY2m0rQLPVVI5KfpQMt5zPTXyKnQXzkPOWaslCvz319QOsIFwYIXbuQgX615K
czqeX2nmpJnt8g2WgIdv5avGSY7/ZIXCvmBoKMkbCWlNK3i4Uc2GDY2NYKuhDCWR27MOFRNwQrPa
Px4UjriMEi6TnTT8qltrKdJeKxA2KfdrJjJ1gluAn9FMPPPaCEcNKYfI1/JMK1oUKIxFjGEMvCLV
ZRJFj8HnanPXdoOVyM6zqfLXoDGVyhoKmDKVrGGthsliIAWg4pMNOEqCWUlGizpRbahZq5on+8Ab
m1J7aSk7G65oFTU/2LHoRW6RwTKjgnFWKtucUt070bSx+dIFdbHg0sydoPEqkdsU4lu6e0ouSrIM
Z75rCfXA5/uJhDTqxah/F6IokjNDn6Y58EnFz0J4gAuTaRobNdQejbr6OGLNAmqQj7alrOedno2g
W70PUIQSAys86sHtFs4lNHdDfZN1wYcqUnPv0cx8l56Ai7mM8nX70rHCmRJVte2UDC3Yy+bKwYPt
eiViZhK3YiUo2XK3FHyDIPou5hYh12bJrfxDp6Pbww0FRUz/WwIWuWlhOJ1Y0hOlL4PwML6JVXH+
R08eCeqDkJW5p8lPwaKjfbuOA5lMWOFO7qDoAu/JTEVEVKNuVWN/WvZLm9/r0BVlI0TG6py6Hmkj
AjOMAyZX7JwD+ZhyVIq4FULeGqMpNla9NAywcschutFooWYg/b1uVwwhc5nl9vCX2w0olchFv0ex
CZ53Bhc5OQX9VSMLUszgxSfapnn4Y/U4Gxbo26LvKUyj1CtEd3uKpgAFiViGUjAc5kUgSlpSAO87
7B29KjzJNj1D/0832laMjyb5KZvm8UkCz79aL9fxt67or/OY2FVBItyUyGHUHeyeVv5mbUa/V5MD
TDhgYq9o2Uipodq/kGFDRLtw0TcuGwp7ou9yxfrF4IwbARPWn1RA2F36cPzSbIJjRnB4kT9Z1ZFJ
bhjhoL9BmAAsEKrkWWfw/4JR93AVtetG4EgKLjTzTFszc+CW2Ng1rKdVrz663xJXjR42GiXj0w+R
uSBeeYw+xg8nMifjxpvwIBf6v5gdih3egjD76lubZXkCAWPYJlp+8sd7RWz7ZmbS/+0xtXunBLfE
FDQ3hQqjBWEkQW6U9IK0fSJVUBJwT6YPb8Y/ZmknLIbUN3XzJXf3BMTmonXZE3Gn3eFchWhKkg7N
6868AtTGKQUagbGYmw8eew6i7BmQZ3DYwwQ/IKmG9Y5ixtLxyszMhJxIxNd5r3GQlrfwZ+GtyHuR
lyZgLleM8IlT2tnCmNhkK/83JV8l3soEfnOLZJzmT1vM8ezX188asniMOTKSIzxw9g15HqhkvECj
46YPu3JREtLrfhICqkoBuNgzR2TjzlCcnZCVm0jiZq5+qzb3cRq8CxIPO9wQBy9m8/sl4xH6yBe+
rbTaC8j2wtu4ihWDVBpIBni2SH1dyfTaM8SqQuBkgRdHsysYDHejBZB8+JxYhDrfGCFgZkay8U2U
MBWCvW9wEaaW/YPYJeNNv0GpYxccb0E+AiPs6zEoJBF59TNnsKS6k2Gw1fZxLAI8J2cLSvLoFQlk
SNRVNy+QITj8b+YNvkLKuo17MDDPd3k0eHQqCl0yuvKl4rl+AJoPLwVSElWbgtWuBU8NLYHzhk6t
GKTq1eFd3+073SpcibdBo6sMPFJty2OzmZ2kazNHaMcYWKmiEkqGvyMUXJFelSzSxHZNzrbH41jW
VzKmKqm4tlhbJh8QbMURBlvoQfIEvs/u/trt2Pjbmau/yislmfdu3CM5uWPsz4Ui3s5qDjuwsjZ5
J5sFyBDxX9+ljGUR3hct2/VWs6K8amY4dXjnbR5aGv17t2vroly99edcK13dee5eILx1bjKdODxi
ApfmRy3ytUdPbKL9xn0I/yYBxRQHGEwuXK/zQHNQkzc1VDg+KtigpVHMnyrEqn2YNIm1Fd09Dk1F
nkWOa2rmzSHCEK/vI0NFq3pf9cgXEp1tD1Mq7FwCsx1eFjvOUN8DastHy//LhgCBt5UBRUyBly2B
O+CSotQCvSF0gG9kdft/re8T17vlV7XpR21VHD4hnuFl2X1Fzwp4tW58mn6Vrf5BafhiuPijMWAX
7nBYx9/p8LBbko+ODYrwYUMoBcJpRpzoY71ZMFQDX8jRsX7UM4lLNOVKkF2DXfWi3lt4TwE93+fo
LGJFCHIZdi4nuPU3mam88w9T2sf+gjMSei9Lg7AEhQ483Z3SLjFDGkxtAeV9eX3h7Vna4xlxcysh
hupNtGxhTP33cANM7pPsgJh0zaUQv28V27kY3X7zNsHWln3dvI4kf4c3vMTbHdNLugJW08evYOmU
KFGfPfaOm+T9VXtCDaF6MmG59kIul450DxBcLlAmQbEG5dU9QJ/KlrG4icz8faUBhsqahapvsrVi
COdUChActlPSatFCPkonS1iNKj8Mq6nbkLufzL37qjRdJlZTGP4F8cmpLuj3bcr3pKLnaB1aKE5w
1Fg5Y0/5/M5FWImB9aZHUw8vDZoTpl2qBgndH0JUS5exQqYhaDxnkXjF7ala4BK6hhh1jVcm7bU8
ARR/lrRvx9+ROCnsu9O0PLzTGXZIP3oxSUVXCfnT4femMjl7SmrYNMeWt0/KjD3ngB/+rh9z/9zU
AYqRPzKF3nYUJ9COnH9BBwBNRYK3kCCL5v/cRu1pRjdyOFa8g4LI1hnaz6e6fT/GBYfCIJNL5H0E
yYtUIRAmbZbKQSYUjGQ++RZoFfMCipzdbSrDoIZUNigUEvpvrKcwdIiS5l/SJ7aBcy/rs49XL/jE
agl+NtkVJZZdCQ6jZtwELi+zWQ7rxRY9jgCbo7Xay2lgRi0SuwksuypsrKBurTJbR2SPoh16tcHH
Gf8QpLCoHipFUebjbHdDfzQToLFZNPUTX+tFHjWpcDw9KKaTY2NfNtkJ0t0jqzmp81+m7oVTgqTt
w57TfDEmO0EulzST9EY9EtlqsrXiDjZn2BReiXaqkVL7j/3CLVKRT5Jq/RKwl7KaW21rte4Fe4LT
PG0x3BAVo97Ou4frEGvtzp5lyaXlEEhRILq+25X7/Pp+ihvG2GxFHiIemqa1XPUsCYG3VZ0EuvXq
TRxhrpj9IkCWeM58I1YPcFO4ZFS88QZf3NZQLToWbeoTPr93vTWOcYoIx25PAbft4rkFi3zgU3Ql
k0acLdpUOkfoqi75mieYR4TVZTdyvzRl9H3r4mZYQOXeMhBqXghAj8uz6go4fdvtGYVgOYlKwIEY
J3JZCBz9RHzmDAZxUZvKWal264hTds1iJnqgiTRH4qlQ414qMGfioeNt97dhqw7CideRSslVqS3w
myURdnVTu7P7dGlM0Ehbl607pXrxxlPut9ALRfIqD13HjdfKQkpm6345Ml4Ql+rbEAacBAnXt42Y
gd+i5+rXS76+zsWbIsJX8oOW9n877nuSn3O9PZych1mAcEGDcXLuWD+hv2I/KFADQT2r5XN7GogL
0v8vQ/LQdGit6zGyJzMhtH6jIqx69qJNs/bQgOR2e5B7yvOjjmaQXItPEhQHsX8+3Xpc8w2lkrx4
u7RPd70iZXcjhvz8BHQPdEzSmKpKK95a4w/LXY1/XuGOX24zpX9W61LDinNCIl28pO2weUAr0Cj3
UcgUPmtEQdnz9sp/DiuDaov/XFRHCIbiczjdhnHbril59YHYDET4cAj/KrRfOMwTeAjFa6ebp5kn
80bPkggMYqI+Xz5E7Qc4Ns9QVbFoUH7hHfMnzYZoPUcnHBua8T+/sb77Cz2WerRHQ8oo+DN63e61
GiX5qRT3muFiInmgCkVNbVX+8fCG7XMvJxy7YQ7LnpfofyT9Q+ZCFUdCKDqXJ0EFn/28tZftVkyj
CM5iZQS7TxjCS3pSwtA3K1W2frs5tD6A6P9Qi0DkUbjQMzQX91mTKxt0+41yd3SGM887L5ZX1FSL
0BFeDZkiIQwosN+TqUx75KP+irWb2JUDYYcz54cOnnsDT1sX1kLfmS8IuM3UIQJAgvbdKSoIxf+U
GW0NCu0Bn+/+bL/aWbvJiCDKvZumYRqi8vN0vZkhp1n71/MnHIBLCDRboQZW9V7Mt6ufIEIG9xul
H3+ItxkX2H0a4J+X3Y9zwiH4z2j5NdN0l/6DR7oq84iraDQ6sSMM5BpsXBc0EVBa7TpcLAV6c34x
t8wE+NLZsOXmyOKfch9pZAfSkBBlJgKU5Tjrr6zCxV5pdWP4YguHSHE2lFr0VvqbtZzRuF5sY0LN
ZDOXngN7E/EFeAZ/bOad5PqvurN0ToEpXjhipzy5pAbFeSyNrI81F7NQqsR8HkBozLUlD+mt8vy0
vVybzQ0xwyFDmddkFvjvlLXxyFcve+3gU2AgddFrD8AIvhBRZ851KnvXvCnuUnn2t2SqNv4H1zeo
MWmuaIT6/bK6AF0jDT+I7PdyY+3eCcjE8shbs4/aRRZABqRWNZoG7iXhMLEgLHTOyv9hduH1uVQ0
fXhLFhF7/+XGMGyG9ZGGk1RSwKb5up2Sv7iSHLqDAzmvYN3il/eYbLBemjZbajTvjyEMvjdCJD86
VydmVK9XhkpJgLfY/7waOZ4FMc4HkIZMSmEduLMw2lQkPw66gKB7757ZGXrQNw945FyWz5Lwd06g
xoGtKSUE/Kf2qEqJ3XConhdMqdrm1XHjZXF/qVnH7gguWMJx4ioqx6TcC7uvnnKgMBhvwOzjTJS1
Iqxg1oZe2f5q98BwWSR53uiCokCRXs6JjLB+QFUCIkvxcFfjp45VSJQgaQPrwpKQ9NR0Y7Vtq2RK
xMUG08WRtV5JFyUrp0iMTEgQ0F2B2aREcSn1NcdCBnhFjrBB84YQvKKOWtz4iN9ld5wNLoXr2xSz
MIndUXJ0CpEZ0xyaVzmOII4L7eFpBQtevdqPOAjsN/1/UK4KsyArRAbQfimd2DKceZsIRwAubvSH
+lr88rQZG2vFw2SzP3UU1nxisiFCzwnU0Le9BJ+5bCf4gKYcBxErXtkeKX/kFQ+HmDfBhZU4Xitz
17CGQkiInvuXJcyv4k/+D/bSk5iMOi/SW69ivyUFsUudL3829I8V3vFxfZeNwGmEs1Un6jVd35uf
FXjqhGuvOsRAKr6uEH/Y6Wm+BpAQJhzFOwVivUKat4Lt4bAOtZa/VrJ2EO8rRUO0WNBHdC4w7Bxj
LSx8eXuFLXWpXdBry9legV3kE1TnuEhJuRGMf5v0NH2k6+Hn0l30qZRmb+Ey3yEpqyCCzqNEEh7X
eQ9xxeDTDxUOtTRkeqgcgdPQSm430TVzg8rb0J4CYPm8E09+KZKI+xQ1XTuOWleGmiXTvW0gpRDM
pJid63kOjPED8fwK+IFkvc7PX+pj+lM9/slB7IL+f8Xadww52C1sBj6hyWRCE/9J500CkjVxI0Y4
TC4mHKGq7LzPKQzGNK2ug2R/KfuwvL4l4EKueHWWX7HSWNdN4+EZIsAUARcyZTK/FFrxPLw2sRqa
JLaJf6swAF5PJZ2l9koCFWnKUiVGnVkCY+M3JgazzChqISyn4UpMA3AWb0gBx5fjV1DeS7A5HB0E
3urOoHYmtOmz7zdeLl10VLrHHrUeEsQC+dX+MaL+KLYXQdKB0OoyFMTSezMcB7rB/M6wRIGWUbEi
zKqIXkxq/WFHqKGthdFXSLFqjH96MnXSre3tQtqGw1AZ62bWqHs6kpVpPvGtE0otyIPrFA1SeL09
tN+wMoUWl+dmbfwCEv7sb/IIv9lumF6eY9BfGqN7I6Cl2to7CH1M6+R3uExLy44EaUHMxfMF8HRG
3PqElq5SMptQkt6h51mm7QcLkfCZxKpgxWgeP5sWcIu7cZb7Hx2H7kl+hpyumpNpjbh7UNogN/I+
wkiufRT7LihJHi8iuHnlvb/oRmAS/maRimPsQnP6aQN4KmhF7hfLqXN44I66XV0X1uWILg2Jaa8F
TlC6RK0WL4NvhLQfnmSrG5lL08/ta0B1a98W7oVcKTB+kQSPW7LQ9cSphgdHUjhGk9HKnL4izUnb
0yrB+/AH8OV/oRSRO8aeyf5DFrUGKsflXJmharBIPS7QkfsK/489wJza2DzIdhHfXtQJUBWp0ill
kmkZwcNerYt8BuYedte8ZRKjIflB/e9Bu8gdL4V4y19KG3K6wiMK8ilOyrNfa0YYkCLBgcyS7OMF
ifPyuL4Npi+spdWYw9uYt/718DQzwEGuiPYmBEkiSAXizvlmqDXwXKJj21BAY5KUBfn/eSHs5W8f
OSMn2X5SC0OnUHMRFiARvmuCTOj9gkSTs5EgKBM2Jb+1CzROV/TF9+t7SnOC5R0r63mSzf4dayWB
3MqX7OQYtt2dM+MrvowXQzSmcCNGsjqXJ8QBtkOmtJ+SAT3KUe49RCyLl3QIgHYlm6pLqhmFKQ2p
uJ/LFF10QNQnDamQ7xAxHVK11jK8roUfwytMoFfdXv0nWvX4M0sSxNTBvmZr8y/0Al7ptJ64GN05
M6zEaF7pwE+v7IHMeYFBXLNDijFsI3/ZDKNTyhGxZYwVAnT/aBBtn0MTCl+vfuH6OTKYqsrXgc5g
XZ/Br87SatsoZOrjaY87HiyYTGbb337KXsVFwsPUG2dWXaDb/Nac5fuYPdMO/HBZJA7HEPqT5Rx0
yhAxyAwVSw6YmNHYA/M6jWTVVnX0Cc7hjzVWiokIZ3vzDFTNx+qwqJf3NmklEYndq8cDWCr0lgpw
Wdr+rxQlyNNOzGc0j2xdiOTq+8pIRNUSPmMqYCvMiFyiECIzx4hRJN0Qm06gsrOP80EsTYRsYOS3
dZ6HWwiRRYBsyPnz22TN1tPP0tDjKHFppHdAFp3pkhMf9zKP5GWwjYZ2bMjWTQmfmzv7LbWhTLC0
NJ/6pChmDRpwWLZGq4MSUDY5N6yq0Rh9LQJ7pIuriTnvpjko1g7SpPHwzX7AQmeBNY2bzNDl03Gn
bQldLmvMc7/pRh5ctcQPAGFyajdf2Xmg1gKLv3Swu1eYe94UCRgl94xxq1+GGNxwOVYsNz3SHoy9
szbbagJ7t8QUqhTBKjQBlS7IXrorrswQFspsN0lC4e1F0e5shTEiL37E4SNg5lM9sVacUbbLr9pT
prv4eczGS170q2OrcNlNP1WFzeapSk+xu7PdIDZ20whGMikdXno556v3B9rFXzntSoEndOE+8cuY
TFMYe83XM914XKYYFW7DKFBqun96SJvyV4hqRlYkBUrbnDJ3KZ6uGhLxXgEV3QVaNwYbS7A+D8q0
Wu//iSmXoWJcfAL618HsyI3XOB355yDuKZm9LDyU5XZVhzJK8i6cTG/2lZ9QOr7+mG88NhpU6Sqz
rBNaE/RuBlkSvw7LRyj1PjHEVJ9rlXv78XRHNo9+MWmdL5R4n7XBvQHVGnWytM12XmdDrDF5AhD7
0GRQIPqAMSBfOfCodZxPWbeKYt+1HCJeC5UcfRXzsuSITPi1q1vx5/9lI12XLpNOjZryaCA903HJ
9bqyPoZqVfX/6mN1DfrrS0v6jax1/1J22tz9TSsuto92s+4yXUD2Mz4AkFCip/88u7txo4ha0HDy
r+N/gmFze7Y2awhOzfq0w5FaQ4f3W6fSMYxeBuvQZs3QJNmzcDKvNVsG2xnyw1vld5SLpOGTruRe
VBOuRVrSz4z1mYkoCSBYP+6r1yBt6UAYK5gOkD6P3hMAdUpkmu1j6TzFWTFNu8ZBDlINiFXt6THl
NZI1vcbTOPk+qAkq5MkvPH2kfXo3ltoTWxRdtc2ccgDEajFBhfRPdeXRMF4XJGEvp9b1VnD55Ox/
FvoPyJenaExxKPPcp6I1nPtb0shaQcIUTPDboCFmHZrsYdZiuAgYddZLh9r5n73h7libDbcr5Kt0
C9VCOh6ZgHhfMi0/6fvzOkvxwbeT8YyuslBqiUMqDT1IDKOUL6LmDQqCpCXNP+R+0sHweWH9/sRY
br/tYvZ/ePYEsoKnxVrTizYZuSGL5zD2TDHEGr5ya+h2s15baNzMTWxk/5ZtMiamWfkgDSzETKl6
uaUNeTxG/ejxdZe2Uer/7tQDEiNoTmtH4R+li2PV2q4s2pUi+9Llom5TURIA8b++0Vn1Ll78yphx
58iobu+0BVqSmmSJwbxDJUXEO1aYJDZudqG+8ymGyGemykSV9D83Egdfhqx0js6qenN9tTzdjUtR
ADMNkTTm61PDzeZJZscwIg3KVQdhNmDvUtYYJU0jWbE/NP4KXD3WCijZBnjWJIL14lX8nJUUiC3Z
YbmVTcF+j107A7BbaoSD+bhDCDQuXR+xbD8up8TS4aKlDlD+V4bVmVMq/Rup9AGNRPb9LlFG0qua
xH9HDAQMX1IZEijfJuufEJtZuxG5WvIIqwFBkMLLqk3RZzxhkI/aIab0uD3VzPxcR+Z61Qfk40If
uAilW9uja94SRSQvJO8fjpDpbtiw63mLga8EzxmA1cqZcDxi7cljQg3DcmqCqFYWqNOgBAhMeSu8
fefvxAgbPY1ke7SN9YvM4WUjZZ17dzSCjf0JJLAhPQXgmQaWIcw0SZrmTjNKTTlp/7XOBkohRZy2
CVAMCL4oxE6Il/bqO4oAmlYp7uqDl64iwNFXE5Zad2wWWvn531cvfNuNa0bXOzNpZTYw64YeVgjh
CRfLsSxOF5DKLfJvhnvWbA0VYCp6m2j9OcLriCfFmF3wNEQCDYoaLLCa4yt2Ofkl3JMD2eoSDxw5
CbspbYH8eXvuxS/xrXifLh9MljOMGVdIzNv8y0f3ByIQNFRKanAnTsJg4sXTkBe1AMrleBntGN9S
CCIAYrSNB2ES3zhYHkgPpjFz4uIPpIEv+Kpl9a/E51R7J+vA0MeXDVNcQ6i/khN4IEoS7hMAUfKt
mtk+oK7v+LB0Bf/8LY+Bu3PVXF640KkBXtfWAvDjwSsucDRqkEoG9874fhMIeRCilipVYa2bGu3M
RnabxaSLJoqmI2JqbPueNHLH4GRAFsIZdw39WfD8mD1O1AVDxhYCnWaIGTftWU59nKivdmPhGKji
90MyPbDhpeUB8IvSW+W/7lkJy69SqcSQ2ZnvAzynHY0ft2AITq8IQOt2a0eCof+iGMuuHLBo7MNn
oW2c0QUc0mmvZuMBqSnMVT5388OT29Z4yQVPq+o4RpB5tj5zjuozHHucVTxUGU9O/rRCAbrjfoLk
kv/9SFRW3G18FzvK1AJasJesiq2zww8RTwzzfRfUfBdBQ5NXDQIF599d87mzYZgK7mDPNM42SfP4
CxVdJbY9I1tmNRpfftJCLkz83rFtfOHMllTNrZg5LxG/mkJhTR8Gh45RS661PqePM4X77GjC38i1
A0SoD1IzhJE30iAx4gzW1TriRGLo6vSpJ3q6DjtijJZaNPOFcVz7Vg+sOkMMUl2EeCoiByHhbHCA
ZndGIACkYDcNEUC3cIP4In6SJklgO7OJMqA/krGmptA/2B37EMVgjD8F5F1FO/6sOiKz0pYi6IzY
VxUGte8vYiGY29I6NvhDSt0ubzdtnY0vjin3Urh2XfuyFsNYV/mLRG8BLwursxUyB3Al8VHeBJeN
owKqpcnx9oK67bjzKm4po5PAxM+xqYlVuDNZiqJbU8ZKq/HhuN85qNsBa56Mjd2a+OM9oDftlDbz
Gwlsr0YxPjEa9ZYSGhu36kyXx0wTeNSUn/H2dtpRKEIWUiCVyeFNvqcDYVgDYFkscViVD2/vFuPW
Ao+YO6rc+HtNaVuWDhfch0T2L5ZGSr+a7sSYEmeiK0Jn94XZ6c09RDHceb8PrvWtf7rA6gWTs2d3
+emaZRfgbjLdtaKonceP9O6uiUECYKKN8dqanHDGwjNVNrK7wfx7Qxivs1Gk/IJD+XEmQXh3jI9P
JLi3YKsbb8DvdeVY7Kg/7hAlVVXm/ztu6BtugqCBimk3H5QiR8mRCq+urCH6mrX7w7fpZIZ14DLS
tfEXczkhXfH+Zwjkd2MraIUrWLIiVBrf4LBchVGnFjh79yJbSiNcV3gSEvxU8nzPIoxg4oYQdQRH
nULYKmOuwV/RYNrZytoJKX31OoZOSytc/lPcIiEsx3Hm7W3jtnp3VEGoQONH8F0Q85/UZyKIcBAl
swl0xmymFihQeKScA9rsHqOIThr9mUS9sYZFGqu7jj0B85epiGYH+s2vS/nCc8wosy326WLagbeE
beq1U4Xtggodw1Kdh9RZA+qfWYysqS0MdUnh8zSZNt/1MVxx9sLAS0XTy96WxrZZ6kt4d0/T0iQs
GRYwsV0jsNHz5NB2aE3ovxxBWUFISYbwzS9SO3Vhw1SrguoKIuK/o5UAHQGB5/yUsCXLQTEb1LOG
NxqCxIMS4uu/AXfv5gRuoujETEHSD0NN13DLtdxE52LvDKo//lPmCFCS7s9erwkuR4CSHPFrVC1Q
34Sl/XfkTPAd4Qzp2lkS5wcybBWuhNrnDNFKzUiJZIVDO8vEg66Bv8OOba+270MQq0HinzabNxDJ
UDwmeDXpLHqL9Ev2l7k7nyfq2PJsn8WDq3TBs+yUCzpYJl6STlmSwijIOZOzcmvwrsAr+cGclhcd
RvWv/5jOrVN0/QNqc2b1CfZgWypQMIdx/gn5Jm8hekelypuQCYMKFI/05eNhotWuJWxEmrjjrVwQ
CHyrfiSKjHxAl2m82XrnuH9IBwP5AiLpxr/trjnSonmbJ9noTThDj5Gjyx5RyqqG2wnS+1uqZBWk
07MXLeiK9RmtIlRDxnPW6TwrNGvari84iXUCY+6BcoxtM/pwes5jKkWrhW1RVxp4QMUswz4bDShr
tNKF/maz1me6uQU16q3GCRrRGAZ4gmI8Qn1Eb2mOPfyxKQOyRA0ZvyQq+EK04S/NqDkzfPx7+x29
Q0FTylwa+DtVim8YZ18IjVlpGb/UgFQ8W+JVCIqfy5rbx0mo9fWiZMbytwQozDwYmrQxiTyA4ydU
wiEEplnbUJbf5DYCemjIaycUAmYv+BKK9Co59GTEXKpjsyOV0PUdVAMAPghnUkkCTziaLCymOT2v
sm6cSUIspGeRL9pby5svJ9dzblTL+yf6gpn6XE69PXRB2SjCqyAfH1ssgtCKbaZd0j3osApT4dSH
JteQE6UW+tsZ0HcfykAP7yH/HwTgQ5cs20/ShwF8NBSGoeHCxbFt/yUXLo8/6qhMjR9f77ycm1G7
jpjLKGURgll0+sDubummkwR24Aoy3jb1RGOHHJ/ZWsWnGL10J29THUnPq30ixgQufJE9htBT8nJx
zJSg7zubGfeZKTUanvBCN8BUGBdVoGy9jxAgO0phdVxkjQFFoEdKxEU3iIkCS2ycJYjfU2ufsbat
0RX+7yBcraYRt4JrZ1LTmudo4rgYNv34QW33GqJA8itemXSW7ZQyEiyw3v+AVQ3Uu2Qsub8xx1PR
KZH+6GfcJTix5/iCmYtJtzaBWzqyrAAn8ghl4GHTcFxcSP7NZtKna1Fg0QOBTr/EcQnInBZSl2Z7
iRxD1mnb5iJqpVsvmeTDQfBuyYxrj9Hplc6Zj+rYNVLw51ExRMJRnIPzyRL5Xc3O1dOs+V4fvE69
9D27y8wfKBr6snW/GxK1bHmj+Hl8CeuoaNuZViC7i1N6LUPRIX7GBMlKjRD3BAWIbTqB75qf25qU
zlYlOygivThtAaCPvAeM/IG/FEjPdUVaFvFeCzTfTigdG/eujWoBHPMqH4cYCi3LLAj2805ZjgK0
+RsCC163o1Rnned/2LXvYYA9ZWpFw2B6A3eHvXE/IUzL6pMqRY3bb5z6n7t1TBbUmnSGpLsbp/lj
28NDCH0Gxl0s8Izrd34EVWeNTo1tjkmSICzjOImaOJrLw2pvT6yilaZH8cTwcicZ47d4nMLrhZ3Y
QwfVweSKnCTcJ1g3i2oOOMp3kjOZo/YlUnfjVVkD0P97dgfZGVFabK2wo4I3gYLXsUNGnLOxGUGx
Co1HW8G/J1exR19IKRmyrkN96alpf816dZ4W+xm15Aoc2ZdHXWX4rtmw3VNOjS0L2IzIAXpL8yBm
PNv/NeAH5G5OgZtLmf6TF7g9NvWxBrJbS2TISdjn7HpvXW3m1yKv6UU0u0vQ+OJ/XmZavXhS7STh
oeSNWKWm2M1ebLcoYcDdLSzDpvUTFGaOzoSUZ0haHOnN7NTePBcKjgC2ODknRJeHM+Gmk+d6F2od
J20gH3VwPMmB0YeTzrB5xZeGGFdHZvVukhIhxAKreqjpHSyNOugdiesewyiWd/ByAhkv9oPcKbm9
nO6gSzLgpzxpfqoAr+7JFjAex87Sz4rsumwRV+5vB+DdFPjD5LdVxhH+TfgO9Mf4YdjBIac6IrzJ
XTAby5WbqtcDeDpU7YXMFHfBhmDoKTZF8zhg7p0/FWkOsb7IoH5R3bG9NT+9gRElG4xejyaNGvVE
MjkoKwlTwRc5tvosGbbdDgaLgruG5KsSeGJTwpT1WXVv2VZqA8T+3F41u2eiJh7OBde4Q52CiUhS
qxn9ZMtemereXa78z4VnG985tHFGvknCWHNmqGYFk2o0ff7KrA9ocnOq+4x7Uev0EXuaswif2RV+
YQS/G7SaWh9q6hS5QM3oLHxfXRse8R1hs4TSfYucH6xPwsKryTcVldcatwH2TEpnOyA1iumQkQI6
0CFzRonESr81RB9k4JoYHUD4wYkw+B+9tNWhT/s6l62qMHwTZD0D9mOu9g1MlNlHGGYcjAKQHHKq
g7qkePtmRuLaiQDY+E0nRJXG/Kh+bA/LvPNdF1qyennHn3DMSooYl0th8Y5+PfsMNxqCPxEKj7hD
rG/zg/xgdjxcoHlj5H7r3hDDQFo+e2CghCxsNB5ChD7u90c5ofH+gU8MxcRqG7KhF5a4y/3i2009
uSsFfLKbsxsoPpBVYEO4Ki+Yz4bPvyMDrfeQ5ljxsrvMud1Zz3oUtky+WVKqKMopOPVVdh/P9dEj
qaU7bPgA4TaXo1r+9AEkD+FNgjHp6q2c0jYhwcHAPHUA0bzx8KLJEjlQt1m/fhQcLxZ13zWSmk7v
MIQZ3fKkkBKAHBgmieNdCCXi273x/8LSf3E39oVfSoVjFzyx9ELjrFhAuEcMoJI//cZrjDQWggtu
9os+tRJDtscFXhItdkAg1uk9gnQpjWaIm5uOfu+01toMuHXxjt6n0zBZMO95O9SA8alweDr/omQM
XfIbvTY5lTwNs46EInGdqvyQZVHWh3kcBR3n1m63DqB2BXydQbs4blEKIX72G+EDltomf0ukgK1M
+rBibY4I/IpBS697A19OpYoE97uDsPM62rixq/TQPuzYDrDpKqeswRRVbD4R9WMfaFhR483lbTaw
ZRvUeTsFUnNGNQB0Yi3+BCSFBlfQVJslAWY2DiCSpHqPmnaeXKl43x66ZuLo9AdEXCd1nzcHBJld
GhDHyyteZq8ceXC+J5j6H+n4MhyjfnWCyjX/k/TOS2FQtG7ufce5vFl4qUNXm1783sS+aIeC4nV0
aFIpMyaM0/3gHjTtB4lqmo1OIUpgwEy3pPR0DsMMwtjTrywAC/Kfg3+2pDRFZ+eWyiq5Ngm8uBtR
thHvxUUWf+ujdBbb4h5uzQSWjBzyJ5eYcs+btfV0LcfXjljtOnoFzzluUNFu+EtUbNtmsTd6zSym
yd/4I1C8G9Z5cZLN8Lzy/Xo8+PvAv5js1sn3C9g9EOFEDV7bbWL91auQBx5Jx0D4rQu2rg4VqYf2
BU/r9d2O0Mv5O2v3h8hYkHV15gBl8ppvyI8tF84/oaMj8upxXZ2JtBvO+djSwzfDEPBqpPMAjm+W
C9p4ZFkF8413NSsgM29+pzVwNvhJQSLxBA6zGOhuHT+I+xEVg00k0Z8Ie7T4NJK8gkNtOWpmXzIe
UNMYM/XVPnzyShw8dggoyHfBgiwIlnDC3nImBDEI3lV8dCdhwW5xCWfQ0JXqKpZmtOGDPCGsEvx9
t+6GtK1yPAYvKZtQeiGbQqd78DHZ8b9KIk+YP8b+4i50Vgr+612pqWtHx63kwafGyJwVMnf0kdoD
k0JBN2rr1tN0DYE4Oz6reJN7vpPne8VhwV1K74tkg5F2cLy/vvkKp74wrAa/zCY/xIHKJhKvP7LU
aI+Ksh0WZB1OsrOpFGU75o4+cZ4LWzzwcFWmM3aCguKAW+3AMudjDCt9g/VcuS/BHiSLWEF5XABf
/FMqcQlsVvoW568lwEiYrdzshe5cQUvmM0Yy+Egqe16aZMINFwwBg4KOOZlid390fHYAwM5Zpk/2
TAvX2Y6AVW+3ELhy5aLd9/BeTur8NacDbCMVxYGG2+qO5raKMBMBojDEAlhuiNWNX9/rqM4akB7q
cZ0uRgf1YhH1XyeXDNEaVsyRILVnAep7EbXOEzjTtlPJkNkr8uKkU9sPTDXQMAPLFFwaEQ/6cm78
FsefHuAjPMlNN48jbED/OWA7ykrjsXKgvyDXb3VQ9uqo3ccAvRXMpUIhOxPi7/Se38TX4aKPW2UN
6AOnt+DykU/HR3GBA+sB6KLrZiVfiSQjhcoglAM/BFNXYr81JpzIUfZxMBe5DYxzsVh53sdTHjty
5mVxqYCgNiucrlRWrQ74TYWo/vPwT3tceZ2FNr427g+Id4HqUmmf4P93gYDgDWAncK+fsn7cMXXF
rSKnwKY5CAAiqshqDfWiAB82snefSC3gvZr83qj5loIaSme/znDTbp2Z4hGirj1M6aHSJ99gIQiZ
2lN75LChqPTDDYkZR1NR8HMrmKs0uajlvyu9to6PRjQc0f8SoDPaAxI1ApKMU74XodZiH3DNGRRl
za1DA5fF/t8fSMBZ9eL9BO0WEr5JqEU/l9TYyIQ0lSMoxXUPKAzY06wiJ0YaLonf8vk4lVqE6T16
LehebDiMTNEYn1oIoel3IQ5n3EaTR4P54ZKxsOdqmj6HcByCQ/ggR5ptrnekBEZfJcn97pqZx/bM
WSnd1vT/kS1793c5iatoyirU6YWdxuVk/KqsoDhFYD9NbmPXgquUzrZ5i9mFveWBwUAcPyrFV4ko
Hqs4v+BQLH/QRiQ5DfrFYHJSZBJODbvsEpqW7RViVBAbjloG8qme44FjvpRNWnlSvJondYpfKBr8
1yC9LI0UlP/uBd6CFt7Lea0FloCOE6mvs2aDxR6WZBLagihhLW9yccEMkoFQ+4358dAsfbe84nNl
CAoamX6SgcWF8i9/ERXTxC7KxwXyGgeqLVCUnk3ImZCvybriOcC9YROYiBnfPcnSVFT74mtxt79+
ZbArcr5uBTRHPhUcnSCsMSYo6D6Hdk5fkA9uqTBfbn6TLY0zxo1I46KLwoY11APD/caLNpE3wUHi
CytFtcyVnXF78g9uW53S8w+cNAXWa5/SiQvCk4xHhxBjaA1+Y6NnR9vR4vAj3WioeR5yK99rdI4x
Ol1qMBjblt1TX4Le++E7WBKWRMVJm6kcQV/fya9b6OMPXFkDQR1hGrNLGn0jw8TQeNFd5GCy1z+G
M+9i6piSn8wkk90TXa4Yzf+Epd5XfEhwGvW+zuMy4Rw9pZxeXxnPmre+rp18rNXjc+f+miS9rM6y
rbUbhE+gZj0QN12wlzmZ+laOpxuu7H/47YnB+FlySVVpaWZ5oWUhBBFYYG/rAjugXjXCJiVxosvy
o1DwXiO7RTwh/Ev9bepvPXJId3bgzg4gcEKRgMVIhUhi3CUmW47i0raalKV8DFAS+pB667yE0bsu
Y4sHfjpsKoIVWB3bytqLg9cVUVad5UqYvgSm/wzEYxMb3Cen4/zPLxw2AG7Ld5UbfBe/oxod/L6Y
SsbJQJc6ltaLKcvrLki35OlBbNaa1RKdP3ud7wgZBGLwLPfj/JMaocq2K++rCYQwGIs3C2Q9FpYo
LAYMXEyyjmPewqnb+jmAxCnXJPGbNlPiYpWlq+ha7LBK3FrGHNXH2kyVGYXIY0GllpZmVhsPDHhp
3KKjutXnAGQ2LRsoCgjBC4tW+JgW1yzXT0fkkeooVVtvF6DkdunOVxK1n1vGyHvLgnBdJtRAYT4+
M/8uNC7NsralBrPfQNBtrnHWvRvjfDct2f7KL+XfN3puUZsAC6EKUmgNkZb4mRrIRV9iBDHl//Xd
4xn3Dm7nwybvLdnMmDQRel6xiXRAZOKBDs0gyGlHutPYXikSBPrik5nEvOJTv/cO36x9Ha+3MjGF
BqjGubIUirwL/WOr4SMfkk4oiT47Gqqw24UtgpM0Gb69AQ5qT7wG+kR/cQ6s3rofXs0B9VVPxOHK
pFPTYgTBOzj1+Z1246zG62zQLmBoseDf4jXPifMBNRIlWKGIWlLKDdA8WTxFgx1GL8w1Vt1SQwRK
90vjPi5xzltttOmPNuSTbxy++zkAg1wdI4XocOBf8dX82v/uvnYOrKAWifCM5DaLSAwtonZNAMal
wki4ec56Jn5wpT97Gl+qm19Z/wu9XNah4I0w95z3r0ThjOhTeK95Ffyl58wUVLbjbVRhyWjS7p59
e63Gy7/m9aXfY77MEH0KCrzSQVDJLH4fEHIr2ulyiTdmxOr1cZAtPdRGfpkg01byZwRzH0+mMyRs
WvBCGBNLTe+JMs6SNCS7o02mHkaymf5ORmvTbzsMmINWUedNhPUFOLgd5WrnYVFXItg4vO1xZR7B
BkLtA0An36YyI+1fThoIz0L4voI/c7spxikaMD2zR/zSY5RaSkfGSXoJprKbh9PYnb/bohBXd5x+
AS5WBmYfItxQm9TGXHkzr/bJgyViudgaJsWNB1ku0hjXuAfyX0p95cvWdEFCPqc1H9oPvgE1xN92
kmiNGVpIAIIGLKNxd8b+rML3zOzvmFWYF7fzttQrLecT/KTLnTzdu3Gw4WlxfFSZzbiOAHm/Vb8g
x4c/WCTfkBFekKEydCYKrXHnOr70WrVM/ZZRMptXQO2Dt3wZNVsEjJuM63PaF5wcnH2SgOh89apG
MzuZKNeLKjsJRivBnCqUzy6RUKrpbtKqek4y+Nl5q1zPRlzPA2uoP+ThHegXKjNU1TtW7g74GB63
TqfxgNo0k4aPn+jt1V0g9x4DG1Lt2GHKLKLH550WcdxCqQZvVZhTyqoaOM0LcFpxHO6dTmyf05uT
63OX8AcnLo0jcPktIf8FR2YXuSeRkq0F+5WevnLs0ZwBAWCOU2yQjtriBAtS6wwPrCpU/dNFIut0
uc7rV7OJoKnkN1cd9GBDm1p0Eg3pAHJtTuklkyQu2SCLDcWJ6A79Ycey3E6bO91KrpdJBHqriITc
m7odRirn37uWm2QkfsDTavmNfZn5ZTymORUdw/SN64LBumQYFZxlbg0dNz3sgE/9/zULMyVFLAoC
sliI39OpDFRmQvjxUnzyGYOKbnunFoJEzpMsaJhvfZ86Mk3awolz523pqpYySrDj77MEc9agu8wW
+E70/o+8UDWNNU/sa6UuKvyROEL6kvBgag1/SwPMQZzPuOcZoY/e5NUB9QecJkgElb3NC3wtBJ44
MPuBrOjaGGrzoE7DaVLS5rTEhafdqt2LW+P8lSujz9bGXC4q2ywdZk9K8e0GIR/9OAs46c84JID0
jYDLqEqKPXZUXEqx3wQVBaMlLXxfIDdLB5xWKAkPbKRCjO7JeOkGeXymXOv+eQRgTRTiq0nIKJu3
UXeEFYil9CeJjD8K0REH32e0nMBJZQbPxfUTIkI8ZiRoBNdWnirVGMgtpzmvOdTKCmcq68kwuqIA
VMEhJULm0o6G8uGEoJtQ232ixAThtYiKsIVlX+vXOxsMIHfmm0zBCErhXYPYxTElIxH82XAOT5qs
zNvvmncB1eRQ3XG/t99+y/e95ltaSUMZc5PWAx+/M25LQWIHWT3F4A2lRd5s+xP31Xs9xxkwUq/5
LZRxbKq1bWXYcwvwXDV5AdQQxwyGM8p6yEyL7Xfc+Saxm0HPLPHNb/OkHx6+kzc0vhT8rKZUlkXw
CFubq3An8BDo2quRANDvdQNI5zsQ5HmkRhf6+Wh+4KYo4w5nvujZUuRopgbbNvtrgIT4Qh9fauok
LYlIkc55eoFruStMWzhz/gLAAi9iJJSjio2W6AdU6guVqAGum0o4I3n0rP5t6Mclvndk1urhnDm7
IwHpBWStIR0x/DkA285VsL5KwzUvby+9B8jmEBIe+KaBxSnT5CRqEel1tiwkSL/cZYUFr42Iihzh
C9HeBSje/dsMjsFXPl5pjSNfsdA8MiA+oAfbSP9rKpL9WH7IdU1MCrE7ab6hZZ5WbIn0w6dIwfhw
2mCctxrFj89b6ebu5zE/F49/G9zCe4Bqc6gNWPswM7kfLCVI89CFTps61xJv7lTqUMep8KWhGNt3
P6W84sEulSwBqie3jVpUb/kKUtldS+wCoRAq3Pgs6GTV4xliivzE5CsJJXDum+tt/9J359uoZGY/
rLy3bTmoONthoH8Ddexv/Cd2nZQAYzIfDdKgSpdPIT6SU304svb/P+lQYzn/g0s4sO4Liob8Uwj9
wAbNvboYebeLDWLl4R2RfwdExyERA65OdzzTvvQ626W/icyinWPVq2sTk8OU4ofub7m3boZOHb2f
Z1yc0FkQ7lLGlbxb6VfmLRe1FkYtJqPUGlZcuByr9pqWuuM6z9nSt49NRyHJXN5LmhY9K8y5pUCf
kb1wiceSqctvVmtAtdoVsx4VmTWz9mug1t8Yp7kp/UHDOB7zJ0oMsteU4eY10LOlULgzSRxViAHC
fFmqcosHjmQnKI0ixo1eypDHnyHfm6+PpBcIOlD3xegC6fL8QSUIO52s4VQzaUvp55lMclaXdwx2
VCZwRSPwmkS9UcgIBZ2AMIBQNA+BJzuiRnOEFpGvmmXO5aeBUAkfMgunqZpw/cppqBd0Qujqn0kn
SyDGsGzXHUD/oOxRa97QPY9v/v+jRsiF/CjWoVWn4oVeerMUMmzXGLa8NqyJvQqbJW3fpDb0saAX
qS7ldtB2ihVPLXkn2JREHAhlQws8e4RXsCgajHNLQjUKBey8YIN20XYUI0yesbwMIKcgDDttgoWg
XvkgPOkSnrxI6BA5YNwMbDEhg941nGKDlAliCL/SOh0r0IksVY2abnGS2HaBN0+iFJD5o9mhcDNt
pWPtLEsiH4SSoxXfN3kU4xoWQh8TcAB1YhD2TuOBAu5I1shRetlWNnbiLzVaGE08pUoBDfv8pV+O
vQD1llaUbATWsTx42FnxHkGGbIMjzzGsjk56w7fj1cAdbscMIzDexwH+TwczCEf6BDTTjtdg08xx
C0g76tHDAbMo/JOtNFm2yekgRx2X1RTM0gSEFTLnUy81aZp3CWxhHlxOD9HaFEEau3/y4n2foZ9n
PmOwtpoAT9F3zxlL383n8Zc66ZtaOCqyFKLjg38Bq2vuGCWwHGis06wCgknAVQ6J4fQcpnFLjU+X
vkUxd/ISJXdfGvZyEqJV63ewTQTQlXsfPeRBmHGcJhxGl8lpBBWUCli6klaj24kjnjuAvLy+SmsW
7pakXq40uwIOS2SvvOC9M+WXtBuBDFzcoX6lB4X7kFhpr9fWgQgtQfMcN/7XsTMTxFguBe/+qT1o
IbKjJc+ZXQNmIg4zK4IZm+mB//wI2nJyzS0GFv7f2Kxw+pplSktTXnk7K6JM+jhVL2T0YU07kJVC
lkwyVfWVZtoGcEsgg8/VpD9VSPjkgoAT/eXXad1c197qP5wQ9hzD+BhlBUAaRZ/NTERTkntPAeNQ
ZZcLLnLcEc6/T2JMkPcpVTYHVsly4VyiKaDMD7OTvObjc2AnQOHakl6CASh7muJKodsjAFTJS22t
9dV12dDOr9urZKYEObIxETPcWHUhjX58ttirizELPTmuNMuDFruDFwA3t0F65Dxfr8U3H0Brehwp
Hr6AeOuZiMa9v+33tnBATuACPshwZ4nvg+XPk2fMxAtlzbb4iPtbG4gVIj5NopReuU6B0NhDcYko
Ov4ETUHyy9qKFeOHn6qAKQWk5Jj99tEwf/jdXPt5SZzU5/yhPK9hg12XAttjVTjH9B3f2IjToRcy
01sKX3EnwZUjscUOUrlNtvh09VLxaQsNLVARadRZFud+7Vi0RP7vh6AHB11uefU1zjH2XpliZrt9
IsZtMqnSK2KQZsHLngd7SeMsxF+QVyp64yMTjgyrJUenFyRD4Vgw8ZTzB05CWl27iEoJHboHx8Hh
BeVZjUar3aYCyTvLjK+mo1cINpUl+rq/0gA826qLGQfycNW4pcBV3QM2OmaH4xhSvSON3ct2Itkx
Lh0HsGcYBGYGSOuhLBy+Cdp3rda89rrbDhzGdax75ij2PPEE3stvFpcMmy6yXtuy2bXlGoGET6jr
80QhSe3INfO8eh8hcjUXokT11kC11KwW3jfPjp6piYKXOTqI6wb7qPBNTbyOH3LTCXZGm2kCjGpP
kk+gGehlkckQuW6c/0Dh4nubzoPtRd4ViB3PM8FlXzWvm09WGPUV04XHhFtxdAGlx5BAS2OD9ntb
996xPUiZHPnTucqDJ2WNE489QY4TF/hFEv0dvEvfi3NDAiLFTeAB+iAtQG9M5wl6HTrg0W6696uP
UVg2weLdnLbr/C0YTOBMvZSKbHVvUi3n1/JGmd6nRmzF29ByTTGdpBNWGvHKtuDoh+XhWYu2CnXm
cD0+QBTAItzWlhdkZ4aafmg5NrSSPIxrE64xnin9KWSjYpiTtqCCD7VcaGYUiYIaPOZ5M97rmdUI
TkKy9vUtTugvvyyQnX6d8ovh3+cmQ00QBajZjHOoZnk5O26cQH4SDrcCy2INjrIN5h5gC0o4aHnm
1LLXijBxzZ2/stJd+Ra6J+5wvvWB4tKfnofcVYFZUM40Ym3d7yIC7oTac51LGRI/1Eb+Ua7CW43q
uqU+D2beZBbrwoDZ6iueePOGdtCBFIvwm0tKccY7eii1ZUQeFMaweI50+DxrVovC6I/WKIOx0SxG
3YfUQVob3yD6lBwiDqulmAdqju4TrOWLwbE6dpP7BA0/GHt8BYCHqOLMyZAMIAzCzjHKChYvYv08
wEkX5QpAoRIuf7bzcB8vnfZ4Ogm40A8U7cFGPMUvVEb9dlMaT+rSWKzcoSj6akwaGLcjerxGZVVu
MdjUIeijqrKI4N6Cnwq5YbY5JBCxc9hW9MtuMSE5UErpkYn8//ACutL5YYwk5WwU5+q54jvDMwjy
hBG1qiv9tu5qC3GHaF8ZuXE05t89UQcF0PnNCzwXnbawMkRKfhMCih5+lwgOVh7zEBv3TtV5RyG1
7yU6Phx6tETviGYqpHjOhtFaf9uJ7JHFVwVZ0Rd4ynmjvBSGywFWMsmGZB7GNMcBWS6tgujLHlt2
g4jZHD5PvAgl2AYRMLENGXc6YIBp8nWu9D9Lul/snhBFMPl8yKCh8kDsi8aRHX5NCEvqhOkdV5rY
XPK2NHPMmgYyqMzxmuHfpFtIDWvPjjyNchZz82ion06cySuXQmafSieHs//BBfFdz2pQvEyyOzPE
Qu0be071iw4aAvauPu7UGVWV8QGn7xN2ZDmSJ9AzSgWWnKeljE+IJ8xI/N+D9VAuXjZg8hYj/Lgj
5vrkx9lveCrFtV2yH3G1YQEfj74/mDj0L9i4P8tqUj9IXvbQkcBTIJqLcxRYVzLB6hfhCUzfpyVY
s0AiICrlwOsiGMxVmt/OmlBVvBXywtFI7PxJ4QEaA5xiv1x5s5mVCuhdSs9o/LHSVqYjWWhN3KIg
MkE2Sr5oKU+VFy56VLNOqOjC/q7j786dYf050R3R94rVuqe3rAUq7MQXX+FQRWqLykg9py5tLq4a
/Culhr3cvhQKB93M1620twilBcCU4LMRXo6Omca4rcDn3QUCsjMjd9b4Wva4mQaETJ+Kk3KbgbvO
6FbT/LsOepU6mPjVFZJr5qh6eKqAHuSnTryhDbBKkLEYlJhw6rFDTuMMZ12Lw6lGWpmKXYJHOnuI
Z3DxWntBkl9Skn9Ck1ygK7Iwmm1VL7j1GLO6QgHiE/LKkT9D4BnPYDDHCKxrgrsjP8KGTjZNHAeA
HGgDqT6nplRj+M6dhiMrnZTlrL1ctha5PzHIjzjF/S56Ja4+Mz3Xxai+WmGh5v3UvkfX1RDbj5Q4
P8DHEdteVB3EMaz7pfj90MXIgeDoMjSoDqwWI1nZ81pDz5GgOKbe1TlCJpcmeePfmxNTRzv+flhb
++c7SwIZPN4fUdVMzkJkQda/HH3Kj+dzOoemLKK+5lxox85m5lV9nqQZ+o3E64nIY3Vodus1NoDV
h1JM9yRaHGTa2CWgvCcX4ZKUDfCFj90NNNrffF/uvjdISIkEThT2Xg85wo6yjfLYmG0JTPt/4NYk
mU771UnJ05E/jNjW2Lm+qDKOeh8oRAiJy/8Ha06zfdzeZPobB/e6WoNAvcHowbIGqZHzfok1K/rv
I1y23WLUQYfZm3UuA2vqFSCyjuMgyPGEzz40zBdNXvdI/Bcp8H8TArZr+KXDVZhqLcUTtDic4qf7
A/rfZxgRm3sM/xoUX28TTOHnrM/63huyV3FhlqPdvkk2VxGI9xbk8IkIOSSc3oPIut4shV5+7Pxl
m5riZalMgipH6uFHCHjpdxjrb3Mi7a4SW0BUbhmXrFc17sz6xN+PzpWzo3ZuPDbq1i/c/o8oR2wD
Qad8C7E+4rfxdc8DPkSoz3GTEohqd1BjTcATlHWVueI5fdKG9Ihd/FB/feqfEs7l3GfI5rtd+Mwy
b2Wg4PnoTZARFbDuGrKoMrnTlYslTDg8hck2hLyHiVtT15VAsBsXwwMUXp3WkibhbC24e+n3zfYy
IuvfjVbyL7mgIqnkrVcajfI2mknrLtTVjxVTCp3oqxyE5PnZJb2g9LEIfsxZH1Lm7FZS01al5F1i
3rcMw5lUpUD5wkYaH56dy23gZETZt4NK8HSXRD6pkPPzC1NHsYm/6QQc9nPPMm57fpDz7J2gD3ke
JNHkwOKsFVS3ZImGGId0fOH9bAhHFas6f6KPIDX0j+pzSukArGNEHNJHim0RY+genHuc2KOqCC4T
KjM95aU4A0y4i791tcqBCdPweIOrSufmgpDMIo+ELrdcx7TP51uMbCDJWOp/7nyWisXmfL02Wk/I
F0tu/GiwAZEF9oO9So4HXbFhAQDaU8a62UtpwvpmnKsyYIrDr6t0/oNqFXLgPeXNz9su0JruNmEn
JrjTg7YXtZaUpyHAGvc7wfvdD4Tu2+WHyGwDIDTSQtDiynyTX698VzTVD6DsIl98dxRHUMqIRNSP
XTJqlq+AZGQRKL7qXp6tOSXOOlqFADLxIwL1baote1c7xzD91tAtjXxutcUaZSi97MWaxzQ/atY+
icg+oOGcVQib0t50ZtZoS5apTRyxv9Me7PwU02EsqiGrHhilU2BpAlL9y1B6NsNVvBkhUE+PUI2o
uk32nP4U17TfocHNe1tRueW/SfiunnPgfd5ojTr/k7Q2vSI/pDZOVAPQRzTZh3CSMoNnB1WDIL8h
SBWaH7EVR4eKTNsqLqDlIg5y4yRKC1lNgVVxA7IFZbgn5oopFGLC3SSvpQkn7BrRWNJT2GOxZE1f
3SxifWAkCoMx6BohzlO16ER3srYHgoCdJNHdmQy65kp5TFT+5viH0cj9jxhNhONejR+p+JmtMTmB
RvlgLYPKqO5/IG+zBiax6jfnE1UJQaXCfuqlX4vBRVgVyMgVg7LYonKc1bSNXsVyFln29NuhAG4w
lXPvldKtVfCIsL4Qh+TBO9fUEUICVgGG6BKRD47JOWambA6Wvc/aC/w2QkN+BShSwLs94wzJi4gX
RrCWKCDRbQUVwPoFoUnqUhScN3sCeopWb/P64xXjVHQlP4fROvooBKFr7LXBh30erpsgjy3/qVeX
JNR1y1t0MBIA1vJ4U4e1+OdprkYfvc86WNh4H3i+2ylW3DmrMq3FkqVC/LPBau4yZ360c8yvY1j/
0Sa9sjacqG7oWCXPummo2niOWewr57xVQaA8DoeQpPF4ZdjJFPfB4xt6B4ZKCcWIKDtze8JwZ+68
/rL1ExFSHK9USh/mOIgZpEtJwr2AGxzzwGrAWU0GpdiB8SdCKVuNomTLszd7CqapmsFqukO7oofe
8dvSl8RN2RN2wyc8xFWgd4t82ki4iG/pRtJT8BKMe9A3tCMAvI6Hc4iXfiUnnx7RlpW1is32ULmx
WAj4T2FGFXwhNbH/CnrEraPPjpW3gYzqGcN11+3Qp5ESSOxU9lUtyTeuoOfyxIMrVWa1rbvXZUJR
t7F09S8pynBMC6nMfEJOdT6i2baogvubW/l/F45meat/+jUfyXOx8Vwzk1fTT+CSWAtNgvozyf/5
WG2IyY/uyXmJzyXV4VknRK0wTLWK67DL1fVOa2x1fVGOC3dnyZFXNVun2xC6N37tWQhJpxJkAK+V
Qwn4sTbUB03M3p6zDAxwWYkxpCWVQvERcoVh/gI0Wbsivy95GOy1+yuB3BANEKR7TRYl43oIEU+p
2oMw5lffLbrMsCierwfcPbTvaOe+5GRh04EMklJ0ZKf2dIFuMkO+XCL0gnQsHz74Cz5rZ8U08jOQ
HPeFwHsdVkzgKYbXTFticoCTGqFynUbkQ1cdUWASuWETIw9DInKosOrjj/f/pUX7wGlZGIdquIQk
dZzy6c7vwgnjiPRCTfIpdB8Tgon51VcVf8bdyC+M1iV2NSsWz1/EalRaT6fqSe1fVFmUYxQfDepc
ohCzENCVqLH2pHLE3MK9XAjiUHXUC3FLTFhLZfdoOv0+RIl7K9Rmc2/qINEvbtlb48sv94eGfNOV
yxblMmkMo00PzRHIoSNnkRIXl/d26lFdpCd6etEZ3pVpWFLNurpHHZrPbL4W8UdGV7Ata7uVm7FC
hL2me+ZZ4KHwx8eDI4b5mksuC99VUreiM7FpxR1mN6OQGzkYLIik8looqNEet/ayBXMhH+VuCoJG
QzwbG+LrwJ3dJRQYSon7MLr0r3Qcaxr97vQaTtolZC5B02FP0sRBjwOacS6pQUSnUy5jhl8CsB2m
HnLDeEY4OcVW8Vk3cb3oBgcyDAFmcuoTeUhELW4BzUR8ICzVXk0uBIhRLpxFOPGRv0uCVPOTATUq
0AyvtC3KViBWPvml0eOIyVG/Oq5tAhCRJI4B0ttDHBSHPhhF3Qb1CRW3n3xo7CpprUPVKUsNv5TJ
U3cTs6eZfVPxyTPzFZxcl+c+TSTM+8iiReRgaGO8p/fN3/OenFxgRSuLEjimBJddmKZzDQWnxl5v
iQ9l1RzRvbZfNtHECagErz7hD61i7tvnyu2C6McRKQmTIplxpDHtUr6qiScWd28mVstR6oIrmmnJ
8+Q3z/Y0qhEGUEt/volN1oqv+AqyFHmXHqx8C/KveAYI3dDeSFcZmGDmtvF16An4cMJ6RAqoMKfU
WoYY0oRhYIuzyzJTxW6/qrtTmujmgC5qu0uNNwDLKOHJUR3SPFaZIkhF0wpZHYaaZ4wz2wLxoUc9
KZ6UPONHMfv1CB6mIzRRvV7SJ98zG/Jjr/dVxtPoCuaMMV3378fJkdpFssrDBSGk/8D+SpQ1dKmu
znYngfJHXDU1fSgDjRNXjIWb9tr/OVZM+ArNgWqAIKvBImG+s6SHJ75GA7rLsbScBxnxUwVqsfHU
TacPIKt8Trd0MqO8CNCw1YM8GVXn2T5yw0o/WWkZjpN1JgJBTrXvEVfUS0LgeJ5YawrjrBrmfJuZ
PHWP2uEO5UPIyNjMbkNORPOOJFgYva8OB9LwvZfw2zN2DLoqTwhEZFereSdKKlmQ74JpIxyQOb8X
30N+i8HnOI8q+t9BThUHz7o6uY86Waf2b1OzcGitJXQcBsg6dFIwN0IF5HUWAtvGPhn/Dmv7KnA7
Zzsd4BNqKdyO4bbCeSWlFIpletE/JiF2MRR8yr2w8CvLs6YI1NI5e79AT4+fX8TYl1KDK3gT9pnh
j6Zb/IIcTQl5F2ldUF5Y3/J6X5KKmnGkFW6bSNXsxIclv25hx2tKJ/2twgAk90S8WAXnQevMq/Km
ar+DKp+U6OTkDpbwr4h+ZzIqygbkX+p2pP+kyZP0MkC8oOvKXJ/FCNTw5cWzAf7etxwKDr31k/Hy
XYXX3Nuscnax7e3hrxeGgRKvS42gk2cJ3sxxYRzei1h4zn2xZgH/GlW2sj4bZhexuisPzTwl9cIw
FuK+YSqs5EFrzmIfbiEH7iVOf/iptg7FTosWuaW4jAtwOQRvU0xZyj4U/V3gHd1XGPIk0NUz5glR
RQtrpmoKyompSIiRmshqdgLeGdKBRn9XgSZjj4jjGDratB14oxYdv+eu00JFA/qzjpNB09AOWBgq
GQbsIfdorqEvBwXBkLGEcdEmiTYYiCUc/4vFG7UOpDGZFes1uGi9Ykptylq6erlDfhRQcvcxD3kO
rCP/XzljAPAN4P1wlOnWB8Az28paP4C6uuWgsN5GFDpocowu0cWfI+AZojaSsEJIqjgiiqbayGxO
eQotcz/M/NE4KdfokIJNcostpNnyiNtNxEAXvAx86iA0FhYDELnDWDP0h47EZjIjAqQ0Wc5QUI68
IPRIMoNZHeO7orXQSICck8JFAfhqKsa1r0NS3OeJaCixEH0iOHSyP3wQVOrtE7sna7k2fF2Jik9p
vZCddWaKVlt3Vb8bkqAiwkE+7a27UgmqAJZeCuZr/f1AkJJe05KTnfm2dGuGtwfa9Ww0QyFISe8p
JIfysZi4w/0QYFtL29wg+MQQwH8TfWGmOQVqeijfMZUVaAJXcQQTZnZtLLkOEt4klPJuHUfPxQbe
7FIjSFbbpjkqh2xnSw1R+sfsOTGviLcBC0orPu4eEVY2vWJY+CJ8GgseClNMqFRhpjEDtR6G4F7z
FVHPRQjCJFIZKdbJRufMt8NEDgGoRbjK8oVUQqa9zYjor3ICQ5T4dyyA8AbMnPqQOAoptPR2sDqW
Ki58ifjJ9it6IOUMhnFdjl37r6tTFmVDqToB1JJBNFxUXj5XJcu/hjwxlYzogEDqQNSwdibEDaIV
oz85SmU/sW9z03sn5Ro5Nc/e+11U3Ch3v4m5uUMEs8vsmM+oiA93aRhy0WoW4+2W0dybs5dGYd6y
NwAqg9X1FJi2GmPSxovEUDyHxw//y1iyTpfcWdqQaHVJSqZ1E/AK4BQymIKY+wINf2hwCRugTFip
YKhLGKlXfMMl5wccst6NmoWXq6cXzlTClSG7yz6F6Wn/4MoegJQaJUrDHgTveyodKOKI7tbO4Hb8
opbTnn+ZkZFd3M1MVZ9p5BFljyPQt/o/jG6nfv5sYAfie2D9iN8WR4kH5RYykjtyiNS+bGf+KnWU
SXQbOkCOT+3kQ6q9RjuCTF2zCdhX+uxBavXc+2zmzFFJ3VvbNXSf1zvg/dpI3zRXBtBnH4OVusOo
fKwE+PhVa7WsmDRIKJmY2VeLHVGVzHEP14Jz8mIFS5dQKrvXmq+XHyv1/UJlatbxuG1qssKqN7kz
uEZBrmCKHuxwz4QXTXlFwkCBBsiiMAuaAoZX8z6GSl2WYV5oz1UC5D5fxlH+AT1ENngu5QZzL51T
Qg32u7boMs4lLLOlA92eFyrzVQ5D3y7fEzPyw7ibyDIEG6HcFXnAFRBU4z+KnMOaxQnJvpnq5/w+
WWl+IaR7iCQ4KgrIjFHSJVZ4JGfzbieUnZ5kYuoX2DMcJOtVID7AG/bCE5H2koO4Ywetywg+taaU
Fpm/Rlhb/W3QNOH0PHpdkfNbeCHmZAoHU/gNfVTE/tiXNOu9ePSXOQwz9W/tu5AiyhZ6tfH7DZzx
4/E6N+pkXBjOsDmjF/AG1rDEBTWD78B8UKSe1aSicQTN0xDyacscSRz2IIpa5gbSfqDIs58qQzzK
7yK5kPVW+a3U/msnCsKK3xh48JtNdLWUGq5YJi3XIev0jGyHW0nd3g51+O83Ijib1ugjI1DgR/+J
Oj13h1AECVzHpiZFESpNxLYgywF5ewWmrH5oSF6Cf3HEiNZvwiiRtguguC3LDQAxHUHlB/lGGakV
Bz4pE/T1x2fXz6W8pK59dd9BZrvQiEbtX/hqmludqzu7EM64WGtb8MQfmkRI8acMYBzDNARh8m2T
b2e3pULus/FR0j78NVaM7LMuGtj8A2C/otEDYUlJOxBS9m2Au86d2CSq7DwqRJu5eTEPJDQQk8rh
zOOJW27s5SLs4wUxkmUct6raP8C49qiL3BPI7BG8ONHpH0ZIjRu+g58i4H0CE0LaoySYT6sns3ki
koTHePSHD3G9WvtYsVSMvgQsoDH1T9ScyAKNczb4qNB8NeLVNtXjh+g8y1lOh1zesAqchpTkCM+S
gdlVRoi4YyOpdQjTG6UVwdp43JozX5wNTMDEEtoWI4pH95TqJ2JNzmeqABErcbzzlhBSyyJbz8or
QPT/DDCNVgWyCUSXg54JbsGVW6MuVkHiMy8dnSt5ZZmo/r3amCrf8SjTm2hLnQlBTTJlB3NekMw3
CM4Px9UvTkwDzTV564bLdozUVNY9GLCXQr2pzE9G9SlSwX+iHjdYN6ka5p4hAvp8LTjAyEE6mPDn
PzAT1e+7zSTJ0DKuonwFzo2mzabFbKbm9RGrxTV9ZxLcZ86XdcXgCI8h3I1wEX8i/4LhELjeoYGl
7aKvZy/t35e3HoB2O9C+f/eWT1YID4yiTgczKxYC0La59AhJFRJiGI5HAPsu2u9btPVarrTORe+w
d0wJ8iQg7URVqlnhpwT3jIgNkHHbHil8Sn+7d8AFl8/9usC8khiQHMymCgpoFdmMD7AM6WKl2z9I
q9NsuWChWzsDgM1xLNwYZEYEiQWtqhXARbo8sKxgL76ewABO5jVA1Xx8PQLtyt2zpVyWup1LUCtY
Tkq6EySkcrx9V0wqWpmKXjIxR/+lSpB0qH0M9j/iLjI+leAwIWPnwKabfHDtSh3FrMP/yM5vDzDG
6fTHiA5+gIyJ+4WEnRtyTuLO/GUSX3gsUxp4m9l7W28QGT1FNpHk2IABRoRPM5ngEQTMMLb9fC+W
5PvjDVVfzylaUAlRjTjpKzZ+LCME6f/ci0BSRypNHIVl/mT5uYMashGbOr1W/IKyQ8h0dfziBxi7
jb9nXm+3R1O57j1CQLpFagjTKNe3VrgI4Qhm4sOPabFTETswTfHIkZmVL5zbfdrfMghut8/pEN38
WsjSpXx/3JySOvBrFlwSyc+vCNOc3+yQ8OIu1WVrTxu6Gq9qlpcOvE4ZUaWXUW8l/tFJwgl2R82u
vqyWvCVLch5A/SA6paJtw53otPUBm01cMEBArLgD6/Df4NR8gL1C7wwCUkq3GKuyWYYtEDMGjySp
rP+dn/7p/MVeaLfaptJUXCvAQgWjrFZehPiV4Q8wf+KvsKE+25F9kff9rwBvQ7Vlgr7FKrFCbk/t
sO/4KVBzv8GqRXFBtQICI456GTeYsWOtBinfFWd8Cq0oxFqA+lZd/raZHK8heGx5R8FKMk3Di+dR
+/Vjmiy6gkI+YZ12XM+42XsjIPPQohqdpFyuACozZepNzVwXmRNTstT7wFCxjqh3fIK7M5Ti52Xw
Xh7dSEi+qFcs++fuo/mXvTiz85740WSLJOQAQcq0tuwcaLKnrG2huU4mTICHlzMYLEAf7pDnVTbw
xDBM9lp7ZWC49SW6q1KIDL6nPElMpy5tcdp8RAR+BqOLpHZj2T8Nbnq81VEft06MX6OcaHZfbOYE
vLMEWL5UH7y5WIQjXs7wyKviYuE/VsnCeMM/RV7HxnovVT92N/5mT2LIY+pcHSqlKfH3ucl00MHI
BeWOWWmUB3divgM+dtrwTINno4mRhWF5W6ppVXUSdtRGFHl1VTyKJV5h20ySBFQVEXYqfkOZmIEk
PljfmqzvDWcr+rRiF2IYIpO1431ITxhYI7DvbtWkcpuh9pOK5I2GAzz3FVr2smasH31WfKp9/m/X
SBpn/E5zNcD0Nokd/1o7oGreH/crSdNm1XTlB8H2bE5mMl2PxlBYS6BmWsqY6MYwFbsIWiRpuPfC
5CrNQa+MKLJOpEFLa3qSFamcNtII4zhYa7q4DUG2Y+Kz7JRiOMKZwf8WiE2Z8MN6+JlxFkA/zukF
ngLQ0HdrDqZVdJyqJSUhNQAnreP+2VI0KPQVLUj+byQM2kfSNMB5DDeDRyvUI5aOcdbFFlIOsjXr
wZSr8lKbX51og7d1xmkp/ec2kQTUxtRnshZ9WcE8nYiAV8da9jfmaKDh6Ss1ts1JzTCI2mk8eT/H
pMi9Gd5EVXbwG17cNsNIHrF3RwyeHlTxd7p0prxT8xg1ddFikmBIiiQAblDsCqq01Te0i2QD0IJi
l0MOKFysyMOvxKyJgFApV80P+3vq9D5lmYNXVbu8KsPq0QUoslabpmkHbLzoUsFbiWxSz4CTYbp5
Mi53Z/Vj1r5LmI4FYT56tjj3GifYfPQecxKD6JBJIQsdyZL/cEl/vs0q9W8F+pl3ROA4bMGv4SsJ
brqnq76CskNG+tt/zTnZYNCkI4hYqGiG4hEFQBQkOyALfes6lfqq7Jnx5Quq5kxXcj740xrh4p/0
XZWlCaukV9m+7siuiUbbaNszzVw2uHtFrmv+Vrqy6FUfNqSVMrXHqa90TjtGci88xRbGGiBJgOfO
aR8lmsXGWMOYCeWzXJJxFsB9yyRrpKIgLUgU4yi01SYYoTV5m5NDhl3V1tPDaBtuZQ+orAPGtmi6
5bj35KLtlXd1CxrnnCUmqEbihutHMWOsPL5Q/+OjLHpYf1u5eq4w0xwWWTOZwupsx0bjD/paAl/Q
KfW32tYprtj+1lulVh+XEGp+x61gkFKdN5NB54aNzB5Uux+ugLRo3DqoE2Ju/MByAHMjwcmjrSpR
9DKZcyosTzEXGQmctOo0cjOUfnDS+CMrZEY7OiTKPjjYo/yOrbLZlB8YPgjJwMiHCZ3zsPr6ay4v
kVZ4pVcFLSc/XLGXsYzuj3OARdDriMTK1jZgyZz7Yqz96WZjhBLtYAnN7wAKMXEo3RyjIuo4bWcH
GM6/aefj9aRPHK6TRhqGykVCEYNkn7e6xPEMOPYAbcwifswZxN8sB3NjTKqNjO9rmggctX7tg2KV
RunzSSfpsvtPKnTP8jo2fCvEGLERCuuZyryI9UOMlJA3dMyAaMI5ORKYZlL1gS+ACbFzZ9LRgpzf
btnPJHOuTPFTy04CR7gOHnDOWVBn/GrX1Jmyy8qd2mLcVi7h/9c89oQL8aH8w6XQg5cDj+0nHu0A
tBqvNlYLjXSzg9Ee6H4kDfY9owfW30FZOqEmjN6coVDsRVIhUChXqlJsbUXR2bAhHgZDN7h4ZY0v
hjJ2rbwG8AOKjsNH0z8qzSL4+LCYhL7bvWdFXmhVBTheUjHhNu/6qa4+b8Sdl6vUp46Z3DOPThGL
RAO6Wy/eVsI/SOUwh/J48WnqUArxbFjrrWiE8MdXSQMUt5bLbU6C8Q0wQIchwlLrxj5N1VNBoRgV
S9+dNH6M1YAn7lU7JcaDy5f+7+xq3nUmsTH/sSV/Lv/Mwn2eojAufIN3jv60DesQMv/hir3ELi8I
NTsaBUxiAU0aWG5S6LaEheg93I9/Dfew1uXxPhpFLPBB5Me7wYrwRmhk8S1JgtHB5uYRweASDJ48
0gIxqWIlF5bm6L4ObLzyYOb4vkhQg9b5LJtCk0iRPpRNxDg1bG4bImbkjKfe0YguJPwTbG03+ktr
tTlTwBfD1ihClaUPwDKkMvacKMJknvYllssR6Z3114HxQc5ofnwLPPo5J92CcuIviP+3qpDZtdwf
+bg0U5Z29hysG1pnCWgA2yQEHMbHT9qwfoDgsUEphPSSbUry8vy2z4vfIXMKociJVsuV39kEkI3x
56/5M+I7t8GIoep4W9qY6e/fImhfcm1SqDQfHztZouvHjlE3Xy2bSL0pbZKevGEZe366TfvLk1NH
9EluIZkZAGe6gX/bLxROW+7o1IM679PTUze86Eq1j9+noetdl+8ARctogRHnC2NOkE6yKoKTeEEK
QAPlVwz+ZZOXS+LuvA1043HehKAwAAhwRjKGmgQuTHGaPlrVns4NnGGep7vG4ckVJeglXBk8DlvJ
2oyGS6342JjLJYoQU3cefT+9Rr2OA8I/0yHqgiVdMclhOUBhoVr3V/w5EcRZaGDTWVfihrGYqUap
1gtIgxbLMbpoE2+pxO2YJbUxCToFJy0w802kaGtKwnKRMeFVA7D+DEZV6LFAQAv6pNWQMwPfZ72A
n9lRPMp4tl0dE5J6x6PdWQMJ4JFF5iibYUweKqzDSEXxLJPZkVh6GrQYXIFAGqYmU2vkCMFRH8+N
VVvSiUz/sLNuYPIR3IAgEJQwtcOQnTKzBkGYkvBtwu951eUJtBPcC34cFkMzWpWR4Bh5mpdrwumO
9Jc2B5j1qb6yL2GQzDMKrmQNokH+zuSbZO+Kx4i15ff6AKPRDJnFzrzBMcOK9WPpfGB7Z3+A8NX6
pUjwV1a4XsXA7297np4V0s2CDUMdzYG3cZ6ZVa7QThwAMbw612QDdhNhTkxb4fKgo2egq98k5Dv7
2FtN+tWqb/uIQz5EFH3IyJZvMe7ffEAhsfa8mISjfUkvJEJkFKf2azEPM7KPnKkvhTBQR3WEc0V8
t27f0OwwwEqIj5D6M+Cn7W6jmgt0uMtmqRejHqx6seGUcLzKGKVDRY8HIWJABr6YIOakORM+1Byg
GFg8J5JNOrj76yMf5HoDjrFBtU3YUMsbbdbocuCG+GTU9BP+mHU/rKG9eCpKQYhgbIo9EFhrdalN
y7FR5n5/ERy6k5qaXHB1ZrKXtIGe/izZ7Ef/W1YLhEeTWon4Musosj685ynb5AZuiWAI2ou4TCkk
l3hq64PuzVUkYjOcaEFNRTtN3LwinLfy+1rVRnRPc9GZ0yQNKFMBNDXyR+8e1aDCBLCOo42c9SXl
xOwVwAsNdwKZ5zp5wU6hI662cKY23zgUYKSxePnll8aXTu0hA1KCwGti4yUMWa+c9toqcy6mH28c
0jfwgfgEqoLMbskdGnn5zA575hPNPZoYosyzeOiRdapqaFHR2d0UogeAXM2QfWc92LvYwo3xbHI1
MmmS7qq591O2wC2Tyv567XKprfHg4BGgPSq8pKnSKpmFjf5H6cVmkJxyrORi3ggxo60eG6y4DQRl
vUvBR+yDTiuDtFdxm7krfWZWqPLhOOq09mrLr9+qg7WU+QQNDvWcDg3wo2rwzGO2pIOU8gx3zjQl
hgOOMlLXbxGEkSaZKbjOYkeeyTfS0pw9n4uYQScxfoaR6nF2jJQSivyIcZ4qBuYjkZqpRFkdtpM2
0h1d9ISrz7CHUVsBWsRrm/r7K4c7KgAIPrNKUqxSzisdB3aGEgE6HjtdE6G0HYBatfcpzlOTDb3Q
DakQy5MU/t6lA0US4Lwv/6cWQQBVQKzp6NGS1QSetobFIQcm4ufTwahbv3BPzb1SW56yuXrgX022
klgn7qJYB/iZ5Z5hA4ZpqoFYUO0pff8zFcJFd/rgfthv0Q92Z2FJ3fHqLY9RJcFgQkGY5rbxVS9c
JToaXIisC/ngYOgvGtaaHM8/V3fa3X/gVE73MYNM+rv7e13UH1ZG4Amkk1eUOGCRZYK4l5PM6mAZ
V5d6Ds0MjuHRYXOzbtETUVmHf8P251/1VjMGUmmCkhj7qfrsMCcn5K2eKeu8MxAjWpu6BCF7FZul
DXKxpAyScBHDsws17LyaxgvcCAiYzhxOOgkcdBYZkniFqNSOSKnaT/6X+amdaPb1tjynFLTCU+Sw
AK/LDd2g3rE0dzohB7ElM+bw5PKIdd6EVZR+GnazchllW0A58G+pnN3qpFOsE4wlJ4LNGuI9qWys
UVx36kEQbvYhFTIOJ6EdN3Syr6R9oZcivrfJ+E8N9F9QGlnoyqP+uIiBGzdRm9OeMon7OP1blgKa
WI8FCFTdqnpauJ+FpuHBEo+5Pi2n77aQDw/53admJj53BH4KALaMoI+YSzJiorKfWqrB66n6P/pS
5tKDsj9Nv7S8r8hMKoZYR+K1sFdb6U3PYH57ecpKu3MF+o72gjvNfpiQJyq8Wl318lbaxT6SKhW4
BNxYgCAupZKqUE6xl8h2PGRmhUmuQarmh5nXPrzv1WIwMrQ3gRuLkhCheYdFgBsXXVsHaLEQp8rL
7JI6JWetn/bp2c4NjCX06I/XNMpamK2FqAawkVm1ByxuWwiFtoiJyqpS0Wr8lwzrvj+77UkzPx7r
k1WWu49h5hGk71VBctm1cyyDRGBlVi040KYXbGpA6UyyNtzZ37CZNClLG+OSKOlCTf1vCH8WoibB
l34ZB9OLavCRguIquHnd2PdZBw9Ene3Fti8BeFTRsQqD4qISy6icqr6VesGxNPuotTEa5jQlkFh/
HktB0fiRz5+ZsOLdI+z4s3ENG74LJ92SksUT31PCOJ17hxrqTfPVUqdyuRkt0NEm+yef2D1djyt7
aANGw90PUF9fLYh+94Xz/MUJN6ODBw/oak4CWfnT67eekW4NnUPDxGIa1OzYci7S1S5pjxlYo5X5
Up5x9qEqWZCkBDyNaxC3D4t06eAHV8R2k98tfimYIG7IV/f83bwl5CitFkyYgAKB8Q3QW72QH53F
TjaRDFjbhutTEAl0N/JbytWk+sZFDo6ZHMKcxbFmKXgN47xhHy8D7LiBjZMCBiv7pEsaQIE+64Go
dTlB5n43IoI7UZ/CYfRHlvtCALn1JJGNQMJNwqE1xaTEg0Z0BCTSdaKbyaCybStR+qutrSmR40XP
12rcahiLPPInmHOx9XhkR2iKb1/wMTIO15zRvtb3/YiVgr3s7+ax1FDn01nYnn1A2ooYw0AKpDBY
ZGnNJTbp2VUFZ1OqqG09Pt6Pvm8pr0tki+03XcvlwNrGCba0y00ZK2wEQB7QeZS9wRW3Mmi2shU5
/9Bi+iFf5YIdv4CNF11yhQhLIKWYgwEZYshxmWs3OGabvWd55bcw5DSnxoDGssKMopwMJPv9PYvz
4ptWSR+qSfR2EWefTHBlB5qFw1/ysrNJUJEb2FnKQ3aeGQmdZEz2F36oo5u+18n+yYDJQPWua3gF
taPxNGrdOpgQTopR/DofofEwA1c6+eCoi0y+JB0hdPa77EAjURbYK2KXte+qOEWGFK69C7RjowZt
7ZTwgmdMyAWwarLdQAsgp5cI1dYJC1/sgpWwfQblrkJKvz+3byT+Z8DX/FKwe35yUXvfwt8HSNsQ
ajC4raOnNOLaBimgOvixodfJqKlvV7NZIhCjQz4ytbAGm5deRTdHz9LbkiWyTE89xY9zXhyTJUqo
XiZQCH7xKu1h60IoSb6KcKkLYB0kceqwjZlSfU3xGPGF3k7cxpZCV+eJUKCePgppLTH1ae2qNQFi
BNiiXqFQih/11fjtQ0ZrpE9PNcLW3Hy1cfBDI1WdIoQG2gtZ0cAh28G/A2adx2McCLuDXK1kXKAv
ivb/hwmHUEeJngvmJMm982ySPomFTm185NMfrsGniaNbKKZMGirOf4sUcjO8pj7fMROJ7hGYYhU6
QKMgybMQnC+xDVE8pEbWur/Gpzf2wQNUigIxOrepPigyXl5kA7l1naO2TiUafKxi3FkdCpwYY3MR
eNa2xrCYIfrIDyrCTPjpJR+D8QFmcHDQDd22CxKZN0oPjK2h+8g/BcCpZWFENmt5bGUHKXanxUAy
ygniBsoOIVzTaRmYpbG4r5ec2RqjWQSx5bQ/IMcfE+0HObP3sbplcC1sYAOiGLPirvDrls81T/pR
jmj/aLR1XgCVq6hsDedUzyG82L0DPUqMolMt7lwP4t2gwEtoMYmMgxoLMwYwrK25wYZ+mYCIEF3W
KOdFAGRbwVCrJZZAGHjdKT0HSMIwOKUx43D7OPRFdhgKqcsjXJ9XsIq2MEmO4LZy0eTCAMaX3or0
RQp08m0W6Vdb4n1CkUapqb2H5Mroiqucre+NlcCcGSNipYXbZAF8lgWxWHOeHIvitaF5SR/FhNVA
4Nb4M6e4gEqiz20Pu7AchuImifi1hJescY1azKfRmDJv72kzw6iVwVrQwySg0/uqLCnc0sS2xOHT
a4U74IM8FDlVpkhROPxpzU3vsJ7HaKyxJesbgUAtv0rW6ZqRAa7n0TU5ZEIAt+PriwGzEqww6CP3
ld3tcwxqZlK4iL6F3pPM9uc8v7Jr8shSog5jYaB/XZ6T6Y9ecYRANprisd/W1t3d1Prfx0IgR+pi
ZAAC2C00NCFKq0Rp0F2lglfTmCbgTHkwy4J3+rOtwX8GqN7kEPOBfOv8nlXsPwOn0WLqU7b281t9
1JkMdfaC/ujAIxDzc4QncqS22Yk5i2BcYHjQO3crIBypWvUg6aooB2io5Wy7kgJquO1vMzDOJPEe
3aN0fZxvIdYL3L7oxT6frW6mYD0MgaA88MrkitQohMzDQheMvI4AohyZkcMpp3Ni6X1TWScG7Cuk
j/djQRBmIcDx84baOJnBypq6OKakGD7TG8K5bkbITdq4agzEOgM/l0SFKFfJKmi6VzU37tZLrFKt
aDPBQRWirm0mmm8IvOVpzbqUKfdQ5msFVGmlePmYWmkInAP4wWEQ+s0WSXTbyO73HQn30J60ejdv
gmK0Ua8aCoQPj2OsXYEysgcqjGwF/bqxxxTitXv1NIBHxwhd6XC69TrJrANOId9XFnlj1Q+J6FSo
4OKFqRQK7ilINbOYkAR9RE/XkuopdQKIfx8BqFZlWtxYj3Ix8hpMUbThuvVqgBVmiy5f+2AignzS
pASY80uslz8kVbj9Rw8wGq2njYapnElxAW1yTQ5qGCQixTXVgeXVvPU/T8cksImuNJh8o4byIYWq
EqLMdyu+/FvBjCvBJOzkDwUUSdhz/TstOEifnyoXIR5hCY3h5jcbx7ozSOmtMa1ZVPDNrZfl8oMe
VKWt1OAxgJTbOmDMPfxjjN8jELtb1aoq9xKHEg9iMoSp9srbyaZCsuwLfDl2xFYLHltQ+WnG4qbh
2fcbYHz/Fl26LXLZzRQNmaJgEaWnMVMIHc6HGUSgRUFcFCjS2X3S/O2FU3Otu1dXpR2vZYmq0cz8
QAUuGvcw6FvGnYYejZOsQF4+qmEtm8Pj1iq4n0ZKauftvBLqP0z3TpWcNjt2zxS0qShcnXXCUoOO
xZ2iUm81LiEZHi5RDfs12VB+8RU0X/+i/XsHTSFsFYogHfB1Vot2Y9wRzVt/84pRUK0SJb2tOT35
HkhQMkz+fDewp0xVUq5U0NrxhEkfhgrZAzkp1qWrFFS5ZUVDCk9Py80f34QMM7XmVlG4hC2nimiw
WK0HvU/OAe3QWvGTziKyw193knBo2KeNte0qftCizlHd+uHMvcNQ/nbzvFKI8OIMlfjuEDnjyMSM
olucruiQojTrQlNdAwSbNIr5RIiEQacork7X5C9r3SIW1w/n3Rcs5+fxIB06OB+YzRIfJtqzEOjX
DlM5/r8TBcvA/WhK4/XDZjMWpSh9Jt/iP8xuBsPoaVDTJZrb+7k/Q7PwG8bJEZCGLnikVF4SQSOc
netn8l1KGQDP2q8QsBCCoD3XpGYc5Sbu2Fz/VP0HGutSQSxkf06Hx7DmIPVvgla17o4fLgBoSpwP
3KzYjqU9U2NJ1/EkBqr5vVPagd8rp0upr2wd+kWBBmqp365biUV7JgiEasvBIt88I24OOFB02986
DwDK+RwM0Nq50aDQtVymeE8XnsqreV5Q3Lpg/W6jZx4SIQibZuUOugdw9lEXnQuRPC1+i32ksCT0
EghsY8ZMtDCmz/OnEK3zDW9doy6sLbsVWAf5GpfTA15BA0UNGX5ZaPeltANYQaFsV1Jx5ZwHxHo3
LOT0ulaKpYEVI6RT/fCd3v/XkepPUYMOMYHYOog0ANfw4qHmHqU27t8cn7H8LKGe4YOMrOfg6waM
VzMLakk79trRQ/Ilh/2HEFth4dHNMuiJqTV2dwa0Lu8hPydzxQ/uFLbKneAeHqFKZNLsW0j6Qe/o
yVet0Ycaey+X5mR2F0ZyxROs/SykNN5nNraimDrvCgTvBqFGLJlR9QEPlbbBYgt7bkAktV/szQ/i
ED0pofU3TqPLdBghVg7eRlr9ktDSaRf6s/D1S5cY5Z/pZD3YNw0CZMrW8OM808kRPw5xWJXK5Csq
WFeKjqrVfzwmKRmyBMWO7KoLCv91FNn9MsObP/N5EIy6riRg+oDnLcL3i4SFclGaD03vUySOtI9D
bBcllFgU1+k/zLhGSpL3XG1fD8xYwwhgOenQ1q3MSHcXOpBWAV40m/syzQdH2LRtUlhFk1tL1cUn
9gKij5j7mlt0HoVWNQ5ihssqOq9tlENJRcH0UHyCu8FGyTxlHUNuAYWBw40PI2Fk4z+xGa8AET1Y
aFHba8XcyNOQC2XiGc+u39jnxZlhs6L3UDSHCDS/AKqhBVT3xnLlb71W9MeQD9/1/1beqCPs13hG
CSanwCEqgj2/2Rsd1SS3ZsE4ACqnnev9jPxiwHHwJyafrpthyIKROTRNTKInukvZ7Nu5w3LENFrN
+Hh4Iurg2nlHkpwF/8BvvlXw9msy072EM5rnMXa8SLn/gAgvv65UcSo79n4scz0YxK/rNmRwzfBP
xflHRMBPfDtx/e1FgtGSe8iGAZtbIzmi/br9KZCtwm84tV8trCBaRloGRepWP3c8v6/f6c/CEtKR
tyl6vstfftqGxF+RHqLqqfetkHtQxTmb+vm+64uKr9b8PqcPdK9xhBFx+BnWlHuLXyhnA2ubpazm
VXbq2hy0/T+L9tDRPZ9BtYU5+HtZujUnBnkGB3mZ+4EH6dgVqAepkWciAq9m+B1bsnxSOZaC9QQl
yxMTEMx0haiKIaAiq5BaZYMyRkdJD8kVP8ylF9WXPHzeOtKRXO4/Ru+t3CoIWQSdhziC9Bnz+r2n
D6y4gWlaJDWL8XlkMPP0MnxTgeln+9ubIR0o1DWwoUJy4yArtz/wgor7C1bsnMicIC+CuIWcQ2vV
NH60lCI0cKfn+ziwayT/muup2e7gpWpJMsiq3/v01KoY9SLqgTxubCUVPrxDMpKSloFQSysOe8GI
bDudGhw/JOHMwPfiggoCVXVgNXmm9F0Sl+gPwFkP8lCXRk7FWx5QWhNXaDlBSff466sQdW3R23lZ
eLgdvh850rvtrtdVhWj41WkF/mc+ahcse1mrBHgUXidTuIEzeNvwhGWb9KkSm2BGVBLyi1rPuVwe
3qVNwCOqL1vEUxKoqjXObbuykTSVGGgUufm8o+2r8a3rcQ11Gm8R6bjnWcE+yg/OzqmFdaj1Po4Y
7PwrbAULQohKA1XoYKP5n4sO1yVGeKg3bYT9176rFX8A5+YInZ445RD4BO0K8uQ0zZxj23CMQ+Ob
DZMT10gWikZQ2MJA/98azd9kjIathbGqJTNelDQFChlfRxNer2JNTHiJM0F7Hb56Tp/6NgEfYXVM
fknp5zozixdbPsnUbnWlfUv6TzIjumZk4XVGii1judmZRdsZXUGp0Gy5J3C0WwryrJ2FK4UjV0IE
GqFMaQTmYPLh3crS107FSwKEP0Tw/upWLdxX4VIVRe3Wwti8EuLVwAYBblNT5xNWQm+NVcYHOzwJ
0BcJLrkhYa6ol3F0j1eALcJdXLVpOLKd6FLxiOybhwd0tbX0XKdPQ1Ad5+S0yHh2ZEjUs6Prt+N8
jHAi/DUJWLWdU71zFti2vJqFf1DHUPNAuSTCh9ZRYlp7OeqtNl1nShStY51nEeYvRYSa7lPqgNXJ
8JjwAtY+tQMocWQkq+0pk4RzOIowFKyOZuovB0SQ3O9xV0YG/yenqKZ65E6EnobqPtP03A8QpbPQ
pMeuhHcPuzvXqXYE5rsE83Jw41+23+GslkF7iX3nKvy3h5LBIwZFmjLL4NjRglKqE6iETQQ72DLE
bVyspsup/EDZ7VPKqh6ndJmxJZr/mxWz8rzgW1kxmp3SoFfvQHH89OteBr+970DTWyWXNGUg/ZeD
DmuLkXuBbig2w7xqpZkFUHy9trd9/wq66N/IurEEzcFsTYsx+uCtWnM1noV4WxohW2qLchyfEC8F
YZZ+ebtbR+Vr12GDUpthcUb30E5hIJSjknhPj/3cdMcRwUyrSpook9tkiQQLi1Jffo3gS6PPvN2s
Bwdphiz/xVsmgNkTfKTHBFxqkOoBMkqJEP1h31rsxixN0LWVJ8KBKkzJPUq4Aio8dfCAxbq8miEt
Q+Gq2jZjZ5FrcTAoMxWoHOt72I+ppV8YlQ/7Ovgbk+dsyZ+kUx951/4XaXUM1CrBV3zkI6KaFtov
Y9dnuFWOpLF02GIO3sO5/vdRSwShi7x2jZw53ltSL88azY4+QjceHhLCNTrpHTA2Q9g92Wl+MBSn
nhehfrnHrCyMwrsiYECF0ofsYpwSCgGHTuqVLafUjjDgj/Dd5dvcDPSUX8703I32zB9KZWWi/5dX
bZ9KNIFY+OAq/r1UbkLZ5ITcepalhdX2i0wYD4g/a8BU5n2Ox+7NnqeXjPl4y1Dkwaiu3zuvzBr1
5WFnOjt9LswnIGNGVlFKQE4jsZ5ochZg3P2hvrgNfevzNvt56oPx99888E56W1t/PWeHHhc8DIzW
1MAd8+Xd8qZWDF6buySX0xudr+oRgquV4mfbVUDbdfOE5olipZqxPI6Sy5FIm88ti/XnJuq4Wa7L
BvexoXNJohGC3K4YOBJKJCFmSzCqJKo8W+X/CsMSg1lW2lbqC5HY2KQhYwwFeK5vj4wIG/drcptf
mzvqY5B9ZI2I5ncGnoFHgXmN05QiIkB8BsPnkilx2hHGDOmgeNx9BgTVIf47xcmejolq71MYeeWX
k6zLccVwdDyDjkN8T7PxY2aveoNIjcjFyoqm01zkjfHWl/pjXgg7iS7Bynz2RZYDKTaesIhGT5Xd
WinDeGRZlrrCunIyP9J4xznZ87uJE6mB3jvvSRSdvQyzRpijrPLm+8WsS4NqC0zyH25F8YYh+jDX
aTnqVV4DsTh2weF48BDHTEGOb8a3JndYSyc9qXTljYzsi0UzVTVT4Mx/RYmImt6Y4BZzaU1FiPCq
hOs0xpiGQF4vQQhy1M/gynTOAOqAgI/modFymFmLazeupep1mNl6MSJXS8LjcTtRr4CqlMWtDozG
6DfT9iOsJ+W3HiIcZczVbTAbx/IyeYLAzH7kqVn5nZgUn97W1X2cm4roskfYsWxEAUwJffwGbTj1
0LtM4ndRdB4mYN/ayahjzZNCqPqE2PQikaqMY3BoOLKf18v3WjDNmvWgrzaKJFo+BdiDsdL3yWRD
KzfurwDq7/Xk9zl6AVqyhWhrbPm7sViMK8k79wxYITb3HhhRw+IOtH9xFRL+RgqPlLrvlP91ipXa
rkc9kwpxrK5kH1uyIS910M2Sh+ZRP9PcMHgfL327fAcSSXI1h4teKSYqZeNXJIBc+QEb2yyFDwim
3nM+xMiLBpNnQ5eLOQd4/26OXUixODQI7LRa3I/ZKVJ3efCXENQGS22l+oDAtCVCX44noXSHaadl
0p7Y4i7aSj5+0FhstjljC0wlpzFxYSAeK/Ty+MEvUySrrZMUpG/184ZKJrK4DvntLYtT/iDW5sp0
5lsaE0FOiuasy7YslkXexBi+kB/mEzWhWsV5tSVZlHPJdGgW5KHOCd306309h8p5YbtwpvEL3OTR
zLoKvSt4yVz9ZvNAT0b+jk3ast2pub4XQ+bPoNKENEVsoETTIP/ePopB04GpMYZrAhyjpdX9wsWN
44QUEcmB3vRE83WeCfj+uBKVI20guPcMACk/UwJVAMcrScsH3VMowjijiinp2PsuZ89EOlgx8I8b
gglmtqRQAHEb5TntQsqMfCwHlChI4J904xIbYXGB0ykVWQYlTXosh3GObsOxU692Q33rfuGDe3+G
dAm0MO4CJk5EzLtbL/0KH3WVZ5uYWDrvFAChJDI+1FkEPZCWwkKXRrg3hkM3MCuflu+Xkf79ajq2
I73RVTnKOgFUXYf5vO8MbPnLLZpiXjZEu0y0u3cfm3UbShhGVaNfBHv24o2XxQK0ZxeE7IJtweZ0
U5voa79p392rZjbIpPC7l8FS0a0msOC5pRTj6Ic2MNPGJsdgiMVsUMtThDVnERSauzuwmDMO5Ej7
ePOFzrfWf1YUUquobI2nwRgljiJFyWl3vgWkHyw2kMctHjCVyyCNGSzkeCrBUOH1iUgIXcIWcpj2
3Ohbj23D/0JHJG0+Ls3SQXEoziWVEQIgnv/2JwHOEXYRgR9xiFL/QMIWUz+PCDTNDFl99g7VAul2
9k1VykHza3dUEJbaoQpFJJYepmvk/kz2ujIxPfhZ4ZEqi6c60KQ/xyvaFZLDIpEGJmJW2nkLtvpc
ibu1n8VpV5edUb0W8DsPWaEZzI/QwJvtFWyf1w+i6cO7OIlZZW2OARVd2/NFu95maz4uokr8HJ3X
02ycOvmEk6u11QiWRiFPvScRn0XwvVeedI9iseBBWrpZSqHmjPt8R0S9fMQ0MyzcXGvxSQ3T8Oej
K10X/2FucS/VePgjhY9JWeDXKHHm0uOomruj8RVyrHG5magxkpGO6hDbBn8vszb2TB+H2lDh2FIQ
qAKOgD5lE712gwAwi5GBClaGvNPhL7ZO+rWp42yGbdRougL4q3OK/GNaywjza5C8AFUeNDqn0dH6
4DAMQBiNAz45291hVZtWAIL7C0Y3WPMA1j+t2MKVGUMjwtVhnGHYUH9uDLunFO/jemNx4/GnlhkC
fugu9pJLaasE2sfFlm7z2C49bhJAcbYqWSl2oPd113IR5VUBPhzkg11siFP9ULpR3s24FKR+88xp
l/FR00eqB4YNYeCgkokyXZpjU6wzhdkw16bV+2VqbyYyOIU9UdBXoKbxmM2m2EvGNzikzQzjgq+H
4cWUyZp9PHl/a89a+tCxYmyKn8dRcubOWAuJCLs8qXmeZMB4VV1yWyOwMIaZFoirFi5cmbSpoGMD
F2nA8pLDvat2QkUMzIsTMQM0f2wo3bKIHiqvNHgxHCe/K9iciaZDhpi46eessCnmhlqwvUCPN/fK
+13bH0HxP6+o6z9y+XsrfsG/eyntPjHmrTufIeMx47lZpVUOP5/yAqhXFhll74ULO/KYsw/hjnlA
giUOUgqpha3X0jXA3gmOIP3IOwGvJUwqVvKMO5hK+PrqMVF2u0KXJIwWQb9manLG0yhdsC1nSbs1
ikRvO485Y/By6QG8mkc+3U3sygclKzXNVktpex6ecir2QBblLUYaLIYuaKmtDDlzINvOxwjx9xnZ
1jvJVrSfjpnEYna9ka0HaX1037g9dDbS6L016Y6ANt/vl6wnyoTN0p1WVWW/I1hxnaTmEuBHAov9
b5C0EtXjL6NBqLMC23W21nsWfCEDK/hBqtVV/SNjm4q6E92yYzhnCDmWhl3dHjlXNXcF7ibJt9gT
VR7MkYx14O7NxxLx5ooFS8k17KwCIIOjNn/tkZD5sTArh7Z9U3a8kV6MhXZqdI2qD7WT2GKpOXLG
cEf23DzISf00pz41tsJIUtpX3xA6gXScOfbC8cxsR/zFyQYwroXq9TPUUn7Bkat5GvhpSD5mY5oT
EFpBGMVGKUlReTbBKym20g3sEV0W6XiSNSbn2kp076Ajn4qK0JI8vpGJcXu9oXz+/BBsnkT8NAqE
zl2O6RO926rNaIykNM3it5hcoct+6Gdn42zjw2wY3KCYm1YJA2CVDwQJnwSM5BYrBxoxnjs9tL7z
8FqvsJi0F/fMdSODnvxAvdZ92ZpwY3+G3m6ZwjhMdd9/uU8M4LQudjO+WRcNEl1DoK06/21B63wn
xR+38qKxphgCN9f2cDRgfyZERvRKU9qnsKseN+dLshIMYTTfqeRM6DUIACZFN6r+NukYuxuFhxX2
1QU2l7iJeB455fBJsKVT52GNmKdOqbUEsCjkDvQ5cBSipDeuaxgl/ECZvSgPk6gOWxImqtrq+oRi
XIH45nAXDKyZGitkGdpRk4BFfRvLtRc8Z3bKwqlnHHnjg95+p3wkuNF3uftFPGaZvawO5hjWqa/a
ZAjq8af9KvtJ9I8g0zUEQ2JR2jqT8Nfh3n1hREjvMcv8c5QWrQMTV8b4Sm3jEwbQU7ujexEH4/e2
aV0LueW5Km+8ZZOskyPsIq2hhCmQ6O4fMWduo4CVrVQfbjd0K9Y/XHC+JfsX3cdKwT/2WdLevJiC
dXEg+B1tGOlqE5UGXsOZl/thym4XOIbW/D4wNLc42vfcwn+zy8f2Xn7XLitOpn7WAVFH43UhfgkU
yQRNrUVhYkFlA9uWf1/cOBewrQxuzx/s2caUVsL9e7Ib4GVL/DGCwukvfBS4KJeO2cDThUTjS1aE
up0RBD3o70277xIr2zO7u4OQjWDJrYjcQCuN/CbLJEDw6QgzPEFrip6f/vDJH0hHOMgfqpRXALbj
U7lCrqwDZcmK5AgfmFkU7kZ5zSn9YExFVnJ88Wgt5hD47XlOwkMf0DtzGOTeHLc+LF9S3X77p5cr
x57R19qnFGPAjdYSqFaukwCMLvuq0/Tvfw6zAhTbVOGxuG+7MQ/t6iPL+FZTvIPsIWydFtXrJVnz
kU0nKk20DwcwhAEusEE5Xtr3iw2mcK+IGHFChKVdc6MVhazI4NH2UMVKWeJ2kCLsuFv1m+yQV4OZ
CNDL0RomZnhYkORz5965sLWSX7iTCknDVPf9w6GdC9k2u0UNPQXn5779D4eRwolKJKEeN49m2LZt
eDRs923qb/r0X+TwTctMiu1fe1pS8R6uCdoO17Y7rmBmjsnk8hywJ42sKDnGEYgL7N5buY6uRn02
99Ce+MCvA0PmiyFooLi0RQlPlFVTILqdl9qObks2tBfjb2q4hYOtbIRI9oyB5DLGxIiK/hiJqxBh
pbzVqAsrIF0HUV3kowmfaDdI2y6o2AlUeAJmgyh49koP6Lm2RpX/8d4iKPV61BjOV/BQzvtKkxNX
ugPUcesOyxjgh9kUAeQ+IW5rO3Kitgu8nTzv8bQDhS8dCVkInTZSzbho9d1/l76Y3nsfaAKWYSy0
ULw4z8SFhOMlRFfNlQ0nAH25AhfDnpjdLBn9xWwxXag+1OgIAK+TZA/XgWzb1XKj1xLjjm6cgnwu
MGQPuGg8q8frJjJ4pPZ3BMFTWG4XnVaZrQl+F4JDk6qVFAA7+2ai+yyVZv+dkhXRcuXk4YE/UwYg
uEIBZ4uzjb5YPEyxMdSxzkOG8FE7YeZcXuYo4DaBjxHMXR6hwaIV+AKVWxPpf9432rd4MKy3xOyJ
Vle5Lg7+KJbKDCJnYmRCallbMb5njsKAR11c8GobzKw/7shOkqNTz+JAIBle5ijAStjszOEL19oG
g9COOuTiZZWFIUVlr/fZUzTiQtf87LoXxiCaImuyd6UPj8+HNl/l5NjplUTpRmFpt1FlnpQ4p80c
i1vE39ucIrh9OpF4zOqbTVbsK0LKD98g92z5WDYJReh5GR1R0gaYmxqpV9CosgT7nCscmqDAWtXp
pSLmaN38RkGeSBSKuhL8azzAB0AS2IrCQlpCw8mozjSHlPGETDVcKMs+QBZqgYhNv/FWkplpwT4d
HHmfBtq1cAOeOdnSO4AZOZ/W+nyPirlRWN2lizU8+MH/UMEfS7T8OiGQ2MOZvjT4VwVtrB7y0wdK
0OnONnG8OvEkbPoZDt4dpM/ecfr7r4qTyEFvPehdNsydw03Hsb2/4ckflqv06W0xoTKgPfQN7DeK
Z4T85HoXDLPvb5Do/AMTALRBips3iVXxD1NzP8XCc62O2rDJlevgtgmsx+DBJmyAgFxog45mRIZO
27niflHEGP3cbY8dqIMTYlUPeOjWGt4eccjCqFyzCUxYalNj6nQirGzwybCXDwBY5TTx8ZdIuE+U
5ABsXJhnj5j5THoy6ZiIgbN7SbvoDcZFi/HYsZViUbDrwDhREkJpcSWrSE/jfic7QQBUxHHokQ/h
NmjxhbexSIx4Bu+U2IF1EoEu/xiJFht8dHXmeUQm24gKux5Pde9TUFxGlLvHwlZTpEZwRX0jkoNA
SsJQZ06P1F3ySq4NgFKw1PJdWgJSyCb1OX4lp0VwyoLm11ZsC9r44nHigGyZ3aaq66cHscRG9sQg
EE963tQYZiv/HwE/qSorZCDhQwWqscjyhmg/XgApLo35fRvmCba8qKyPKbiMcNjjYfgTMlZryjVJ
xBrzVZyca2/BA3z31gwlxI2+P40c8Ea05dMwr1LIOUKYCAdkqsKH2QM5AEL8UoQX6yJRJGq3otkt
ZbQFWfb+d4Z6Q55jpFn2L84t8K6jWnEMhK6XKyp3AAn6VY+eG/iRMyeOy8Bc7Cv5q3hTj/qDfuKV
sPbRWoranE0dbT/oNJfjXlmo4UCbltiO9R2TeizmTjaBNCPMPLq4PRAY6yxWRzYT5eLdGBwxDerx
AjWhTaW7brxxSZvyEcD1GbDY1SobWQzftfyQeoCCKfUOuHUPBgORRrllfl+EA/isQewiFFjLDjYG
ENZBd9Je17oPEvbKW5sBYtcbV2aODPQDpy3F6QfFP8A4zmiFY0r+xZcaUnuYriYvHqm3pQtWWTEa
5MfxXaA0LosqJaoqFKWYzq2DDoLqT3qfO4ik/CQdiJH5p6BK0+6e554+jP1CHlfDVCv8F7l0Ctef
0OTrvB6zlvl1Pi2wce2Q3m6qXMGCqxzvSajDPlE2qEVTOupGND2s17dz6bag2+FdT5SOGyieml18
+BptVb/OM0GXp85IuWhD9zzM82R4EKRFBARC7Qksy7XciuneteGlRwkLz7zsNN0n4RXAqstmffhw
gMDH+kxKywBef0M/inHjMbStmjJrCnQFUZYbO7bvdJGeIEtGQkRE2d0R29EXIafdXQSUSgUVVNlm
kW9BA65Ipu2TG9Y7Pgrf1xB/P7hrcecR28NAqUTqWcnZSN9szQmDLA3340ACASIpUcG+QIrMuCN5
Q4YeBH/H8fRjYd+oULTsayylxBHwp1mS18nSCrlDXY3NFLLonbgEMrhhN9ErL4WviM8A0JfEIb8h
jbO5sYaaHX40Rm8WhUW0HCyDcZFvSaDuQEZmMyfBnmq2sHvc7C4DAbVZl4lwWW04BNek9j6+TcCd
wgel7JYfdt+HWbwW7DxExwl19WoCOWDA4saFr3We1eHYRReWnzjXOteEEQ7WjFSZAp5ltjeKKKAa
RnVLsjNRWxatx/dlyy8RBPSVOwiU/vvb7ez5nZBjbLCDJ1rw5+W8OJ1IjMNk5ATQd5ui7SdXSM1Z
Upy8fJ5ZfYJlSu9t5OO4wYqaA8lhrMR1Ya7FdDU9MvApBQSLgEbySUBjFdwsO7cBahxFuGpKiSLE
omst4p3Uww8O46cNnDLq8jk0mZMOG9hTD5J17yUkg3M3T+ASIuGOgATTPwLPjN5T7JRSWEUC9Mnr
AQ8z3YjxTLAyoDlmkgnt38x7YhRqOqf2cig3KmsI0zMykFnv4bLQnXiKV3jOQoCPV5uKAkOIlI3e
Ul7Bf074pl4hBQ7+xYCkA2AHS7mC4Q7mmEVL0TxGtAUbpEFwohtiVBhUv5Oz20cwv8fvJyPzvXpl
VqdGfh6xKtfiQlvjXOVbARN586ldjPYarNxJFqRZCN0PxR19JvT74u2EzuKsXVfZq1VeSg3+Y+LV
ivaBYadEnJK8UHQDvBDCE/Y95BEBo63ON+59ZNOX8RR23yptUjKaA+KVKZvN+jpQmdVB+Px6BPiP
Rc7lfS0it8YZHbno8wdyIvK+ZvbtozVBvn9lg6dKyYwXcC3JQrxobfrNlg6G/4uhrwjgWzw/UPlA
xDNU2D3p8n8lbrQSZD/bNXnrP/8a2jQ2IoWQHx9RdZBfFxmlqMcnY7ghgqdaDzHvkPRzXMfzjH5Y
Gr2j3JBLbkeiZV0/VMzSTpdDnwHr5MCuJaNNhSd5GhCwkuauJsTAdm4Q+jEb88F1X9X4VeCRAhbD
CLk5giJv8lJ0Z6eAC90fwpAcgm1DmPAvzAnTfn21oCC83TPNAI9AV3IRV8XR0Z1DYG3qxjQbTg17
aVNYvvGdNuZpAubsA4vB079KZwqLzsYLb/4Wt15iEdhn0DuF0hnQ0gvlPkpi5nvEe6s0t65ToIcb
LE8PoKeyd1R/ASXEx0GRpM6EugOq1Al/kJl/52PFuQ4m7uB7eqwAP3sfUmyxLclugP63khk5kkI6
Bm5cIRqj91/N50UGk98Gv08uGjo7bZVFMlDRMOPt6geKtViB1k0MAOijNLrOqz/9swAeqm/7zmMw
lwX75EkE2VPzQU/h/l2bwSOQYvQ/x9JwrGJYtdn8q0GRlz7QWlb/QWkqg3v/v4q5XD2ZntiLQIkV
ceDCqwu621vRGFIilTwlZ9lF9AHh8MCa/W+RR73xHaB3emeQzyLcxSO6t30wQNcRqUiF6uH1CS/8
vqDUqg0RySk7Sd1viZcQl7226vSpSuGVIF4KkqIQv/LlqsDvSdMXE2IORO70bW413kMXrQoYOYQJ
ta/7JqASOVNzvSiCp8uW8CcGt6S0KFi9ritT6ibhxae0TXvDhJQaiXit2oqEIdqHQP/H4RbI2cFf
Xw73tnKTVmJY0f2rHWkQrILCoOZCUxTc67yaayoAWn/Bnfpb2Z+4WFFg+T77/Wkw7q0O7WDMNeDY
Jg/Ipvv4q7dB/GOfwrk5iRt5au8/3/OTxCEMOgf5lTIMt6FcKLhLmTEslW893QdKXbN/ag0JFCv8
67Euw5Hm4Pqt4hJUKHVRmzAqubWE1AfSwOAS15kwS/gORlO2opVz8V55tRuLh3Zh1D/u9EwUXyrw
8DC13NQU31z/wiDajFU9H6Glq9TO1uOMq/XZwkIb9Wf5A+agGjBOFXuXdA6EDSw+2RHVdDDSJA9k
orlEaNjunxyi3rqkTAC5pT9mXxxL5eGUZMVJS+Ebc7PoTGeOsTqu8R1GfW020UdXGHRXmCUDa/lm
fPiZnLjLT7P3njrlx/MeAorzsVN8jfDXApNHwkeqg9r99p7SgiFFt3wSPdNruBbNwaDcmWY7g+y2
bgRIa/5Zp6gYVoeOJYk2q1X/JRXDLyaTAY48ReG1R+Ngi/l7LaIDiIdW7x5JSKmFmY7uvyfsSnO9
IB0UQ5OfHdyRHo/205GzuyDjsaK7boI27/9de1OlxZu5uCaLLSeHbztBQMnSYrCsPob1kHO27y9K
WJ9MTprgMvGWz0a6aa+N5F7yToePLGeY1nDcdWBHqP023DJNb5wGfUxN/2cdFCKGRux7lzsZBtQ2
XmLVON9brfNpIIu1FLha3q+ts+RR+cUpvlu3hxKAjzB2cJRRCjMKNaxYjVyQOC+32b39PVME78L9
0vsqBbgAUIpl9O90LrDhKnSXo0Fnb42VDPY6bfu41E37lR61rP6LvQvAAZb3eNwi4XBgfW7P9VWC
PE8sSwvl81D195P0IFwiRUR6ORVbSF8QKh4TqaEklrc/firrfXnip/U7Rjn5Nyq5CrjVOowCYO3l
dvTIrmRLqIIg8oGmIbBs4kACor6BDYrYSDUXy9bREnqQ/qzkXQWQ4DhJh6HsavO3Nnhe+1xn4I+5
MLwh6LJHtHZkK1kNoaVAYL+DsODOc3vIKJB8p3KsxTHKpsZnG6Ls6x0n7YHdBG/UzxcVLoq7O3tF
LbcyA3lu5HEZHgK19v9kfmmPNc/E0jC1PLB+F97b3TUFYhR/FWKlFL2XyFVN6abfnFV1dhv3tiNZ
HrN/7MCPK02YCcySnYtxVYLvgrLVvC0P43+XDW0Drnsb4E7EfmHx1EF0oWNiXyrf8h4czUHHi6FV
a+43GUP7PfHvdROEobj6e+bmbDEWVOC18d/7Dh0VfXfgAUI3nbV0LqDNDTa5YNgYnGRBrS6lXZGb
rR+XnUBKhH6GsLb6ks/G8RyTr9o0zitrz7EEGeA3i/O9mFvhbMiJd2BPt+npIU6DN5PRhqFDWRgM
4ecbsr+xQLcBdNradIsLMJ/bbhmd0BRDwWSoSneHedN9Wqx+4r8BZWx54I8ZZEpnqS32cJdDWmVK
+xxr8Fp8Ih/Gpp9lcLWKKNLrhKuNqLoFPW228P5CHbBrHW5tIeAKN9CXt46Hyykyx6j0BJb7+jQN
duVmrGlSsN8vYrjK03R4TrULTmwEN+0NLFe3NEofO86QakxxK9tIZGBUVIwJ0kmdb/2bDePZ+puS
de8z6f4xHH/TQlf6kgdn2t+a83ZqgItObToxC8+/s7HtaqO1bLj4JUVAmi60BxiCPOZs219vrFD/
28BdN3SnM3qa9tCfP8bOEavDjk305xsfifMO13lgQtRL2Sd47pyvhHb6z8COesQTzHFoY2z8yryM
vVI7rNcrnK7OvUVGQoelPtVCJch1ZIij2pNQ9wKXMfG2YkHjlmsS3e8O9Alz8KFSSp/uedtq3kOe
jj6wB0RghHA96ufTO7QSf2P6SMMPakhYPGYZsFJbXRYEb4lg2yox0l5qiITBdIabFGxIpAMNjR6L
T//f1oqC0TZSyVL1wK3wrAqnaBBZrcnKi5PbPz1YXlfwJgpJ+OCwwagugARTzdTu+wrtAyvh9q6R
ERLsORsajLj26wYC7eWkR/VwRlF0BRJ32s+47x1yZjdZf77WlKQKQcAvqE1zFe2G1Rk0v/ftGHb7
MLRSFcIM+uWvieKfK+FY5DRe978U9afO1zHyAp7F96hGk+g5wM1BHg28Y9TXZQuykLOXGjgqVt2M
Q+33KwX64qTIu8Ns0jipvt0SGGtKheE0alXoOITQmGf0a9udcA/PHJNqyNU94WFMmAbnFGlACTC8
JLOrGskZIUtI6q0sHhrDfUeJJ2Lo+dWQ/QqW43g3J9ZcbhgT97TdVH5HQFR1z4a57V5Fhr3RZTjo
80iAZECnJsQxumgTGJhgniSfI5WAe3WTm7BdQRhbivj77O5zxlhn1Y5kGOfudAK+XN4cYKFo4JDW
FyL8VkAV/zM45MVpTjLW8t8/VlH2anyHY02Uly2LGci19u2bFjfLwmkGtHM972YxBfFbbDWl/o8m
FkXZoqHEHg7MXOxQsjeNoHQ9gyrgC7nd2AfrBmoCwxG2UbEZiqH1++WM1EeBI8EVq7P36n64+/e8
Lhemh5QhNvkNhgQ+FW624B/AtZljqWCyhJ7YGYdXmyphuvLzA9BSQ6qX84LJ4lt4H8PLYW2Kuiik
JC24f2Zv4v5LxaaJJMS8F94Ipyu/s8uNMV2hjttJT2V8jEJzTTYKpD73AaMOpjOrE1K/luUeYIT6
nC43yNYteHorkgqHrHbtE9a8V28Hrhx+R/W5T4oaPuTG/Gsb/T+mcOEnp4DzujG6bfk0D0oOSyWB
ZYraLvaeURCds0ifxUEVWn+HA81VMxzBV0uGLRG3uoaZPpASR9ceiAz9DJaJfGksNamxmxYp/CyI
dv0oMOlvajX9kayr8ulqCiPWKl238b5RC3Lzsrm0rMfNhlrPOFHH0kMhTEqNbFdTCg5sPiM7/Xzh
px7lxlF8nwp2Y+BHzD1UcH79rfsLa0BdeiVVYJDqqRRimZV2BqP93MAYjJKept3YnOVowL4LnD4u
FCsWTIN3E6MlJvLojGBn+1FsdoTnm5fYXuX6xWk0fA0hP2Q2za4yvbQHYQatu/5mlbmqT4zrS1xl
NFy0aY71weCsnBlF0Ka8/F5Z/nQN+8a+yskOl633gHvVBRotSpU2P/kHP0K7KzDfCzcd9IEnaSb7
Je9SozuqJesjoNE/61o8mIch3slcJFUQVhYVrd2MSFYLQmuvM0NQOSzSAdc/ERnbXu6ZNDuJlb2y
//ADEnLrry7SE7SJKFZ0de6X6Qcho1YvgRw4MyTEDqeEyn0u5U9UdmgyNuxJprzOeFp+ttsWpalG
jKeQOkgnLAfNEaItds/yRgAj9K+W6+A2DG42gqCFoMl3IHWaQzZpYp7LA8fb7hBKdY2V00HlQVAX
1CaakuNTvZH3fCe4ZpJAGKsDrDczzPQKzPz4zNuXqhOWawFui03P6pVaeQORE5iGRKrD/Jj4L1rm
AtU979JYBfEOOBiPVHZzrkuNi4XMMBj+rTZoOhV0eqQd6vqm4wVbzGyJ6f7KU4nk6+7bEqi4B8N7
E5N9KPTNQuGY31K3zMxFz3Ty+U4u33/gr5QlYQspia8aGB1cOq+mTg9RqjBnLAFXsfwsoHdS3A9U
DfmT03xOQ52U6qy6O7gSgbSFtyBu5ZrU40+RRe3EiRxIIzMIVD+UA1PXmOFk/dXPeLvNuqpbX91m
i4hKiEURKHBJzrRxJoM/kn2Os7vkUyFJ0a5uxUSOebYRWDbaAgNzLFz+5Rl5Q3taK6bTRQVJcnfR
rdPz+dfK33EchqJ2xXEsMvX2Bl7S/CAnLh2TZ2q6n00SMm6HXSQ9kmjrs5V7aYYXN0lN9qeRpSCz
3gkzwyx/qMGQkzyE+IBx8wQ/otAQ9+hxJ29SZLpHRq+ab5v1X0aLMXu8IWo3RkELN/l5fJS8cAhB
xM/Voc3AnkACOZTEacFVmyECGMXMLx9SwOSgU/GVTMynIbzx1L0WM+by6+nGKVMc6GnRrImHRdnW
bz23ErklIhKpiVM0QUC5JY4E+IPEvS3NXka60/vUk+z37lYsoQnqRVHeAGF7xzpRXMhbMR/blPfd
oTyVMxXm7tQ0neK8J/XBrWejOyPi8fBrJsTVg0YdP4oElQAVSEXBgZhEOxyDMg9SGSTdHJRWB2cn
RUawJWYotMvm367nAYyn/qFUmZGsTFNrsF+2Q03fxwRTHFEvv66sd+0KAF+UaBMPlT+odH1Zb9bP
6EouCt/bkIEfPEf7lYiYD7wKZRqN/u4SRXQX81ov1MDW4WVBMNKBD624TXdZQjpYkNqj5hy315cg
hR++hHL61V9w4eeHM4Sdr5h4EIUnxcY6uxS6Pp0RlDr65rxa7bYAntlaA5su9XrWhT6jWzjWN4dP
4NhwjNIbRLtQpvhAZTXFs4AFz20o7DVmO5Qgw9sAXESlmqii62jAGXw7kPiG7NlbKQfNE3BwwgNP
qIk5XnLbt1cxvLkFC8y8hyQcFnztC/Y/Bf8xTvDavakfem3OPiEU59LYi7EYMFHev5UK1Ue83b3+
f+NG+r79hVn8DExBf18AYSYu3BHQVwo8G7uGA9eUA/aIPVxXP44M5GKUbfKfNsfIHq+eKQylLvGv
X7UFfGy+sxzkqJbokz5dj8KUj28nwECSIeIjpiHbbHEOqwN3pYj5OQnkXatsgNGhDvqvPtzJgPqV
7oPvECiUmdsOig9Uxz42LksGKjGNNbQURUKsbvAaYmdNTMiRTaf2RnZfs0RXqaM85IWf1plH3UJF
o88afRSWabH7EGUtSyJaNavGLe9GMrOeaHSp3okZwDmuDCMEDaSWoVD9Ev+QwLut9NNa1msezCyb
aIzi0vlyd3tr1GG5uTC6oWIIjxDGfVfVpp8fWglWN+LycNnrRlt1OWpuvpswdvEdq1Laj5bFY8zZ
U7OkxreOONYZlHF4uzCqPXG9yYG+0/KC1Vgk1Zmhw0Z5Kgb+KZS8hvhNqKT3GHRrTcCgQdcAw9bb
GN8xqPnlRP3jXhDYYsES7U+nmnDqj+274DrcEoVXlkEigVAA6y3ibi37A9CJdfut/LfXFdJ106/0
r5JoE05JGrnJGt1XGcmkwuKtnNxtWfcBV36yFmGGWww68SIFWZXo8C5rrFvyT08K5Bg7gjFdN7ww
iLeSc5+1bgVPxNgY2pvFm1YOkA7ws2iTI1mNLgbIWHHoDezwkb5NcV1O5lmBzvYgSQbGqqLPJlYU
VnojvrGEw0qvs2p1R5Iefjr0tMWO5q0tLVbLnVnHkwnFm+SmwT9RIiNsUvsF4gU7iYps4aVGGYBS
eB7xFbYYmFh4/xakBnNBrlZ8L9sRuF/2RhCeQWvfgIbVy2FJmV/6p5gU+I3tTG9HLgnuEcdjK9h5
+2UPATil91ceknr3Sy1cP8EvuITvpJJMATjCG/iCNY0KK4Fe8h4CNXWyFPLtFI6Osm/bP9VPM9wG
ze7w2a7/gTRonBLrZWs96QrNula/rLks+5sJi9/kKCKvRnQCeuglxgMKaS+/0toZ1wMVX49xO/XK
CTMlE+YFZTc3yXBLhyGIPBiKn+w+NBgkukHgtSvpuVYQKDAvoSzItmkz8lPHeFv3eY6DYDslP7uj
ujLQ2ahTUfpBfEHyLxIxlejxp6dS0vorAV/YWaKw/aED33u1uaVJR+bibjQWJuiNnpfJ01Eib9qy
XZZ0Rt/J2r0lxmGVyEZnPR/k4PdD2WAh8jV3ykSQC+o4Edj5stBMJCzfutVob+GK2cjPkJEcSwjQ
DhWxtb/ZzO2u4DBH8tWv24QqdT1WXbDK3yD45UhUrovv7E3QamDR3uDvJyOOZMbfqt6Clexkm/oa
hK2+KYKbtYQklOm8xZGNkqZkvpSNJrFBMZrcNLDwed4mKDA40q0lovfMdmbvdu7lXsLL+3L95C0c
eOheLI5CdTswKpXKpsJRpLw43BzvDpgZxSbdFcaVEDdrYBeN/EMzp8JFLpUkgZ6MIuQNMilTPqpD
LPN2A3eAOYrmppAlP9VGoDjsUH44EYezIvhZ5wE29HmBFsgYUl/O81pgETjATOszVTyvcl3nwR49
KMIvNi1qCEM0W9GiyVkBCPidvzgkq38kAL5FpkSXexkWbBJ3RSTWru/UIO0E1/F9XK45BJ3dtrMk
KxmKlibxiOffxe18g2vSPM9lIO0lATurbcvFABoqqFnIweSCDahsHKdOFmdUlacmgyEAtoSVUugg
KNJkT2cLqBvBum81ikxq8pfmtEYzQK3syNog3J2aMsIO7gc8zgP3UkWTNRPOY3t7pF6qxTVaNYOH
C8kfKMzYTmeh7BjtMEyFG5RyfTHq3CxKo9tZdvlXCmjQGDwGOturo0s5W3fEuFVYLNH0QcYSRSqK
lDVfUTFFhgFz6ozR0oVtN2S4E/O5jdmPa1Vblz84c7gOYMOLtmd4H11cURkemUF1KA2YRGk6gs7W
HoEl+AVDn314M6fF2lEw1UvLQLJwOT1PtxcyfUhXibAyH9ciWihxYdiUVs7sdhhPtQor7PG4muww
Z3nnHbPuRIPvqCXEKV3Q6CXUVGxixObT4rlA0xFSMk3jcXxvoEfvtOkUstaFzHwtLY+uXcHoFfbp
RwxczyuUQt0FA7BgdP3g4M2EDHHusKvTow2CiZeQJUTYBQKPAw5aO4ZBDxQSwrpivMND8F+1mEDX
hxUxk+0rMPZx/+vM5QSPDZwlgm+FPQos763lCWhFXZBrCYkRA6YfShY6TGBl3DUl4JfGrxrcxtuN
xQ/Ff8T4q3lFycnr6BzILt7OKY+iQCTtyZOG5Y7aFlahNSN5x8MKVXVW9y4uA0LoQ40a3RgQtHH6
0sX2YFFV+5CQPSM16b2aYYLZMeXyf6Fw7UyiytCn5fG/BS2AHAGsjeRTDB2Nx+Ex59y+kFGh5YHX
oI4oSyecSiGwKjk9IJ+j0hhWg2c82fqZVl20RwbOZZy3ZFGLPtwSZTonoNqON+IMAe71v8lABHu6
pRgPYXm030XTZkuSlZ3id8r+X+ArMvW00X7WLKYpYVDgkDIhvYCUehlNeElVtBZ+C0m36veuG4DS
3ikO5tOaAGeo5ITuFgO8E6KfnOrxnPEHbBj6He8SXoEVFdflt/QwrXsA+YnLA9RKHzXQ2byNRmMy
FVcepIT2c/0D2kTdVQVcH5alFeq7cupWIW/gIer2sv/CuqOE6oPsyMGajxim+3+g2zSXj7bEndd6
ycfjR4kidB8Wv6BwMyNFQ9gdb9O4lruOH5zJqGzQ8l94Pv3WF6fmQYZHk2VvrbN9su6I7/8WUWrQ
m124BrWofQ/bFwdg/KelV89d01lKe6wuIHfnWJa6pUVdTSJqMfmBUt5JEMeaTHUQM171jWz+PIKv
Cy252dBlR2wIBK8DWboFrVsXzxBztCo6sVVRFnYgqfzlwT8RmBPCBt/6aN9joIVKskUEhSjG5YXh
U2JEDE/xwT2iY9GBGCrxQrAkqshubgvXvqIZUUEEAaEfOzYZDH2sKDzRP4xHMVAlN9uKwTadmRbA
nkATNIFnkhKU0qdNZrZW+SocWwTl9yIk8sCfKQmU2KEzMEIVhJ/4eGG54zMlG/QSJ8BgNUjGHrst
9jyBmHNCMFW1JMaANHyGK9p4HL/Bdd0PC4R/0qHusfrFYPGZpV+6pNj/eZpw2jsNyhSD9pzbQplD
CxoS7eTolCjhDaEAGUwxrSD/RUZ6fPmfNdRsBU3goerRmMOFBGI0o7TjDHoracbIqwknNjuHlHMM
aDQR8ESKp7BLKXzWddC2p9kWfLhoiU3oBVXbCmNxKBRtPq4F3hUtSp9nbydOGc39dN0HsNGTZ4Vl
E9r+6LMwW9rnO4AqZ4XuMDqQ3AEqMGbcPfnpJBqwQ7aOOuwlUOQu9mOUIJF9hI8ZUYe26RBc+RUk
Jz/hjkgHjkTkx08uCHOw8Epos9lcLwkzWksUWVZ5jC1PJfkhCpcRM6lxg7mIyEAhQFIJ3k4PCu5e
PkcEaZuKWqZMtD8dMRgovrNjJgLqMgXzgTZboLh1qKp/dOwlDPilQ6/mhhDUmaIuV/F9ky9x7V+U
hf5kJjzmpiTOOjM32bS67CxFMAPEXd8WroB2rXDoJrfUHx3qJa4FGokHt+XdlYVNTyevhlnezhXa
Y6aixAa/bbRxeTy0BiebNxEg7TSrX8lNlbR9OWdv0E2kd93VxuLcWiY7ho1MmBHLQUQvqiYwJKDx
OW4FyYXLwntleZs1X5XG/O4bQmPI9Qr3HEevLJn/3SwtJ0AyeHsdlU311fEhS+6tDRyiiHH3YXNI
ni2R/Jy71jzbFiEvwNNd+VrhDcrL1Co9ax9PfE0x3YJQb21SRYXldqXmxbjbi5RTT/kF2bIotToH
BiuIxUjr/PSQH6tSs7tCQjw/LIrAF5SZmvl1hm6fQqkJCrVvGDrdLrIssMEYanHgI2xC4DWKjPIn
tOeD44GYHuy6lEGpi65v6GFCQ63laCwGmP4DBzw3Jru4to6qS6frq0G0pqT3i+hrJLiRemc0yrDh
ZWysG0v/9/Rd66o/wNwMsOGSVX3fPt1QBtuYOwCJqTbGDNmyzTwb0q/id2GKAy/Zn0xWzKv53gnj
DMOaXC3pcH9IuyoH/xslFw1xTHioDx3sHYrxq6iD/6//djTR1XW8tmEyhPAXPsEf0U6CgOdVlqvD
YB3W3zIGA8W2L5cS5GV72EUvJRXHnOyQ5S4ilA+ML4yNTQxrYyjBqu5I6QGZGVltJ1823XitqJwt
/OsG8UNWKyc64S4XtuvPvptREWl+8sMohtmIKETHBtSXbwZuuIE7LZjH04hUAF2zTqrzezo0wvER
bdp49T8nbnxFK2Cmr4+7Xb4NF/rBrfLeZZWlOPylpP/6ciYFEEXlc4kJ9GoeGpxwTZ3YMLpy9IBa
TIIMx/rnT2J2lT+FqpGalB98u/779B2XQ3x7pUTTQvyzk/TcrwwrKNsY3iVlcQNv5Nwa4bAZPgbi
jGSC37RFA2h4gmL/KCo31yyKLjn+Oe7gAiZOMkiokZ9v34hXLuBojCkPf1D3ERvxAQNp7dV1Hilf
jMgTIJrnGm0BpupHzItK52gX/TgllrUbaKfW2k/9g75CFKfep09SNoIvnCsGF3RexrzeesGM82h9
x/S8nMtSB9rBosodAd/SF2pBIVHHm23mqKx6lFYmKwGuXE5pBa1L2Hv2rJZuPdVTY8FJU9pZ1Rrs
2RdnpOi6bLm2wQYubUdYQKYBqEWqr0ENV9fMmmAAhje14es5SUQibobfCNgythpXi2uSg3D6CkxX
JFTtD9uEsuEfZak3g5Y4z/0mrNiDKexevNVbNr6Pan4/90JZbv7/FQ8UuCqH5HkyTAjJDL8hw9E6
/LMJn/8pJ9qcXVqOeg2zMaI/ttGlS+cxSjQtxaQSrT3E964CFweEqZhq2OYOaNo7nX9N3qDevOqF
+oJhHnGoCTcgl9r/RhJO8Qhsvm7/0JRI6z+bnOJqoyXztgzi1YhDKTz9B8uYdOsUG90uTHgucsro
BMjJeDTOowJNO5qwZ718gnN5X9kUa5W8t1NG7P7gzw/MTocZKrE9Oa8dNXBWGqzHuJlR8LelczEL
2FHRAE63UMhahkq6/2R+2mKlnuV1NWAUt5K988F0pHVIa+QYCBAbfNv86CkQwK/JUn8M+4hQAPoi
UPwVvenJjdf1v0pEIpgZNDQ/cBhV4zsjH2RhfH3Z6WRDJXkv95T4qsU5Dh3Ra1uKEPZgCtHusmOX
6E73wu40ZCWv74DWvV7gRE8/DCc+umzaJjnL5dHwIkYkdzR46gBd5g8vU3HhnrmuP8DYWDY+AIRJ
OgAwas1mCxwHS6ghjSELqytLl8i8iAB8pRiarDNQLHVzlDpSWl3V5OisSOJP6WulHHbNun8bCWMT
WpBj+OmOLc5E7+fWosSwy2efAIGYl8zVnYUDtabF1k+E4zgr/eYap4KGtR3Rjy4uM5yxH6kIV03C
3NbAqf/0lN1SPAbawmif+HJbf/9F4xwIPAn+1UWJacreH1fo3dENqGUitwuZ4fyls0TpUT1F98j/
NN5ktHcGPtzhG1fOEd5I0a7eYrClhaRYM0WiuGo6TLI/X4NPivChkx5eWyLIS7ZmcqseL3jlPYio
K9LbPPc7rFuPd9eANiG8uxY6GBAjC8asiyMRF/ZCeoojvPuquTKk1AGutFGeRgbQLfj0FB6QrFHy
b/+v3hRULcksT9ZOI7gSOqnSkR20kLK6vMzFbqoky1LOpBhpXlvEKwLSZGxO+VK4Az1kTN0BLZKo
z80fqRQlOLhaGTC51rtNyy9zIouinAMoIKPd98CBfttEZDzHshRkF6NfZYbkSxRJ8TFg0KnFbW16
hKFXCTH0hyOj1xOno4UIVx5BP+PaGssf+9PmZ7NBFycNyqSRvJX0KR6i2xNYShSCcIxaIZsP9cQO
JUw5yfahHKKA9Sn1hhzpNjKlq1zQGIsRBFQllb2MVHousf+AsUxQtp5fwhJK0ilNYxiaB3yeCDaV
4QrLCHOYWh8ChMuMQDh1DwKk8TFlnDIc7zwQgnHimNMgOPPqWOe8q/D6xFDW1Vax9H3/zDu/nWJL
gGMkGEyku/uXvB3P4SNCOpBtMJ0GUwrKkkTZU8aNq+WC33sJ+iP3DoYcR0bITjnQ9GvH29KOVHss
LAgZ1YKSeqH6hiKOGCiBsLN45rT2loSA0kYO6J2W4UTw5026kRqViPNRpUJ/0uOZpXsvviIO8Bdm
nerrpdyFlAVncWIT6JaLyfsqkwnFQgP9ysrp3gfgAESs2ky21UZfQnhvfnNxINV1fC82rh1BCGDE
TH5KtQS2Xaz5qfXeSMTgbfYKTR7FtrkZw8X+fgpLMmoRe2peQhG5s5xl2QHTfN6HbugQ4p0PU5+0
wNE+BxKwKQbnMGZWPISR2E1kM/cWuWdxjNNSFEPs6iKlJwiqDn9xPpb4pbXMgFmXeK5UHUfZu+Tw
igmQC7gMVV5yPuav1zKweRJ7Y1WuBsa39E0TgDqBNsZuqWgGnfmtMu5eqcr2/Si0IhUvUEW5HYo8
c/x7bIu5zdwUw+nfLJTsUoZUocAFbS1eFdmOgEHXztoHvHpnOeQLh927ED1OGTXtZrLmdtyqfMad
Q6PB2g4Nbm/Oc92N10F/0YeMN9hkkJpwZYeKYU7gf99EQrcLw/7o0rCJQc7KWX7/CpuOUQYIY/nP
r8t4ZBMe0kWHfhO86ToZ1+A7LfDeVQGj3MjI4nHBZn9Gs+j8j6fqhrPTdHNCf2i72c/2dnIDqOvA
wRcPNH9tIfgQ8MYjIYAGTyPc6rZUD3aRkHC95Lkp6ZuOl5P23ieVidftankVqNolgFUkJc+t1glA
ed/QcV3n8AJYFjGfVCuA6dJYwq8J72olWT1BZ0jVwkkEXZ7QXtAQCGEP5pYU37ex01IfWjSIsTa3
e/YGNeeqOae2KCdOarjGSCUN3rW3fwLg48vAUAR65ZR8UlU69SbEHQUS6Pdw402db94aMuG5Dnhm
gHgkAqmWMGLAZY+KM5r65EYbD1LSlUQQenTiHH179KVuWnhjHujtqRpWq0PAhjMaJMq+kNAjPAeX
cfURoaH2Vybbt9ov38kavy0wpw2aK5sYOdtr5K03OISU96Hm+DVbOI3mLMowAc8GZ3ltsS9KCZy8
m2Iip4NDnXD07M0HMae3w4cH9W6rqJ4FmGHuGStNA2WbhXLx94exLP+BFsx8Sbsmcna9XVsykbu5
EfCIr+ch+Ky2vW+ed449eeOTmHjuR49tQRUzoA5lR8MIHbVktCdlD6/L36/Fzy2+o8BGZx3Y60Hp
csq4CjvlrjNPBMsl48OBZ1DnhslLyoUXpXFCaZ34+e6TkzRaP7Iom043dZWBhWQ4dGzsOOL0iocs
y8fQmlH2lceON6n+N3o6fyfY92nTUVNBzoLNj17CcISZmPEz6bYou85dXhL+TP6P8enDd8s1O6ri
04N3t1aM5mb+H3ghHemFXiWRkWWXKhMVaRdZdghd6yetnOj0pK5HbDESTJ9gqpaMovJB8/3LuCC/
NojdrafmFTv5iVcNAFpmgAe22FAKh7G93LZ+DByLBd2C9lYuYtKEWi2bi0tasN+cboPxJRNS3A0B
EhjWcH6X+v7GJcKgbtXpIOTLallHSGQIxCwqpg74rjFCykXkIBfT84oa4+nyAwLq7+QVsgImzGt1
ZJSkHjC3xHjR561NP/j1mp8PaNNbBFNLLighORTJpWha29v/KXHj5eHWcEBvg6cMekaoizlbDOSb
lWIoNDm/KNdzgu0VoNwsIaHfD5582W0GBNIbHStBNOKcsGqZgfY8+KYl/FpfbB6Cs89zRvmZ3ufv
pd1CTPJei3aXxrsptPwEyKyA7KX+TepB8rJJo7OKnZ5sRw5gnYtDJJKBFuqyJA6Ca4HW5ipQt9eC
NLj27RZ95OgvtElWxwV8fdE+OUbmWDU+RvKKns+aJFvRzybSpUmc03ddX/YT7tr20GJc2qs5bPkl
wGPztelpxXs5q+Fm32cxU2kM7BRWCj082TujwpNR4bfzFPULqxmeTj3Sy9PyXisGqiK4jTQBqQKW
rzpUjquUluc4k83Aa/cRwARzWdWtrf+jQuyvEbcJt7l55wE68reyF7NLEryB/k39HxdcRmv2f1Hr
9fSQG2Nhin3Fv5hvoxhbDXZUAL7SsvJiEpRA6AGfMWp0wQRSr4xrZWOr5m1vRUrFk6XdAsYUOdRZ
sIbIYk2iKTGbWQTPkT3lCPIau8bGzXNaNQ18ERUoFasNWPsLPFTPsq1duocogVbzjYzWUNfK0l4V
mq3JOOZozCuOViXZqiC6JZXLdQWx9U5wrr3StmpVbAsNIPRPzf0LoDlVY3vPe3Zyup3lBCjBAAOp
huKGKSyb0v4zMpZtvGZmloXuMp0xN/bo2B4x4Q5tcSJ0zgaZUmix4El4VHygxAeWAWEQIdpVdtOt
IdD919jhSb/NWrk0gBsiyBm2FuEiIL7LSVIhnteUO3pp31TbzdvNkCbaKVp7aqwJ+snuUH4AIj4I
PWnBLev3e1jTz9sm7S5MPr3XHGt/imr12h/vXlzd79ysYQkCeJQ7H88pVUBVlRRfDpNfLn9qJXi4
OkWRzAR0ZbOVlKtS+2WBtB92e5Tlx+KQuI2q8tor/VUpslvDjFrXQDRaom174bF2k/9RCLHd7Idp
2wiprdoyH7Vj1bmbt5g09mNnSc6RJEUrcQYWvB6Ig3yEMiUV+ic1IMpsq3wBOfbi1xtx2FqVrTuv
9wXB1rRAs/aiK/UvnmJxeYsYd82WGarE6wjCFZNHZcS4qO+7CZiL/ta8rJ6og35kVNpzxGcWLYmj
lGjiiCN02ldu/cBrQ46Yu1+9XNFjXNh3InkaddxIKCzfFASAMbhitXt0TeOdSIY3MZx/tq0DzmTe
OeI+tP9OUjlk8IsvGlIaHRu7rKp5wmWwXCCGkpyf7T0FvRe7uk5sXzIh7K8st74earSMqc4q9A83
k97pqQjcersy8ld6cSUptQTimUG3srGdmRGtBMNk1yKqT7zhcmE3WMiB6igLLFs6o3yHWcHLyykS
3R6SvnMOA8YMKrZV8xK25k4T1j9GrlWiRBYIPIX7FY9hM3J3p8yGgC/3LByyYZFf0sfu6f9Rao4h
4gm819BFNaIqdpGQbUkdabloyaYjXqTCSCBy3IStgpJGm+9OxUK+32DSHxjxMMgwbrSMwP7AXeAh
6b/36QgBbxsgWbCNbdPmMu/yxhicQ30Yk1Mp6sLO4yyC49k5XvRIgFSqQEkz8vclD7OqBwqerVuT
nBTTYK+uS/zQfbgAxyJTv0T2L5I8lx/31jx90q2Mt1lIgvGX+3ZSKlplACgqeMp65r2U3k6BotC0
5+Rivy4ABhPSsjmIzbHpsO/zgJM2435477r+4tGLwXRyoaWCcIj6DITLuzLekNcCXgf4qKrMRYtv
ronnQQ5MQUxpAyhCcxR7W3W+mNr2WMBhYMz498UmoXCcgjQlohLQ0r6rX6UMksfBJgvR2tjlVVsJ
RT7JOcBY59ZzJsDG6cnnFkZWU0jIg4ISM1XNnFxgR/wipo0PbXZPy0gXQ2nQwt/gULGbvpg0Q/i5
WkNitOgpqYgF4QnhTXx8Lgc5oWJtQdgSvxeKcOd5Pz1VG1J8G4MG6GBQex5DbtpuLwlxEh9Ij5XU
XyXwydzOPm8icwGG214rN6UXPXSPNVxt9VOWghTmCXxr7aPy5HKzIowZMNNvybFRsReeQRtFtHgm
Q7J+qA967gZ9r/0UhJzyr3K4vZU2NFsaoXtyEktGuwTyGXR/VEvTSZWt9tsv3jfns4NrAD0DlPap
YRJ4+0bWsx5Jik/HKoHitkFc42+82fRA9E7psxCgvM4+x5VVEvRD2sStUplwjZ/oYM/g7t8a9O/N
CLkEY6h71ocCFp3yw0pHF46WKXpqloTnQQmbUDnwWADeyhOuCWA61OszFweZSlBbjkzTRJYIZiMu
ZX3fzoak6yaV+NMVkGrq846MbK4IsHDhJ1s9nPWJ/OLBO/44G4BF1IFgqn11u3/vfiFuTh7B+kWo
WMH1yGNiEe5O0e2Toeyekt4+dAmGNOZnH2sF+quj3BtFMpY3isvzcvYjQW5d3W8oeKF1DVgTIh4y
auQEgldrMQOtHLq9ATgOg5N6czXallln7KbCF/m2tLUSgtC20mK1rEAb78a4Mpmi+eQN2jPi7PkY
1CfNh7EgUxxyKB1BoRlq8OcP++qX4UuOI2/QyGo8UsCuGjIwwTp6wK//a3T495Mi/fweCUloGLAx
AA1iFXQmmgYk3cpeur/+gnGA+cWyYBk/4vhwOgQnQLp6iu76IDeHaIJ/HtknyWu0ZP6gcYrgnFcC
dQq0675Wb+xJ1us4lblbkf/wjjKa5RXfLoJdNS3O7vFjAlhmJewcw/0hFW5/rQm/9ywUnsqZtE8a
gx4a0xAD7P/map8TR6fxMLO15HS+i/+lVNM8x0BEtynCjFWTsl+k/OGZazBw9vD2SB9pNPlVET3r
K5mAyPAXdkaCA7vgbObFIX6+CuJP5tS1N+iMS974CX3w7Sf/N9OryKEuk8g/d569plroCb8gcwU8
WYuXggkrsnyNu09N2gS6sYYMXV02UPYK3hWBjOj4bEARtS+1n27XQ1HqnxkdsTNrx4um7J5/+4FE
t2LT2w5SlChd6Fl846Itushyvx1eU3rIsYMNDwtVDJmSqUrD1AZsHbMbU+X4ux8l6POahUpoht19
K0UjLncZkDEz63maJ4z/4SYMEhWfLoixIqVdV30+wdx1AHzj4PUvhepGduQeNDYJu9zNfy2/s+NI
YMKNwYxpiLCkznrBu2UyhI/dXQCyW+5fjkbZsgMHE4xWJ5juixb5f3ytFYwfJT3Y/j0aVtEooYpE
JSU/+l5pOAr1Kd0eF3O7QRdILO+Y0tmXxXuWnNUOsaxek7DycZHP8O/77joGaLsBjVUxwtf4mOw+
j0fzrCciQEQPT+JZy+chfVE2DplEY1gFHKF7OEHg+iItkz31JAmiq904yqRagJLUfPJPqAAqt3N8
YsvI3Ybvr+GvsrP9cxCPe4GPGxSlNoj77LgGGmymXh3hOosSGb0v2WgGuiJYELpugAkkUjUBEr1C
CCU1v3vJqjPMOi24gDK86npaKAUNNvkVCHnh4g8S/SYQQBgEl4WbugsuQXiK/8ypHBazwY3uKUVu
8zQ9A0crbZCoYY2KCUdRlGnbw6cF567N+Z26qPCrB6mSbomnlwUnj+o5txgFrssekbnIhqP2KUpJ
j5Rwp6jkICU0KmlwqrUkGCnaL0cCIxNQq9q5Ht04gXwtYdEoLskfFAr8YC1f86XnzBeoKDzqxycw
ov2xGc8buXNVnpPIuq9dcnraGwGuxslZeGuBpNuwJccj1wCYz/4Ia+yTfHCAcmkiLgdRd10SJ4a+
/e+BJVeEgobYDa8VvS1KiXkyHX/A5dQwPfmUUTmKUDFn8sKYl4j2Irt4iKiViuRIHn3c1A6a9jsS
Dow5zDpAeSh9qC7w/eKf4m1FvU68CBnJRHiMpib2twZcbVDd/MYAipfRS1dXvufNbk9dG2Of54/L
yETd4HISsiwEZ2nDhPqQ/6xl4oJ2q5nEttYS3SusiAFSs/x7bTrLVHYFvOuV4aqBcnPqCUr53Y8K
ASbrR++/6TZ0UNeX+EaBKFfLEkDKgt+tfzhSAQZt9Lxbp2AEu30TkOXDR5MdGJ/DuSq3wRYonzLb
YAZ6nUowkCJ5wD7fjhZLHF6gqy7s4IGbp43aNXXgqOdEKZXFQBKGgRjbI2HpXDPfkcQRvFZdLlu5
2FJiWKXbi7c9RI5IHuEG31A6DoUqYVct1Qs3UNgYjlZtsLUUhNph1MSjx/Kg4hL631SitcU4YG6E
t0tgbOil2mUJZEZkmjk2wH5DGM/rREPJxoaB3XxNjsfeBEjXjyHFCazq2nYaY3cacrvm7d2vWNrX
Iu0Ql0yBG6gw0dy8BADzvoqKaHgEVM1b3WKwUjeHg7WJjIm7YETBtx4IzXKBz787b75k40QMLonH
I2njzHdv5CA75kUJz/xwzTDME6J4w/xE54qPVrP+NSWdZuvdpRaGnNRZ0nkMQJucTeC62WnmvK1k
lhsiomV6YeIUHEnT+dEsSrwFpsOaZSMep5leXnt94T6iUvyBfo3chVZUwvbz+n1C2m7fMIHIeK/K
4a2QR24dfxwjRcixPG8gxW1JF2dg6RiN3IXAn53YKEZbdcyYZ920ctGZz041zxsdVjpQX9PP9rGf
0D9EIFfQ1iQZJ7Yp/EO7vgloCUv/6ZKPqdu0iLaxvmw/OywgQGIZM9Nsmbyn7bwT9s8fb5DUNzha
8bNkchBIJoEnbrwTZe98Ovn77DU2RUvpR3OV6B848N/6zkbxWkw36OGoDXNskKwt+KqXObe+PN2+
sfHdHdexUECqAnGaqRQXQ4y3s5lTLKJFI/wXxDXoE5T3YrpVFS741klSoxPZ0v/8U1vMzz8kEw4H
impKnbESUSxZGKWJYUQPxThge2TiEsV6P7NBFJzmzOZz9oT+e1Ohe0j3FQUiaUpP46y0jPG/dQ3e
OWM05Rc3opindZt3w/ntSFT/IOAmrKqE4yLOqgiGG9ZugPBasDY/NaVHQMpzvdP4ixMc+J4qFoEG
QxIX4qydT/Tn7vwyY9E2sny6eJmR3+3xty5dmoLuyVomB7WJTwlDAKH4HBo7K2wXnh6az+dQw82K
oJAWVmRt10Cbcsy22BAerz407SRb8alIC9ZhCISZkzpe/f9TgbtEUjJpi9l0Tv5xkf4Qs5Gl69/v
sR1ie5cAtzoItI1UvacGKzxiL1lUqfCrqDPmim7Fx5EaeA1e29VIo4d0EI6V586RMvVmdPfJ3gCU
m3JDoWsMe45AN6zos1ps0FvbokPIx46AjvqHUk1U1fzlw3z60oMuLv1J8V2hihEKW8ZMTCfO94yw
yuoM7aw301tvwyfZY7eV9CYMcC6wzgCjOZ/O2GZzG0zR+g/g6vRFlEGKgTLjcFqK4TmTUN3ogay1
lT0X1uNeFVChaxNO5iDH2y//zm9M645R7uyQwwrfGkct/qVf6V0NaG3zyFx8/Us52CzxxxMyTWI3
ztGZL44cFdgoRSXAU7xRrY6GTLz91aLCWPJ0uO477jhyoZUbzarVv8TT8nfvYUIzUs3lW9aBYKY2
/p4DKw6ozpCGZdyanwDioG0odssbo5fkmSZ1n8IoSnRUQUFi6I94WYNdYIV2XTD4FdbDPrvUeCzP
62DyRTEZjuy4BXIV7l4HTrv8dn7pos3+TZ5ktf+k1029M/vJxN9r/ymPHDzoV1a4B5Yo+qTAZfoB
5YDyP21d6onDb2W8x6Bni/oRIv712tQGg6/xAdc0iMBUTXobyGJq/Iulu/uBSMar8+fNWawtzZpg
qw8eCHzIR9vFSUJS/gWBVtlxGv7BFO8wtHu9351vrveqBYUP4c9ZdX9f79xO5XeAtU5wgl37R19F
OYVDkur9iH9sBFktrzgRqWSNqmNwXB53EoqU9cuHf/ezOtgI/diQaDjlJ1jlAfRpJGy54qYjpCIt
duj8zf3bYhz71mcfOCyuWPbcDd8H+QoWcaamcexy0mzZ5x/mX/dVmeC0hbY2RsaHnKoIEka20euH
jKL79JNH+B3Lou6YiqSkq7hsXXwo5jtG/rMw9poO+BoABQ5L3BOaqQYqfQ9ullRoZSLz9cWVfvu9
QRdQMuDAWbjSRag7I6D9MZwDI6eR9wTUNtAUsk27YgUiC69HOuBGT6s3NkA3jKiCekZgCHa22Yg0
rYcYQ6KXc3JzlS/ckV2cX5SZV2+IqN+W88A3btl7D9kEcqPCTVAuRB4riVX9sw0FOd2L6FGUnuFa
8p+4cFXxwnzeAxRfvI41XNyMOfalgI/ShPL5ZYZ7ZljZBImrUA3B5rjfPDZE1wQCFI161uiR1zKA
B7PZzJzRwI83K618vcpPMUCpOvN3SweIVPk6JrItkRsxH2bzNiROv+Aqtf2knfTGPJwSxIHOkFCJ
svWAkc7QpcrS8fFNHyYY3s0/8O6glwHHy6gXOfkn2uEVVxFqDUAN/upckHmPaaEQGqZPpKWn+kO7
oWqapPoaZq76XU+OrH9R1efIO95AFKNn+X7QQPD9wfpJsjJS9dXoG8RxdGh4KQYsSxqT3doY5kSH
HTfQqj4vM3dBP0Y12gomNiZ3QQhAxwV0Aut7sZCjZSpLkXo5rscbm57IG0uiW502Oj5I+fzJUnuc
Cs3ccKYEK8Jhbj96+BriMG3xrscNuQn4IF+Z/Gsxkp6ITtvh3UWvFtvjbZx/zH9KukeWF3QZKVpB
Tjhk+gSgLdwdGTGDQn5yakTxZtJnGp+KIPFMvQrRhXqB2VBPLpwjpqcnaexp4MQjvdRmk/5XvJdC
EnRUoUATVNew3HFbI5EisA0wtovedjqUM5FZ0NgG3wOI2ZNp/Eoir4LHXthVdmbxB2hI7A1NETgL
YD4uyVOBf5nYlOG16/OrAHXlz9Mup2Q3Pv0owmwSvsZKiF22n0b4CI1wMggNGqKK+U9ZFR4rOBLU
W5bH6OuWRwdcf2/c+NoSIsBxqQOnghX5l9QP9OmnELWCO8l/uMQKRVkorwx9XsQyRcWTATZ82V6o
mXliUNwrJI/aLdu1lwqgBQajzKV5ANbpgpPpanSOkVgthy2fK3dmmPcQEWjF/D+i2MZcd6ILSQV/
VfOx9vHlpwmXsOrd9m1gimi7Fo0/RtZbEfCP0P/2lzkr91/QXPc+UACtITESAu7aXpam3eijhBWg
VD+An2zFl8DC8EkfgGJUdQAVkJkAT4w6miBFvRNCzp9SP91mW+s2Wl2+1qCgmWLLhPhSLgjO1H6A
4xpUNCCc1f/IfPp6qLhu0H89qLlenXFN5fErecwDbhGiljiIDTp3hidYv+D/Eh3HHBcVOSi64xdQ
P2CRkB9Hd2YZIQfcJqssyiIy+stbrcC5FspggVr6r9ItC5ZWmFRoyatqCItGYc2KpwmXwzMtf1nW
xHYC7XWjGu+O+cyG16NpgExum0nqQWcQTCzJATGBKP/BPzDtqvpk9X540o6VY92fXO1JVxP4zoI5
HkrRgkqQRGEnGnbMkuffqwA2IoUGO+cBr19Qbe82ASMWK3bs7Rw+ddUPktpZ/eubrJIcNFGZTTrE
mKNB+vsMagr7NY6WPDVN/gcXx6iLU53ecZOM81Dp09j6WPOJkOQYIiBnhhBdwzZBtV6xXcwdMncx
cq87Jfpq68/ZdBVj/WitaG97fv2XMMGHNnIONBKdu+ZXUs9t9tPsbooHrEH7n/nqVPMhdHoq/Y4B
ZB2Vg3BY5ydXkzlRA5Ujf8CYLyAAkWNu7chBWLZfMr+1dfHsYMBqFnlYiyUKm1B8Bkyg3TZUqIbh
5MkGrqQXR633UdR27Aw3gjvDLAFPPyKMIjt1aVapW4spFhKuqOwPWtu3QHCrYNKqyTIqhdQFd9eX
ngBpZI3HFJb6kO4/uuoQq2k+lmoSvtv+23emN2QojL+bNc+NHwyhMZTBPDqoEydGbS2DfgPH0cDA
nhslLjDkq1m3X/z+0AMCzQmNYzd2mMpKUmy53m0+XMI/kajUqVWfXXRjHe92qH4htYvIxWOy38sG
sD8sM9OQGfo2searvf5MLsOfekp6Zd5SxVV8Df1XMJ0sKYZ1Qizj9MW678oqucystHwrZXqXOMC9
HTuEPQEIh2UlnL9pXQcF3zM+1uGHe/Ub6UzqQwuzYRGA04XjxwpIPQfma6Wc8Nz/cceCh8M9XK04
Kn4ehH4OwJT+IHs7NsqB18KhPrgnNDNo9FLsff+gya/QTyaOXB8tyCTc3nomz3iHkz9LxlXVNUI3
aqs1KHDP/3VdBZzUQVuyePMq47YPiUAKgmmQc18CSNwcO+RnH6uS72C/3J4wOFlfTVWZiWcvNRbL
r3pBVDZyxQb+vV0LA7+kkKnRAMBoAJzyTzW2Z9NGHNvQTJtJK8Iz21/BqYj8aZNTU0VrCCzOcdeA
dYmQi2hGbL36TT7eLdA4Pe20I/nbs/Ayr63VEUHWbocA5+SCPI06oUxtNDwULqR+H0IE+6P5b+Xp
PuMKmDzGgQxsxLSt5mjjdXVc2QL+Y+5s05ZL+OlfoWY0dvMuzORlbier4MX0ajq5HEaEoq33jTAP
S7bSuzGRJWMCQIp3zsQkZ1sryefNwzky0tQoN6od8fqnNhNxxqOrKR+/+6SvZl7HtrkDUoH9KHib
Cgv54KblOCk0WxWT7T5FbS/Ch1KTDeG7KOl1cOcGyeccPAJKelOdZEtwT+89At8jlMmWX2ajgnQq
B6UJdhEtfdypk4y3ISzwTwc4m1xvTEs1PXvKUTV7X5oRPKD2pTTdyeKuVP5RabKeMp267yKJd9gC
EFs+QwZd/tusXMHgJHUWDX4rtdzwOBps0xK47Whg0I/7vN/O5TEaIa5BMh3neoivZiaLOzdrg+Xs
Zv9P7aJCySd/iXEdLYiqDn2w2MGWKu0IdqH84E76+sriYpQpYhLRNiFWYnU8/dMrkqw6B5f9B2Gj
nPtCNTP+U/Nzl4gH7JvAxyGlj90mCYviiejAXb/nzoPpomOlkWWhSd6cuK32KTz+t4AF4+2N/qNy
/DRXZk17/r1ElXQpAyt/VSOMhBAbtOod4uQ8Mu5gS6DHlG4LbiabFIpfBdHhurV/GBtgdG34qMVz
rBuea7OBizW2KUjg9GyfRLBaGSp4NRNAtV/x1nLmQ1E2XniTnoaDprWtxRKQ153u+NETZ/hVCt3q
c9cALcWl/lzHwaclLYWG/m6DQBklK5G+jjQRTjiXzE1JJamAvql7seYYRCHZ10ZgYCnPMtPUJmEz
nVGS+frBfQHSjHf4jqZsE5Bx8Wy17d3eJ08V1aQiCyKHhquKzjHP+oKSCm1NJCycm7I2obZzZOWc
/gKDsxw5UMzsbjk69o5rCNtSLiZYyttfVpCfO/IxdiphEkQjEp65zCkxsg9O7/9hm/FNB2g5AHuY
cXnPxwRcF+BGCznu8rJ71T7IxoRMEZlnoITFP41S05jBjckA8xJq3+bgneILeNRNDVnrFnmB5+v5
0sBp89Obm8ijGRlFut9YMA79rhuOhF3+VjjTE5RWnqNmmX5GZv1qFJHoqDr4K4t348tKLDv3ciFD
Ly2JYQL5YWtbkPtfJzgRXpcOeyKU3BQoK20yNp2R3At5AZZpFkS8FDci0B8RTi09z1xOXTsNQ0SK
846qVLZ1ipWq38w4LfJzpUoDjNl/p/RtsAn682eGQVyLPtF313rpU/HILtLR0MkKzeR+j5o+pknb
fyk/6UQH1KAlXxghOMTNUpuHsC4R1/9xRlWTywd47EjF4KhSClx+pJlWctRXQPV0Gb0BxIwDhEg5
v9cnPscZjx7BEky60s0sBGYhMWtgDRBfJrFRnyOb7toH4OoQu/L7fI01Smicu7Y2ZLKYIcBdQ4m5
5bt7QTQ8AY5YFW7L2A2wp9Pzl75SwcS/0G4Spb5EnGzghV533ArtaeYcNSX/vXGZe+S4DDc8BL4j
YueKD7HhrhqXiP853rbgJoxxmXdlWCqb7CMqh/nv4UUF38GCc6Yaog3wyd95WtWZFBXRTUaLe2h6
ohcxpm/eU81ipyKCjjf6tetlGqAS7HS8+EEOIzXon7TIEr+INLqHyLfch3v/89THfcpofMu/1VG4
C15i9BxrlguM7RNMdMG1ke1cZM3Tuhnmao6bzyXLqIcKxCkO4e0FrNrZupAiY3nkuIr1efyCKXNH
c+Zt91oP+VUh2DoPthz4TC2ZsJGGt4q5oxTn60uMxjhpb/TtJq/bJUE1F4xEcJvDXD4SS7SpD/Mp
c7KlnHbUxQJBQ0njy5sbMQzKjhVBCttuBjJH5/1yuEzuSVTDPKcdDJAgwCe638QRWxNTgWTsHSvv
CPJnxmaitsSC8bA5b7J/1ygx6raKIIiUV7kqe/zQOM8xhbL0pJho8cBhW97YoGRl7BesbCIaIFTC
cUbLCHqVvC3FQbUyjg+5THcw8GFJ123ZQjlpvkyJkE211qMsc1EvRVkeb1PQwX86yNsyzyEjeXN4
yDF4LbZ15AfaK2pr00RAY8FhuGnGKLeJRmmVfZBbRvQJQxNBJQTO58UNMMme6179N1QsJ9g3xZra
PGvtN73Y6WGqHrcZ1Txbn9Pu8K4HIKt+DuQaFcPTgkLD0PIIFbXGGNlVoq0szkYTui18TgF5i9TV
SZwS+aclIJI22Eb1lvefEGkeyEjSyUEf8qR02dc/vTQTYpvhpz4nYCEe/pi5P1Z7zT5TiqjcN+vD
Ovb84/58DGigcP6Wve91xkFqs9615/e10QHf7COAWdic3D6gNOScA1fuoMuWy+pXPS3qp1FUVB5Q
M4kTxB6IA5r3vde3kgJgruIkLphV2MngZsUNs2XGegElNe5JuTSzzG9xSAz06T+k4LhhKrabvgA6
ukPPoysCwMfD5n9N9Jx0ta9jfUHB5bQgQcIH8QiQIdFkDGGapz2nK66Gu2kyVp5HpLvEsnL5TZ/x
CAUbXnFK9fabqNr08lE+SyX7t+IQtK8RdDNNsxY/vVueqIWaBvEMCO3/w1MeAiie2dcWhWeYZook
CdsK5tme1wKzYK1rufF3QVQmlhrvsDSJTMqJ+auUKw7QEou4BbqlOjkoOYpXyFWYQ4Mc30IxAzUd
q2/1RCKtMhexE2iiu48olD8fy932mNzdqKp8OU68SPjQjfoQRdtdFJ/B7wnFNkFF5T61yRRF3KyY
CXbdtw8O4h7kx1+wEndf2Bff/HHohZNh/AGYD6abTK+LiECrr68XerO1aSzHroSbq/EF3q/ALITr
mctnHtqvOUkynXxqzTccj6hXnNk/UliZo3w/tEctiMWRKD7S4P3aha5bTAsfnoh4+urUK3tc8J60
X6BXMFjOZG4LWuPEXtksUkhV/aGI8VABtlAHAGMZENqQMODVRHUl4x0Y4LOsX+L/c5h64YQMulGI
LY1P0kspIddIF83cQ61K0CPnxrs4IpK+ytBxI6C1K2GzjvNOOqUJE/5OkdATvTeDM0WYWj7IvO9v
KbecI+/j8ikIZv9/NKArzM44xyE2GSwd4m/KEkdMspThAjSxRTGA1I8e+mmfP4ysq7INCZWlYknV
1KL+yMm8sJLmysaYZPSDfDEYw20k3lIkPd03dI8pa2AmziZDs9lD8t2gyrAkS0yBrcj+433MhoXk
h6Y+7MBzm/gd0Je4vbI4Y5h6WGokM/bBc9dR6H2Vzkf+xmNbgUxFBOSVFYbH3WbiK3yPZQi3FuLc
iNQSZYamON1PF22MXox/OOd3BVBddPmlcywMc+3lz5P/jB3dO56KR6nQjsv/rJX6yHKX23tLFRN4
ieXFa5+dwLkgbwpi64Wgz4c6dDBVPZzTwC+N8Pxq64PgntiEz+n6Bu8JY+pMMrAz6/45RX94NmOY
T8vGbodhMXTsWruFXQMd1vH3TEBqA1wriDhONErWLsDt83ZEKpLcMVGNUZ96VQnZijEII2Qa01CZ
1QR32hiUZJD4wTY7PQoVSuHzyK9aZNdycryPcsk//Du3u2mAOQO65n2lbRVXiIdYKdFSYmHP9GNh
pGca5rPooK1Kaavc8LFX0Zb1EoTL8ve6MnIWTWxmlPyl/+woYfDIslZfrFZ+afMh2bJ9cdqfGEtk
enRe4wpFbxWnLEIUNc5WrZr+W82LMza/V2ZPNRTRmfffPB9n5qfVhqc=
`protect end_protected
