`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TMlgMKa6CuSsbNQSPY4ecLOxPZgc92einnEy8etO//uXlPIvQ1qiZ4g23RpPqg/jXfZRDjshOL3I
iDxV6dAc4Q==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QoKGldyGaOpttUQin3e9eu9RMzKXeHPbSaHZNwQTGLOTXKwkjNITVZJRdlmxHDn6OirKu+rRFQ3F
wCZ/4vMuZ21Gn9+sIrxJBbCwlkCPvMFFfEziD5VC7duz/o0t/v0pjBiE2UzrCzhX/zNav5cYf4tH
pwzDXypqiGs0S36N1Gw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HJLvAmdAUNLnaTOjYW+iUfvPnE+/PxLm7N+W7utJxjX5Mlrebuqkl4ewozWCwYMAxkpmKLhSAl3a
ms4RYNng44+YY7iX4QhTyPNA5H6q14SSve9TLLjNnVMOpHDy6EhmjXFD0ryIP6utmSfn9p6AA+yf
zhDKL2zsH+kDKsKIu72NWKFp4KnVk+Xri3bxYIV6Pd3Gf6paNdVvXFwcGhVrHLW+gnPz6q/VgJyV
oWed/PzQcYHE3xf0r0wBnho9/uc+KQy5gdGXngVVq8Vh/d6SyTSjP5are5OOHRPMgpEBMYtF8tZM
FCa4ZC7a65iHL6+pFFUL2fRYA3IIpe/Py+e2cw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q7v23KsLKhkl86iLzwsfkiPrw71r4zeRyKES8JFS3Gt07O8z+AIWU2HBH6QgwwvnBx9nvA8MRTSX
5edZIiNMjf/mFinVNOH/G2bp/LQgJvt053/IOUVz7cjLPG+l3s/l9q1Rnx6brs70YHo9hg45gqss
x+p6rM/APyG68KcaqvB8z/+7cIaqZb+cutuppIFEghNC7tteQoKY4D0VW++ec366dBz5VO1UPZ0f
rrBUhhFkja21HOGD26llSDryBKZ7+ZR4Wnzt49OUh5XtJvEOFcVkzYnwm0nRKqxIdR0/1Hd0rTKl
lAJR00fTrSlBX5qN+NVUlOA8YhuqsPlse+cCMg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bzyTMVwbJDyYq52SCMZVo8C175LNITaI91UZF9rxFP/mj7Gd062gcpXncoT9Pu1J7xSfbZCJiADG
SAM7iIHZCSX0pYnVB2yJGl2C0MATQ34CFIF65YaJ/DF6vFPgSv+Y8d6wBhtjovhSm37gF9OlxAEt
K48UJFqFj6iqVNssGgH4iXrQXXyR4LoLXFupFAtcywZuqTMnZ8xGny/tMIsilWuHtXBOsyHFOuSs
Qv+y1c2psPEb+7c5ttZVm3k2HHzajvTB4dqEY3RsYkKSVlqdyHCtwVsWS17rV+yPUMr6+OlV+Bma
ePpf1bY2rBHmrtFKfEVDhUHHzHSb3WDMjFlbuA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jrjUdLS7qwzjwVXA+zskeYgeNFZ+g83Z6osl9Iyc5gmi9BGkG2U2gWJe47dfsOO9oxW6X+L5LzMC
sq1MUPLrz7A+9r4Uy+nhmgZ5liwXvOm/W9RHAiYNNUQaMLMgEqYsUB+mk9WrJLlOd+ltnxV9mNi0
a890FqGtglNhIhyTxMw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZqWgCo80iBhH84p0T28/3oKgMSztFg1E8X7O/Xq46RRhDxSJ/dys4csu2sdX3z2XYylb7w1jzwBU
SELZSD2m44MHI2jPm0dFUSjAvaUwaMBps7rrlCemPZQ/4seZkfcuA6fo4itXK1nT/y13qEQg4fZ1
5sKyfJdyQ1asfyVqPtkAhTSBZ3j7yyp76p4+Iqf76/7cCK3yzujObquHQ1AK9DRmMbEXPegD+NX5
o5XXxW3KAfKxXpsbTvGJVRbho2zLbVRpxLKUVCZJ5XxLgtxfVip415FJEAoS74URcfZnqbzLjzLH
UsEwIXB4KMj+ejdCr9xsvmN3Ikdz/j+Be16E2g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
jz+bVp/K7kEQv7t+d4oVaHWRFc8t735tZmgeU7dp87sH+frR5X3zGlfYIA6NnOaOl/7oidbLnwoe
giscO6xuNgNnjuVrWHaWVUZ1JbkTsFA2cEcMlYtwFEH1grMuNPgj5PG4TlBFQ01/izQvu9IAXbJ9
eBMJ2QY2pxzDqvQI6qbxWDyitqoadyyidM+zc2rcNUBDsfvldybNMEcBetIC7BiT8v8+0J7MUMrX
4bvOFIMG9XTc5gqRPlw36rZ5L50xbUNybebmZXngr+Sm0C2TuKLutPSAS2ulJGKScMtp9gxpFxma
xNkYdEnXwGsiRXhOetOrxlYzpP5IP1SpDtXtJXSy/UPbcAB+S+5kViXsapebNBTSjkLTZN41uheC
OEsIyS0GDJC/TurhEF9HFZZPVkijfsLnBq0q53URChWrwCR1Ggf20ntcQaYLqHkC+H/sYmg/y9oV
0rU+iQCTTnAzyhcmB5VTzFI3b6dOlLg1n5U8lv0ukv755qfw3CxNJXzxeql0lG+qZsMKZDfIDaci
okHJ2VwgYoyO1mFO3FAiim3TKgcyG5QfKRk/BPkEJhJAEdOf10FqmdblF7lQao2UnlgDT+2I1pNC
ShVniRDcVWzFkva0ZpGyWAYUQAHV94TMpM+pbQ9mpZy5uPM8wqwlDL/U02seZxfzy3GV0fA5hzV6
BDciho1syur6d3XCc+SHCeKgEQpT5H7L6igDKaJCVEec0qOo3wsXAMOCgDIbCvasYVB0Vz6VaXd2
QyznIpjTQgonanruqGJRJNEXl3nZU+dhdGclD4Jlb/eV1LdKJMc8JXawHcKwEjI8xO/jHw1M0z2W
VQSYiRKTIqQPSgDVqGMcbfKp+WjT2spS5Fj2gqy0XFE9oSzNpmmz4y4AO9cYdzWKlAS2NGVToASK
KdnKeH1irp9aTgdpYp/bryl1uXAbYinCCtcRVWpW6W5T7RxUZqTeng7ZIOt5BF72fh7Dwem1pRwP
tueMpFIqcfJJRDPYsuArTStzqDWfrpyOQ4bZYhTdAfOhjfBy4CilP26uASOtEj5DTnleyr2H4o3T
4TUXpVQ6bJG8dVFmYSXBdQEU3dHfRprCwmLdENSzp6GCycj510HuHcRmppNTDI05d+ejHsa1MZ+3
6NHUEZs9nlBO5ZEFrJkfWxD1AmBy1TEZhmrou/amMeIgbDSm6p4YobK6RSmw8+vjXTxWq8OAUHQ5
wNjBw7YNAvpqZazePzGLXcv2KVlvZMoyPXXJ8D9c0Ec9iTFsW7KBIAm6JNBQ9Jkb4523nT5sHVoR
VqWPs9Mi7uJPyokYmF6x5tG/cY1bxOu8VJyMjZl58RTE66LX+38h0UNghUBjSb2BCnlvSQRLlrHo
IeB6kzBF06GTcioeKjAE1pgpS0FXIPMuHZZ6qI2JbeorunHJUMwSNC+oGJ63XRr5QvabyrS9IKTW
qRrcjYhVgC70vGx1hpOFriTpseCtFDkMV6U9YE05e+25jSGQZexuGxPc8ep2aq20gB1jGBHrDdBA
L9DXqjRUbJBTgAUriWPi2NXYLVBUQfG3Ia2WL9vAct52Nd0H113AiDw8sSucN/vuy81nc8p7lJDV
hLhN68CU6T8CFtpnaB5zX3COjvZUmI9vwEZThRQikeMeU4wlGowYUQzq+ukMEnR9lu6LrY0/UPEe
cbDw45uBddNvsUmFF2FmLKt4uSNmAxvGMVuSjpqdusftEhuinXzcUKodYtSsWAgOJin34ci1qMAB
5k2rWvRlMDr9LJyD4nVpm/8eys3bn2p1um+as+bL+6CCek6p3ZeJT2Duy3kXXdfJ66r+hOjl8QMS
5LZur5ezBq9Fw2uHUaZGlo9bOvby6Cje4zTY8+lV343i1xaktZrkpiPI07l3tG/ZxHSF7BHkmGqd
7jiFbqcPgsYFz/NDj1C8JKi0CkS3SA/beGleOexHNSvP4Kn1tuu/f+1Ip3PovLUZYlRqRuNmmJCu
VG2JfhyH0IQWYJpiKP5ZIYquhioXj7XFx+MULe3qWjD94JoSSzZNFHielFzKTk0vBbKNpjFbm+cI
CJXlyqwjPsvrqh5hDCAvu+XivOtnI1+pxjxZ8/2Z1ZTZkm+Jb9YRHGLuuM/5XWOzv++Envwixdk6
Z57i0tTS9f29TBDYelNl9ieLgTR5kIp40BAu/Ogk5LHASYkhZaKr7OtZAcpizv0XVYfKAW+NcnoH
RIBebdTPX/8lF/2ZOaA4AQjjJHDU1/hNpLOpZ5Yw9qlZqrjz0vo/EQkgnfuGRSZCE8DDn/hBdlrf
sGE+Gr++rp1zBGV1WlodItPeSo5f1vsCrFNLHX5sLpA0KQiK7ujNMN+MOpkLAgaGegB2mC5cl8MH
wbfoGx1nvZ2Ohl5l959QJJ0eYBv9gx+Fjh84UbXRRvrwwKRBCLyPyx/Vuu8f9OHHAxT9zUcSu7+7
BheVu+Hel7r+g+Q3PV9xbbNA1wtMdPy9Daz32db7AInr7GhuksNBk2nHQq3OWVtrUkuHCg+X+UGd
r97+9/sdTRmyOZKru5Eq/JG5gzIjEr7TKEnndpoHzbuH+TC5AlywP64ypW0E4rgtNb7W/9aOBtHi
a4A56Hv/lXs/tV3c+ZMLjvAxgO+9QzzE04yBeybUIsXlIZ+JemiXz4Nes4uSCXeozaWlk/e18N1c
XXVQBXo7qODGC4qGo2te97MpCg2yI8dKiOBsXzOYoc038+tWNJzYqWQUisdljD57WfrRfC4ETcTj
D7frlQaT5lNFuQg2q2dR50H4fIYrm1ET9XEufyBI2/A4eKRViUdvob98EwgpGF0aRgOBidDfoXHd
h9EyAmd/VwxUkdko0PFAE9SYD+X/eWw9bZ3CdFm7muJO+L38Ai0j3k5j8ueh2B3A+I3SEM4Kpm5A
fyaS59X7TJuxgtBUqm4I4xZrBH4QakQXgD3LCqFBBWnHrQAr9Y2JTCFotSbqEipL4T+edux+UnEZ
/bw6NjrvrXii9mPoXNH07IaAAco8U+9GbexGztUovA6Zbn8XRZVxLfOQEIei/v7ORIT1Le+KH2He
iFIaah5SbhKZF+/pKnAVMc255ibuAyg+Ro/573q/XalNPmAKhPmGHR6oJMPavhC0XEJ1P8oTZdrW
kA7n+yBSJHTGX9cyYXzqfVvjB0iodG1BG/ExC/O9jUrT4Cg3X2bZfZi6kPnYIJSTBdnA1nJUwHHT
Z7ScAAIN61NrH2wqKjfu3T1fARYWkOMwHkuLqIqiUEzg0Di7rNiPTaV0JA1cZB/1Uidwjs7WTWjd
YwEDENIaEVHfXz2Yo/vSixqv0sXcJRohJ8MjoJF7ssVG7uG+Wgfr70G6xh9nWC53+hufGLz5cHur
5WmSBA0VqK2o2KXZzgeh4jZJPqzHZH2wWMqzOwmezz/XcfuhAYUoo3YF8RFe77PciS0Uv31Hv05O
QGxPN5pb0KgbW/Zn4ankKQgnhPjFl9kxpZFfXoF/NQcYOSASykw78evhhudZOpoQlDi+PyWTt15L
i8WYO7h7bEzbWw1HmRdiT7NF2VoFwkCZMMWU3eJ61KA0AJDwEPtwD2gSaCp2IF94Xt0YJe/2GXl0
OFH/F7DoX9igrlYZpyCsue0QYgF4CAAwxpXo/q0uHi6MFof7yXKQVHBINrjslVTa2MkotX+eFMs/
/wkStn9ge+TQHFQ/5E71Gs0lBqceg7YqBCZffhE5w6pc0drEmo5Iy7o+X/DWAgulA6AMYytWXmWW
jBzCSoHAlvLBCbXe2q6PTHLHVCQxBka2l5GzdICRmWLAbBtcRWsk50rHUwkIhzynOannwyI1Ypoo
sSkOVq37msb4dvGXmG/O88mqSh67O8VYdtAMQIcotFp6hkN4VLfusllmJ9+Z3NOHo5LE4iGJMlTY
VK4pzGmV8du+1SQQtDbTwVSl4XndiCglf26w8xZRfGjqWNaS8vLuPpGFIes3gHc/bFFt+7KMA9BS
OoFqnnn5G7QIXq5MP7BjIfeZ6HYKs0YVfcBV0EQJrPZzdLYD8FxUPO6dZWs3YH2kJho05c3PUf2A
QD9ADHms6fnVEzlbaOsDL4EWiewdNK05TGXgTFxTjqke5XxyqCxGhhmL7l/jpk17chZ2Ba2DyeGy
Y+b8EiCdYYza7E92Cv5+qFEPSR0CuA3BssglO7u8Sih2E/3QPn/SaQryWW0iWUsEHr3OdT6g0VXE
rzm20OG8gxigkkXDS7HS7+OSt6XmRSeK6eA1gbRDkMs/42DBjNZDsOXzDdKz+OswWwD418grNFfO
RpReaYCgK9+RruNS4F/JiPs0bjOJ8HzIz15Uq6XuKlmNjRitBJx6TLBfDtTvVKMyUsqPhxYHfTZK
pbN4+yGxCjEpoLlPEdx78fOZTi0mPK0QHhx/Al4VosBLZwp6M/eeqWy9iZzSXsa6Zm8Ib8UCNGJh
Ny1HEoVY8PItJ6xexAZXPbx2k2LrYuj24LfIjdWAX/dwMnbamO4e8+R8wtqtS32mRP/R1Ne+oJyD
WWYBcQuSHAA5M5yqKe3mPxob+huZaJ02j7Mx4BUlE+rPmzNhoEpEEs3sZEb0KHoezXn2GlInNqv7
MxCfg6yVXodeU+jj3Qjel23oGHwqcuIwiDoJzhQfKQBhK+wxj6Nqacvr67VmijqGRCv8G3sbOISD
PTA8iJHBxiiDugysLKerWHIWfOJFrf7PVMqaCvbeZkUmxhynCO+posIIT6NpDx0CECR+wiKq3mBK
T/MyApmgUkZMONnDIdDT9SFmYQQ4tfOV7gU9IyN1wG0WVfSJ2NUu7WcZ0+xIc4GzoWH2yIfmxlfH
vQVYyjrsp8guTgZHMAF2KFhvCH+a/bDRWxCPawSXxv0pvI5P/NSLLGfl4qAWEEM8EdUZGREYpMtX
PsiiwoIhBESNnc7eRkW7fJHyUKVsJSAASPRHgMtDkHu8sHy4irqOEsXAsVVCaRy0sg09LJlT0adx
yrk2sVScIqnP1WQ6p0zu4auf5jit1/UXLuuf9GPSyiSOwPDesY25t6cnsih38D9A74OPho2zvsZA
M1owwiWatRiFlT0ZL4B0LvP1yxHQOteHSpNCvuwi1ypSZNamSBY9KJJYdWPY5JcOqpP8l56lswZE
2ypZVNsZAqcDIl3lzkzqYdaMemsYoaOB1JU8BeepVUqGnS709H2CPMzXGf7dYMDz55+6TwGjsPnq
mogkk3qtkoIVYA4IIo66SAAR/c/IX+a5ovupDaX5Q8uVSHxf8GfIDVbRZgGiZEW8SIvgq0I77Vdu
IxJvSdYtP8nnwaSAZL2rEZOjDbVLpHgiMuPTd6iNWnWhZpWGhGecfF0SPtz8weP65WOkHfKmEOEM
Gh1KPeZcLkj3KGQFrq+yeU11xsZORkf+rZ0qS9xaeyZIzCnVAWsTe1eBb+dme2JVhySFPvumHlA1
YrRrNnREH9CK0Q/9NkQQauWJYts2XEqx2M4sKCzksFAGm1dBzno3xYOKVlBjE0o+6EptLnMpBTjl
4RJ/2m4CMRQ9ifidwoVkpqqm+RWe4yZDJjXp7mU9HoI/K+NM/fUdPHuE0J84u5CkRYba6oBXmTXD
Hn/TDyECF/cuASPv11RCf86KNk+I4iFKScJsFdH0nwpxcT3sUsYFmANiySCN2AG5UMWzODMFoTWY
rqcxkb2zkALEApQu9qMoV90j1Er4cEns31+rdFiARcieCcyAgLVVEVIexkHi5ZTO8k1Vd2KCOW2B
loitNaJhrLz9qjcm/9U2sx81nA8cX3KDRVosuL2bmBoBvLWBRhEWf9xIOFtInNgx2jXHzH214N6/
AXixH8Cb3KYGcyKW0dtnP2X7fHAiiv2znSOk0GoShautlNlOcfNETUiGnnsI6fj5fZL2H9uqy9dn
eXRFxQ5v9dlpDvhL9vbzTb/wydNIrzbt4rPtJzwlOVE6RL1v/uY3q3hR767Bl/XenesStIeSku+2
GuBcWAflkqY99KMbztEp+gQSbNNCWmHgvcJCo0C54iK7CBd9BW6ICh5ypqPavi7nYOm7lDTCuUTl
aeHikihFyIpREZ7IcH2nhSraziJ2Q9OsmhdvHOqrjM4Z8suVjTfvp4yzWDtA9zhfgfx+OYdP1w24
NCD38vBosoL0QigRAWGM0ULX+4SBjzLdfWnUoDiAuU++TXDUCkSp6b/k4gNFgDyqN6RYLI2o8vWT
npr8F2uHFrBvCFCz2w6pc2f0ROp6whJ+ifU/chKqPnV/0JfqnAYatKikytRj32tE08u7HcAkZRzM
g5NwNQZBD77ij3F6rvRH5jlkSHOUBmdUZ7Yz11QFJUhQ04ctMEZrj1JCmVff7k7QKl7Fo5+ZbIWw
HwA85UE0mnH0d/Hd5QOjsKBruRK8NcrvJ6tm5A0MD3N6iq99gmdXLbbaIEgA/PqQBt51bVp7flLU
tQ6HpAEckSHBTSHE8Ygaj4V1hpR/tDNZw27GjTc1Gg5Qw6VrNVCEUc7VBuQsnOom+zIamuVlJ1cR
fZn5Zyuvo5e1XgiQLrg2AZq/ZPWNmv3/cASqMv2dDgQ7fF8bTVpfDCa4DwyCfm3kN56Iz85YvkkL
r16UgorIcEFGjR0RxfY9FsoGGTdA03mIxcOkv2NkB4Nfw29ZtQgrcOvlQvaY8v0pou/Wi3W3nIRy
3X0gKCJ0udivrxUgswm1zY4cth0rciYS/v43745CS9K29j2duQYAEB4l9PonUF+F2SUYjXlZU045
uZJimMh/j269PbHF7nnMAcVvKiVnNw4U9ZAwDKeUEpp35ruyFVbf5zLph8pFz/4Fib0M+iC9iPZz
FyYZXvSOQbk0a8YcvDiTuLr1qAe7nNt4Kv7vsZUoXpXZ8mK84hIpOUtVQ2v49oRIUUMRXhTcX1YN
igV1J4KEEmAJ6BkvXsI7tsTL9VVLKGdouXLuyy+nD/G+75iBi28P/7jGdXfK5RbNPab9oQfV9bgW
oLfk2fvJcf0KKIL4oCXiYLRGmnh0wfG1T86YMAf9BwVYlyo4GvEZmK9xqYw8z80TOrabbq6vKUdz
yVe4J/S1UqeOPnlJkNQ36TVlpAtVrrAvThASVSRV8alA3C7+q5xz2laibM87quHPV+eUN8lhVHvw
8sJM7xHX8ryrIs2boYkMaAtAj8OI9aHGlPy8LAsW7kAAIB51TKxqzbhZ3NqENZAn+ExAHy+D4HEC
mCCxluRT5KXyFme807I96ZWcvlutcPZSJcsmHkJ1NezElIyEOO2rig3ERRl5PKyICCSHY1ykiwHL
XIGSxIj3t0cCuqzADTwI/kafI5PSPqDmHa5m3HB3kYJ1pG2/NtVJjwAvGmtsdBTQIcNwlsSZo4hF
JbqiwpmptibwiFUVnWG/sNsmdy8NtO72iSPdGld2PVYsNSTxpUjb0As5gzZWO5FwTHeNWexge3x4
0se2Hg1JQe18ZfYe3WefyO56kJzkveX2zDGa91VPfqSX4VD2cb/Bqk7gVvX6KriqegDSX6FogWH6
JLG01YI2hKibRgoUjwhu4pxoyZso3vchbvEKt6FEKQVL50bw2hV2w38hNX8Pz42IgFKokw9Fravf
s29NFANPkeDKDXlDNAYT/lDydWoe59stx1KA2FtXoaBsD0NQ6947WU+XuZVZijyII5zR8tD6EJfq
+FIwU6B5hH704v1keqPUMmp/e1eY8UpSzHT8Wl2DL9YJQolVkB4NcY7zotV3+YR0Yzqr55S99wWc
jzjuXeiWCc08fWq0OwlZJg4Ize2kPEdYunF1Pc0SrFK0FdTISiOkYIt0L7kWx/H5jQWPqI4Sk2lg
hniHZxgHRT0R7yH6tHc4gXblOjHtMoiLJbXa2Gajxj6ZBSvWg4Xw18RE4fBKpQ7LXZoItu18/PH+
mwROpiixpd3/bBPmJjY7sVoy/r6EPp7Yr53RNh+7zSQk2BqpiC8VYmcr4ENqik+k6W+d36hRRr8u
SXhzWtj58lNGU0Z+Ldo3UUmqLCsYRL5AnjJaIQucOgQcSddH56UoZTsvUVo8lSwRUpW+lIrGnoOh
ZRrgKyq8MbmPnev0OANWqEaT70hyQmrARsjG0pxQRXVRCB8EYzr4u6b7eu3e7m2fsbKZVrnQtj8a
VRt0Hfe5WchKpx1IRM5BUuBTCZfTjboFaCleOO5mp4OgnXsIwfV+GotJgxJUYYHB7EL/ZwkBsUmd
cv4ko5rw66yMiGwsrQTZ3rmfwNb+DMKO+FIdygdjTTTAgsuYOXgZ79d7e16EUZPgPyo3ZLT20v5j
n0DhJiM8jPN1QvAh44O3C1KJAgCUXdNVj/IC661WXCCjaAzlcZIalyYrfT9WUd7EH5SEFIpRyRjb
dthdB2yLLBcHGUoxEoHLJSY5tN+Xv/KBd4akym35Ld/rujsmgDfPgqyptKEryc5bJ4Pt101o1Gim
LqreoG6d3IxAyl/01l2rwT/8QFQa7naGEPj+EWRG5cWY8PG7Co5vCHGRmrprLUQffzADMbhagCF4
m1EYMcG1jBqlF+40FVgs27Kz6LcjZ6Vom5ENyhhak4J8uxZgOO9uMeo/DzbNBjpxenN6UwkzdvLm
vTFYWPqwSMpXEpQCfSX5EM0Huibvi7w5L0dJmTMMVySFy9U6T8uHhDX9uqUFOwAvXeNm9dLlack1
mK9tWXsy22CzED1IoLCP/dTL6ON/hiSH8+v2VXMY9SCpDjx0E3+Wkeg3xfYG9jJJWx3ysWhRnhj/
bqeQFNANV30kZVqpPnSKb7Fwb+jNL6OleoQFUpeuZQQXy8Bj6IxQG1TgwisBwfr74tqDUU0aclcL
uQvTU6F+tVXGen5o5I7rAz/UGOmWbSxUS51OAQzb1srXdpTNLwTTVtEWzhV9crWEBFd7bSuVwpnQ
mxpuqTVlPuqvvy0lG6htNNIx6WwOy/skz9jKj6NLnyQxfc135yKae8SxzhwTZVLhiqSuwPHdstdP
a6QQAqzZt5x5QFQkmtcYi/+X1w+k137sGNKvL68oLyCRaTgl18UCOzX1I/O/pAW5k9vFZESIBvOn
mwMX2mx8waumHhV8+is7cuKJ4qKUDLUqNWXnP+2yOEDJpEcX/QGL2isunbVVwSKdAfUFBPWO1LtR
neMl54q14FOr9Ytbqy0Ok+zkoyrhN1nCzdO9rM/+kmp2b//JM6ZUt8FTRuGBnUzWDSH3dTBM4bQw
wvI/c0+t9nzJtg1ujBO6TB+zlmbcXjGP+0ZCuSxSn2B/oLT2WTWl2emQGSLcNpczeyyIlqXehDjB
e8PJqiyj4JtTeKfiPS0hqKLmmq1Nc9iBUaQETya4ENO2idMSQI3pNbz/fTXkQxG0G38ESqdzFKXH
tEwy6riw0Crdj7gMqxCRgVFZMVcKf72qiL7AFr4Fy1ko3zBNH/0Lu9wJTRKYDFBuQ8EnCavsdjGH
/sBYzXxPmFKOLEGxr201G7DB30EgzgEtlqwAYNm23NXeYwBF6aLCwRPzKzdALlRerIZYa1LrxswC
Q2ecxCTuXI7HpjiRTf0wAbXv+Ds3YXAr0rnY++c/wWNQ/qF69xGhD/Vb+2MG3/6HwsxxB+vBuAxq
7Z9vpmd8blwjI8zDIa0ETx6RaO1Z0wtRuYgdWFvR6hAY57q/JQERKfaDaNoLck4MrBlPq+Ir4+OL
+6b5Z+JSCFuXmrcLvaBTBxzHKMCfIU4y+Gq1yxL8UVp4SpoH8ro5BlHbHWJMsdSFrQbn8uoh5mip
oCX2W7pw/izHpZXKZvCiJGBZQgvYIA23vZaJrRcW0pubT7vQH8blo7VwtoDgb2cpJMJxxoWiddib
uJwFO5yCZsK4qdZv/jOG+JIkmRFb17PaZ+kpWe2zP1f4H2rsuSuLPQzB9fO81HspDIP+SAts6uHW
u+yoFvdN7VqOJ2rAiwiNoYSgFDmt8e/naNZaSYn3ppMrsPrlyM8NY5p+tlq4WqcucJ6taE5I0i1e
eCz3geA+YaSKysKbATJQKHTWbMKE25SJ+cRaQSp6suPzB8F6/2NJjr+KfhWDWXdLR9VfjiMWJigi
0AM6RQ6RVAKhqOpw2aMzQ6h+tAX5MBHBGGK68Ont041qhoS8d7gT6fCOkZVMpa39XwT7pOnziJp9
riBsT8hBaOUHd4FMGi2NZO+0gbq2VEv780GnX9BDPXSlF3z8NJzZR/0f2fMzvyIj2DDHkzXURo6c
4iL4QTSYK7NT0e6Cw/KYV3Fj9rnTkm1Lj5Cwj3/96vacVnVFHQ2G0FlyhYcyBKNowr1PB3uW5aQy
sAAHHq3u2pVp/xAPGF4BkJbUFhLRkpAHKRD+YClKz9E6UNZdz+fQKbxD+AxRohvYKy8rj0Nt/2ST
MmQAArJUq+Ts2HT4Tqhku1Uk+doXqq9w6GDEkY8Bt/AP+kOSaubvprcU2bKqqRxQXpKzoZisp2WF
NMb+p0oDSncqsY6A3nEHAwQtNjuB185fRdOdA/q7ob3fgTLlg3PgAwGqYv2vInhOEn8SuvPGh3ok
foU6pFoyTxOawzUhKUYNVmMzd23XIhwp6ZBCtfPCADJEkiz9UQloIDi6aynE3OLpViys98lgjn/x
RL/YhxDWA6QXnRJsXumx/u2MqGRCjTNh+ifxuvJkQ2yfvcyvA7j5CA4PkmZugjAVKl+EFhXmei2R
2/c/DBknv3GRVVKDXjABWZjy6pmY4WDmu+mp5XaPeajhTsTiMc11KmLolpq1nQzJstviyE//B0RS
yka0WpPPh9SFxWgBabmEnXk12NLDpp4uuSVJIRzEEoKq5YKo9PJpsLl4p4ZeLn48HAUrS4/3NbLH
D0ODHMDKGOFiSTo3E8JlRxUPaJKsYNw4zzJ6UJQa16MMaV90uhd73TtCW2iVkVqud9sARNe/7Hw+
ynOed9h0CQBKere9DWxUw2I/gBE6kWfLV7Y8XEDptygm+I7/tYlGoQ5mfBBiE3tijHNjehgn/ykw
c8Q4ALPWwn0tHYQ5D0M5e0K5U7MFrWf+gOwbfrqLsCwLnBFVeg/SWxyNGquH6cxdvaLl9sgSpzWj
XEwIk2qJDuRzKjcntxl8qyEwjWJyAXWBRFnyFLrTGQbsNJmsyD/3eIh4Mk63Y/00DrdDq5LcBmTq
hU62YJXgkrZ4diDHSUxAMn0VafpcNb1/m84Wp0mq3R+4tgswI82ViCx/k5+SIdsI9gP9Ms/53wHH
KIhRFt4CymbFZjoNgtP3mSCjwnW/RtN2oWsX2dH4T9UKmy17PZNu2K9lpZSuiv/FbHss7DuBduXk
M2fGPLZ6NsDSnCQxFV0X+Tx572Kha/DRZiEwY3yYlRUe+FmucaGutVsGlUfrWtmVaY/K1VFvAaN/
BCm8+KDfLD+Alo3xqUgmTqaInXAK4RSdn30sohpITjgE9cRQJ07RlZBJ7JhfXDV+GU/MicO+g12T
hAziZROFXH3bsYds/++Or2iUR58Xi77V/IcAJJN6F/L+XNcGsVSTMHRsxSRSDzwtS6OPEI+Wu6EQ
ydGLWFZ/HQIqHTo55PmkrswHzOyuGbjCvJbIHetkEbyiXUZpjVdz/MluJdch4IjcW8qMOs748ll1
c/IA5nke5BCxTlE/KFXmxv7IHDN+HgkKBGTsfPH1PZQZGKG2YAkmVTKksrptmJvi/echk6TJ/z2m
4wefYDK11zznkw9jcrp6HHcuPMeiylBfTcvg/Zw44IE4myA/kMVpyHqrvaYSYbNdPnWOY4DEI0xu
sM1KQ1JbImCI6Xvqjefx3O8vTpA6hCclk/xYqYvYAH1lo2t304yCJkR2t08R56PlE2S/pzVnNDW4
JweCNiedXcmv859m2eSYQ+nkmZeUlBYAFDPEqW1AwG2t9mqOOmg2JY/o5zrAsIyzJWZrUjLnkg0I
VfyRJusp+sG5+tCTo26pKYpe5VNNJ+4zPP1CJERJmQofOQo2MfTPg5V+cpuTCwnpKJqxu7zUnKJH
b0wbllR0uOs7VgnOXjAk0/6DeuBu86AWnWGmJMeRX7P2ZGelXp0M3+F2sOwllwBy4nWcTlBJRJA2
xsaHzSbNCAUgTdlAZufQ2ypdd9/EFNXQLmCrYKlL7dgeeqXpQ8lVuK6LgjYbnba9iHrsSHj8TIc7
VYTs+OCevEsqMQICVnGFQ9hSYTyj2b6+QTbfLTDD3hkdeZnMU4TjH4+DfVtWLgvqczL4c3hP0Tki
+3fN3d5mtTQmx04/UbVp22xaiRDcswWA6piZ79ewU72DxzTrmxqzQMjd697bptu+aq0LjWu1RHwo
Y4CyPdM6Ydid7rt2DFK5ol+JMWSgq38d/pIok5mExisGW1QHJ7ogfJV/1S0ISJwoBHh/ZHNpajYx
tOA66Y7grITTGFn9bt4r5086MCOf5QPg5pxXdi2hrvwFUEFzT21VUcUgV6ATxaqD09d5RpVIDAfn
WmbHXt0mEStOlpExb2XoZbbk+vp/GNjcd9O02xCSz8wbVvOB84nDrbfIfVu494B/3fYkCekCXNmX
OAmp94yMOybQgv487rMZG8KHP7nwlLdpIcooVzlWjtdO4KYQCzkqnVR2UM8ogYpCv5bgTZwD7WrD
NlAwKwqKPMm7TnwKyLoJ1OsuVv5ETuIugjXJP6dmpKiXfy6j8Aln64SCIgh5h/RIdWjMPCGO8wCP
ptnUMOiqK6e5UByo86R6d6lQj+TF5b/+WgNACjCJwyKv+jsqLQ09lu8MH5gUsSb0ZwyPS5gpPQa0
lpLdTb9GIVSY7FH1W4/aPyW3dX/A4Lx1XTagi2iCedZgPNhAgr1bKXhnvbgAlOdefEQLT8X/VqnD
12YxHxZRM7jl3ojY5WQnstfRIeIAQUbY1igHfcibINNANUu1NlHJG34GtPSUp+JsXK8BZZBQK/9Y
/gtLUmrha4y+MVHqtNRHhcvITOq+YDkCg3rolNx2qnb2u8RGxYWns926WHL/KTSxlVRcyMrNvQlQ
L2IdI/79Rw7x1JLCt412Pe28gcVt7Nx6ZKwdBwVENljmGyD2xb46UxVvdk6Bob4mX+zwL7zlSdEk
qYXRYfI+clG06o+xAMgfI22HvhwAPINEr27hYitIgj0F9IjW4lm/br4rc6y9zQa0w7t47uicb3rX
TWDLFTEdsIAtiRSKn8946S67Fw5uPstb3EjTwrg97BPi/8W/mUgVGYdrXraWhZ71edLXVqgXc/9z
INiZOuUiAI1oQmZotaSE6TFeDh/rjtIdTSa8eq9v7WyO5FlAVeumn+v+SCCXLRnzfjoydrrNhwpw
mjJxdMqUZo9bJ2xHBs3jm5rJFWz+IUo336s2ZLSKXeEJZrgKhZLqPmN+xALky0jC3R5DB6GW5ALe
d7v/Zr9FXXzBMP8iePZMmC4sQZ20W+VJB5H2I7ZJai1ZznXgtUt2JEma8mLjJBNtNrmWE0QOyxP6
sYNJ/9tFQTqbjKAM9Rl0kERuZxK2+PrJtGO5IkLCxRlofZksanae+E8OUIgVnL29buvUDwxTjSDH
U+vr7eUP+alp8nk6s7L2W+leoBPbwmHKrU8roQv9/p2hOfQNogrSn3Wp5w6vuWXtkdcZE4LM6wJ3
3hRAIzjhzDwbqoUuyY9pikaBn41Hp5ILg0zTyDLSteopsx2LTjrtA4JyfJDmRi7Gh1g3lycEOc53
W+H1mlHEF1E1U461ilIFCUHEt+vfKOfmYWaZ4pheWecbWRYwyAZR+62wR9S/tcAHSN8wAYJ7AOLp
yDRwDcHUYHfYzIGRZ2l4BhvuzeH0Ls0aFMWOfr6tE7cEwi5mJ3XNy7ftUaRf8YOdAVVQAUjwdG4S
frUfcTemOybBasS+LgHZNvbrHnZtscAet4LiTp9H3USyjuuSJ/vO0qYP7VlR8cstrlzYppCtyQVL
/lClCzLCUMEEBhEZokPO2V+ROze6WTq9MgIgpBJpAnDuoV5gTwoR58AwHaT+/wa844JlH2MDHN6a
EBlXC1VTt+dlsA1KdraEhjOhbph9o+Ls/J0+EbnwRR1gnT5q2m7JOrVKVztl7a4k/1I1oIzcX1X3
LgjaMHa8O6D+DGu8zgDhhwVqqH75c8rteiRb/F/x97vP3ld1zyhwEEnROXYg9rF6taAD5wMIfBki
G6HVmJL9c7GfG6oFgEclyaXYpaGiH6iQb645kmZFgE3KYLYhJlXt5ptfCAqrVlEi17g7lyCQXoAq
FqZE9pZ+c6KUI7oQdaSplpH+KGxUJZ6SAga29IgM2ZbcgBkI0KI+C8RrsxQreXYzTHw1UdtiXKe5
jyzry6xA725M9S9/H7YOcjBUTAbBVIJqh0kGM01dfiVbwfXPxpMPb5DqvGjVzQeMYErtcUGY/+AG
sO0imLgzy6Pi+T69js4w8Tci694pSmmCKP/lD3ojU5S3vMNMEHccj2yujkw4qhHnAu82oec4SLVP
Y/XbST3L2ihf5tZxZMd/7In1bbSEyGIUwHnM01fT2ivNwO+kwdcpEIUgXS3GQWW5CrtvuyfAIkNu
ctaWUAO6yMSobwko3/vjjww2IQoYWbWRkJn+8b8zqB9Ofjuo69XvM/3rkGimg/xSmB+AMhbodZv5
tHpt8Zu29U6RWSKigVZcX8GRBES9GKExdv4WHLzVWkUdZUbB2DrmQ3TPUtmUGDBQxNWBrwSFK4RL
3uvN9qD+MA0DbkckPWx4lEfxLbIyBwAkqt0ybIfB3sitaGVsoMwAQKWSVK4HWl0MdBMtpCw3u9wk
oJmWnTzZ9whOpoBlzNc2qMnIvOwai4nXnzuQTDaLC6vRAZ821ZnH8cmmlq5cnI+l5D/BKsj1mgJZ
bCMJi1hr8/yij8p0j9FOPcnqbf8L8bhOcqGE0wQBTvb+BCUI2YoIqOs5W45hIMuRZs5MxyZNeYu4
DhCbLnn3C01ZTfuw8+pU5B24CvqR4dNoMmU3YQoSK2PyH5ZL/N0VqZsPe4AW8QZHXxd4zlFBQe6s
PzYS/DIVeRV5uzU8u3PLuPgk3qdAtLEvcp9go7AjheZZIFXlYMaXDoxuKFGLloxz0IpJDk71gWxj
2zzDOwtIV4wbI/V0zMSmxJq0IcEyBrzQk6EB88QTawhsGBMKqe2Cgczt2anktdrZIKQ2rHiaLhv8
plca/IFmoAxXY0COPCaC3UAR0ws+irfXKOOAdSfsEy+TuzmrIm+O08mwIIT/QS5sjpgJMUZCK6rA
w1gTRCpu34F6nB0y0xVxxW8d64mqCn8UDNCC8fqCEiypIQ8Z0EtPSFIf013FP0QShUz02/WSkJCD
e7ospkE9GeJsJB9iGiWD5A/KP0dEOQyWbwhk2xr9UcRVLlgOv7nfWNrG5/a7AYmrIhUhwJ3fPDZb
7JxT3rIM+np75Y+Phi1sqYe9QDotlOI2toOpTMCcwz8lofufzh8J+/z2Z7nCejWadLlmvoyGVRNC
76H/KWT3lYTi0OXy6FyLT/mdpDTL5bq5sSK92uG4rI1qs799N5HrxlzdlBJZ5BWUH8b1fFFPzazi
WaWfrPe45L7TrF1XxKvVmsDRraUs/NdTvCPe9EnihlEPDJgXC5LbCCbCiB08ggvJfMCyketOBVvH
gjFtV+854mLT36XcnDTusbFnXomRKzU5oHeK37zvzdhi9mrNXEIQYKKoJBp8/mC53MxLzG8T4OKQ
scfDflYgRlJuRFREPKjyfUxEQnGtCAK0qm+TqhztCYRByv/yD76dCTdaB8XXiz243Wji5FjHVrzu
CJH6m1iC5715ICpjjukv7aNo4KS2DO0aGqkQNVoLFFe4w/roJdl2iPuvP7mKRGJFic/Cf6JjRm6i
sn7Fok09eMnI1BU9lvuCwWe0DjeVU7UJ1UdKy1uXx/tT1L3AWvRZt1CIbZukuVN8Bx6gY7x6ZsiM
sMuQDEW28vkk8E3awUKlRwPZLJ6BxPPk746rEaNDywtjAOspTvfZFLgKA/lmJ1MoO1OEx6DwxxGq
2Fa7W9KZrMTE6LyACKBorZHyD2Of3lbdY1yFNPVLJy3flgALg32BsS6NbtZJYWATOToDUAZ1Apci
lV1Qzq9ycUNnFqkhg5yiYOoXQ2Ybq+VtBteXm9fWMXlcXE9uKSQi/eo9KOtGivpA79P6Y+QPrpKl
AE8teQ8yIF0e8b3buZnePvzP/FFWV80/R8cKc3fI+g3R1EVSnZ1cCOftnskOFNxLBawYeerVTJCX
ObLZaTZVnK8tvaZ2HAFKPIL82ifVuVkgh+eqCCUZidZNspIkKQmS2sfs9NvPD1ZUXrb9rHmo9c1F
+Z+r9jBdp8qWKNcq5tLRaxS/kO3ADbOCvrBTis/CK/Eg+P6zgyEk/sXRx6jnrLfJvyaK4sqrr8rK
f+QiiCqJcebaOBAKLJV1QETCQNP9Cavtmg9qsX3OaccOGW2q0QpNT4Ns031AyA+31jrnR3Pe/4dv
l34q0Qc+mIOW4Zbn3qzn+fmZHKZQXHdY0bfU8Q+KKqoq+AY91e3lSVonhoR/oZQGM6b3Vm7d2/Uv
riVSFaAYaLVInRYnFGAA1gPYfGfhCVNFq96R3c2/vYEYRZWXVlw7wLFTSoIddErUtI+nisgpfdIy
eS/0Eq4gfUgY2mAh7rcBftVWm8/Ay/FO5ZlrAE6wepqyGma8jeQrYIEoUGFowcPaVkrdWQ4YUu9z
98X5ZCzowzV+okrC+BR0FLYW9zRKZdJIR05Nn9v7sxWH27cboGPxfZfGujsL6IEqIMUbOP+HthRy
/yPRYUegA2vOsqxONtd5PWYliaLb1jbEZoeCtLz6aYhGL1UWd1I2cvxpm92J0S/CN9CkkHAFfikj
Is2CbC+EnC34XH08joJk44+5B6xCtBnz5DzTQ5rCAkD+uooIFRdAs8CaXoHIwdOoEJZDA/sqyiKf
daGCr24dDAFgeQ+7k2w5xB7Thfmf0Sm/U2XamfoGr8gEfGG5mJx7cSEqTvA4lGG8isyVO0o1yRdP
bBUHY5SyC7SWsHchdI53R6MKPGJ+y49cug/LoLJ0mfOZsRQCGXKKBCkoqE2Q9R2ByvZhLUhsBH31
RtH5zKieTtckDYWIFKrroPe0N7qWr7T1UGwrr9GsmSB0VdymO7Wy9eMEqzseKYTBTj7qQ72LOXCM
L29m7w35IbIVhBkilKV2ygRGtjjOfhRrMyovukBVSlM7Q+TgW8q/Wdslk3IFhbPbjMb3U+vozCC7
t2k8wtsig3lYQFjPPlnbQhgMOlIKnSYqEE1D6yPz9SosjqP1hX1fyw0pWvF6arPCjispAsaiiEFO
3eLQPh49Q5rwmCeqPWViHb5XXBXfzcsuVnPzjDYsVv3JJHxbtlKJuq+iNvuI8czou2JWrYJwUjng
Oap6BLw6rnriy3CPH60v7fP1YKKMd/4hRXGXzpxVJG1xf6Y1Y2kiFRdHWfqPkN9xCS56zbjj4iXM
JLBtK/1k9MdYqWrulHh741I2cE6uKjEsGoi8bTjf1QLJEOlhmyqCFcfvTIiI+9ZfWDX7XFq7s0Ad
1r62y4LzdlRGG91omwEe+B4Gx4ZJfKMbqdUu3huAn/qlZIcab8u1Z9JhhifL5aWpiC2o1AiKWgM1
M3995oBN6oJcskVmZU6opSPMYgXo9MI11vOrvxN50X5Ywz3mJMhFXYCeSOjmQtKcGnNfkvJgbof2
XmTFOjMVfiqsYfid8Za0rGHFlpHhwf270q6dr524YYkUek+kQy7hk0qg0ubus4aURD43wA7Lo7/1
I764+gcOIH535Pgu6Gq0iiVubA6HdGtHL6ZGWVSyllGV0QLdjTNQ9TC/hP/8ct+yPJS6sJ4x4lfd
GziYrrrbZn3WVB41nQBTQ+0vv1S8ipQJQLHgAy5Eb8B6OhsqIBKrmR1xUAzHsDLKdA20c8VLkDVf
s94TyU6cqu3FCQtQmpCY3QvgiV20QyVZ8cQgSNUGP8hNZApXHHa4wUKMU4Uv0LfT4wx2KWPHc2Kw
X3b+V/KyIvbafuSJfCeIVR6KAYcBsOUoaK7XR+QjX3dD0OtL/vD9HkuOrOekAfAitdtt0X40qZu8
n1tcKiCqc9sj7jtxHXis+NQ81jwAWfC2GHQFN6/1k7vm3q2dWPRkobRxJRXdyHJ+GlauqhmcYjTi
IMViSTTYjjQObuJUWcXjWjmv8cHoB3TNUb65H36/lvRFlqcTBrZdcjUjaOAW3mlrf9NzIXc0Z/cf
rAmDvLl9EKbqjubkoIUejz0w6X/3yP3rIdw0rDFAzsEFig6sPvne25R+K4BIGBPeuO9ocqoMf/jb
3IbI83l4TuiCX2b2qzQ278AbN/UzDH+ZIdGSXOoxW22BTO2Bj0CccCauFqFMusce783g3cuucece
rMwKY2BMXsvpAT8ZJdmCyds5IbeHYEq3c/iGY8wslLX5ticIcs7A8wyubWaE4AHeqHDhDJvaZYZM
UykhBb8cHHSHO1HtLsP2zUkDBNw6X/gEl+p2STL5rdNhrnidakuub5xV6pMF78uBGXpcMxblywnY
Ok0eTpYGfWp55rBE/fsmlvz6t4A5SGTVuDF1Ug7t+M/rLiRlvrkaIEb4MYyS7YHBl12LK9EqHvUQ
jEmC+T8XJbQiWoxOWHYXZKS6YbhsW8WTjzI1LWFm83FWZGiU4USIVNn5bcyEcVXegK63vZMxBpL3
ZuEK24LAgFabP+Fj6f3gtwh6/LZ4XtzCry4SsDGaczB29KWuR5vB3Ch06UYSiMwtmN9ie8slsS4+
RjyW74IToMjqh/pLA70Un2Ox3GQsdFi+Yckyab/LWeiazGnNqP7ox+qPwVwxbFieCMSo5Yw0uHuA
6e2B0VvzVib+a1MI+C4UId4EenUODVEn0ONfHaELDiPL4AgUEyUqva6XEbAN4k3TqvwxUb7SwBMZ
13dDy5TCy7+BmRbol6LfNgKCaZxaXPDStohi6xLWAu8w1dCFhUwcxDgU9wofMZaijR/br273nzEk
8eZyfeJkLk7F3MjnkGM3TmxrMo417R2aeAz3YDGxg6Yqb2J7AGnn0s/FmP3kLLx//6pP60+0hmpF
lMrtpGQD2X/4w7TmWlGLUfwnhzKjcenvojIvpg0DmqqOSDRvkOYlImIIwZQZ3HB++4MqQ1vmQMuw
UjnfsonjpDXBQhYud6rZnsUR48U8GtIkMGV0faM0FAksBSlYgPNCOS7t+0CC7IyyNgpBFm7Lt+86
/DllEWK/puSOcKOlDN35+n2uiKjvg8wtpemELWrNpxudblXkW6gNp9ymVXjHGqgKiBHoBtsxTMuM
0o7BYdoq5k4eA7LQlZA4N8rRr8Pzq4IwgdYoiseUQs9uMDTEhu+l5yIrX15pBWTOucs8a2aOlM7v
BkE7ALGYvJuhmCA5G4KM5fxwjYqEJHQo2RJQZZoD2XHl2yctds6eVz19zVNgkvXGCvM71AzKb95p
95D3uORgt2Y5niyx4AgPCuTWINizkVdnqaClbYUY7GMUjPSnQsSTBdqxqWy/R/DMafU5D9BiHSK1
a7s0N0dcaql8Pw5mquMy1tKCx7qaQRFe18HAF4xybQQHjsMgUwq7lmQU3fxu4LP+V/U81W+SisTk
jfEinpTOCZ1k5l0FrQT5avrZXXfONHZN1g5p3bkakVXglVxHwJuNrX8nGmRmEf0kqBW5kmNs6qbm
eScrkTP2zwAvwC2DwDsfV5d0v7l4D/jW5Fl1cGCbIdf2tzj+9stTM+GqWoeP1xtSCsLyJt58uoib
PUj7Lk9mhlk1BY+Mzd5Wa0PJ8SkucOSd88nwR0mL94oztoB6DLcnMx/PUjdSvwmAz0vYsSZb0QZb
/CVP/eZL88LlljRbF1JvGGUWSzB+7KAIN93QQmaMJPZzGtP+G/SDSkVySCZ/XEyMXN6sUCR+cNMJ
TNhm9iO8mhS0A7PzFzOG35toxINur0RA1ZNmO950JRQKT1LM7Vph6HePGcRjGnpUeEy0aofStIbK
ABYQLYKVVWvOjWySVeju2mW+YqZkX6A6pUQqFKg7lbXhXYWyUUqGv589H519STLeb4bnSghCNsdf
LCSZNrqxfaOXs9H5KwcT4yRDLWyD/s3bPphFEHkKoUjBEXYsZqTPj/n9pTL9EF0q9rGmhsFraiS9
gD/YtzMzRVkxZsD5x/PjBvK2+zNxeBh6tfW/fmtBrVJScqjXNZup4yWPZ0WaOQv4P/CajxmyBRpx
QkOISr05/JaPAgxlVuweF0C2b51JXwWKiiUFcp1GIpyY8Qthi5fT7jU4Hcd+bRQc/T1DQUn1U6V8
eGBU2Z8N8SYbozd8LtCr96Ntx4iyJuxiC4J+EX0yWghPN4ZMLntRY7+VjUxtQ9Q+i+fvc9PUKJT5
JBOW90VOvDh5FsHOKFFYIItEP38k+UdO3GB/PYfGmKMgxuMSmWHd/1pKdTRxml1+9TKQkZ6mkDrz
qzKWZWoBBmN4VhlWiYV7E4pDjQKz5bmM6jCvxA1pb9NsQhdRBaNAy+iyMYCUiQr2YgjoZvC2/322
NasZ1AFVD7k0Hx6FrgV88TsyRJidDIkpfjxDe3dwnsgb/Q6aYAdPIQgyfL138MqpAS0OK5R0Oppn
bQbLGiCcW7PqatvoGwofyTPo8AkBt7EEx8N+2yY0b6d8lxj84Tn5NjZ9KryKoze4M6Cy6O3HJe75
TjQ71KMdAXGLdbShjECsEghxf19lVAgKy7KYJG9LBAkonr1yKLFxDBnq5TKTv4Gzy63M397MAIA4
Dlu8IKqYfzoATNDA2YM9x4GX4IdZQM8L+i/8Vf+iZQK4yzaVG2OlSMnvaavkVvakKmWg/kJ2hLwh
auzfQo8BTZRKkvvQuMgtJamGer+4V4hXfYTMpo0lkL6tAAWbUanVQl2tMBD1w/cIRmXuAvndmJNN
IJtt817xldPjIH4eMocHM4Ri3D4qv2xNjvCup2P/Tpdvq/S05dSbH0pg71oEY+KZZqwh0lVoX78l
JDLvnuueXT5zMVLwPpkKSDdUbls3CaG3M4cZ9LSdLPjHnODShRVhyubx58e7yIwrLVQL9a4Rg6uC
hkdBAkcMGZj16nadVr+PH/wyLXFYQt9fv/5std5rov6akNYde4qzbnTFNgAgUVMq6yFtrUbtl3rU
nUIZPMnlwzojL30XTLpzWv6sKpOLawh7hq67lHN81Kb6/wIAOYjFTn7hUIgKBFfrMgjd3SNZqodM
h6gM1rvWCr0oz+LdIrErH7PUXG7DcEGqc3ePzL0hs7dYs869SxKJJIOo1888lPSbLM4jVI18jjNz
+8mFcaU6IVqXWD7bm00aq3U6EA2IaT4bcREreY9+kwV0V+qk3cCkWasIB9a2KLnheyaiFXFQs/uy
NtVevdnYzwlA8yoiTkeHhodqu1DQgS9lFuhRVWzev59aQkuHG6wuJPkrT8oGE+44tWBwqDTWrGwx
8Kc9dBMbVnKWf2ulwyszknuUxwZyBVNNUnem9fysVi4b51wrkAKL+CEw9C/wsZBjFWRMhFOvlbC+
M3EsQ4i4PKScXIdXOP8Le8Riri+mxvyZktxnW0ES8HxSwkww0gHGVMilsEmHXUPJUibzqtRR6JFf
gRFoJ58OP6dyb8UjcyMWz3okJhtbdGPgPV9yD/lj/R4Dw119HzbwmgLnFBG6OPEXM9hQ35HhBVxU
M6M9sKno768ifZmEegJIRaSMZI/fFVXjpkxQrIqr6wmTQ+77BarLaQ6DY2wqo9ro/5Yont0DQ1mc
nGGTeNzYdirsyURVOGnzrOYzelEEeUJzjyFJd01ob2miYSZxN6IoJcVLH55ovt/yGaWCKdr3Do0u
mTxsFjJLEDw7o3d+tRKEBgQDXyH0eOoxeIoD4uMuoXpg97zjz5ssjyjYWUgn6g7RbHDx43D+6gVh
gvtnIMu07XZFhMZun4VstIZ6SOBUorxJHITK6iIggF2KeGssUq0RSvbSp5aBhRfhr/M/IHuP31Xp
2fmNUoKtoz7zBKTxU9gtkGEpWcrQWom91HM9n169keFu34D7wzihO35de/Q/M1FnBxGl7BvoL8oq
R8Hs4a+Y+F3AWBdjon9Ro7SblMcuu2VH4hU6EfNo0Dqz9/hKdflnwlAbR6fVMtR+jbAgOxyYnWzR
xvhc/G4Un/203kF6KBsvJy1F0zVJSK5FcugzNh6sDvL7pCGvmiHwuG4iXkjtpXgwJGJ9sj8ipezn
IVa+7lxqckUzXmiC1iYftvs29EIB8gvXV94tZproakCLby/mEXKdK8lm2Sh4bFuE1dv6M+1GJ7LP
hjy+QTUlbKAiABNqPWqIxjLsmw5WJmkWtuymTAYhSIcSU4MQSwp427bDmrkF+KHr6CfDjLcokLbK
Wv4Aj77ZZonlTdOsS1BFWSnQ+rgen3tV/LyCej4BSZONjM9fxt2WK2DTXdKyyC9qN32X32EOf6SJ
YuznfWnlUZ/iLdt5u8EJBmreJA4btSqg2d7AWvtv0tUaxN9iOBsVLOTEwNuwYBvBWd30YtocSps6
VUqVvYDSz5+QcdMbqpV3ze0Yxl9HILx+QMySu8m7OBzSZJKa43L1tKFjuPVA2O1V0I4N7rEOLMvv
vJPBdSOPr/6+KoEsO/7oE7RxQRP58oKnI4HbVXpg9uc3im8oSIjmctlmmFYXTc6KzxUkCLdpvxcP
jGtvB1EUQhvP8dnXldhA/IylfDyPyRGQDZpGbA86Xb67GDyHb74MkYt0P7yxr1tFvY0KyGSBuUQa
EiqsNKUJEi1qdYWqghx3iAqOCGAn0Py4qPwjovI590vwpflS/1XQ+WAJPM/wujXMHTSVvyU/HEcL
LXp/w2vYPFRWAWu797OXb8nS6o01qx4k3NUtjIOOxDUnj2ZvjUHECgoPUx3IO7z3cs2c/1vghCcI
M5rWYXKhLeTozcXZZjaWNhMZt498eRPBoZ2ZVfMmX5TmpLHCZ7p26jerjMIsoRG2Aqv9nHW2CRvL
R/bTUAIgXBoCO5kJXrg5E+TqfoDeqbgl0wlGV5FDIrvXIoII8AAYPTth1pR0UGBl894g1nJEsavY
zO4xAgt1ms9c6b+DyAcenFYu8GD7KpXTXrTKXL7SZfDuie3I3PGjr75ouankToPAcGC5cwHSQvgL
9UoYD5igvUbJmV7WMIkmu0g2brNKBAooW445DacZW7f7NfI/rAVaCQMCCm/rRtZ6hrNh19DraBlj
RiHcytQtdMvhOkYBSYeJOZCDY3S6NHKm+YzbTk8NJ5PE1asA8W84qPLAlzJLWn3BTiJ8lFty9NkJ
zQAky1/afbQ22KKUF8UguFbW9dcanWv9gau/J4/gCpvXSxMr2rsPDosYlRsL9i3oWzGJRdWqGZoD
qD9PzRpB8wOe31bbfmzgT5lTEnng0oVStEO9y86v3viF480+QXqQHw1qcaIlEdbUZv7yDQGdzi7L
gk87KV5js+xwyTKFNFXbeSENTke34bCjY/TKLK6xeT4Jkytsm4HDV9r4PZHWCfCmmHWLT0AR9Emr
wtScoIRXfNS0dKXvbG4D10hZeGGze7sON94mfnIcMAz1Sw1GknCp31yybWkTgle7vgSyAeMzM182
gbgaS7R6ZqHYV/fBef5OZYVuA1B3/exVL/RISay0VageqFr6D+47IqliZ+D3bC7tbAujjU3TLDME
JniqDbh0wBVHsfTDa6w4lT6G59O6+pYjb/QviaL5ihdAwjU7RgDz84Gn3flnAh8DIRiqMXAfqGgw
GSoG91dE0swR0yXNk+wCiTkHRZAs9ckEO4FFz1UnoeY+3fu/Qf1a3i8bEKnC7MqBlY2pQZQMbXFp
3Mx+NMpYsyXc/rIKxGOTNQn3g5cSGANM7rtKaSbJ/FjQOIX4A5RtLkMuAUUGHw4cnHokfteq0epQ
LyRxhRAdOwsmWzYVy35ymn/SzRzdAdDX+5OXUl202ZYQnqUs8NU0+N4uu/EPYn1StnsXUdk+QNPU
ynjbzBQUmJEdb9Znl6OwiegvdXiAITG+LRW3fbUa2g/5oN0l6UUydCcB5P1gptovE2lG80i08yrW
823eOFyE8J0ndegkK7PXjbmMuEQhh8mncs0HCDHfxoquxRY9/PycnbCH++vA6KH4PZZ+HMyj0PoW
zxqnSydZztufDpIa6zdeQdgVEbKyQHl6K/K8+kvUuOd4wmmMoAZB38+5VNCPixNzqUvvBLv4gcrm
kJHjJZV753Lc6Uu2sz1qlA6pxFAaII2u6OOA3SM4f0ELKjFsfolmv+67bDZVok9K9OrGjuajXVGu
Qo1BBjvrNXTc4foxWKFxYZv2M13IIvTKgGc3f6z269+20EyAMXzIZHY73ppH9+ROF8Nmfbi9Gb+X
JndcXDrBf8ZTvvw59O62ks3kMChWj8qSCMhyLhfaoDusKNEETaZDsA7K43q+ly3LdcKw6fZ5N2ZF
HR5XDRX1y06gAWMgBo8RZ4IyA6Gc4CdSKCDDzrCPGILyLcCrdydMyTRek37kUCR3rTVYm4yZyssQ
pWrjWBs2ZxpL+pCoFVwaQ9U1spmXS3qLT9DKYmGFXSCNci/fX5AR3Lz3HWNATPOwiA0ErrpGieqE
QXlzbE1n3w37f+FeWD6Mtnav2IxKyqUTU1OX1un3uprocgxL0T14bUQviLu+hmIavp4TJVc1y//q
MCnlMWeDPkX0YcjxDQlaD/c8LDpqsgqKjTKm4K8sZPLgetEsl+wnctx+KXBryWrplPqkYT7ABDDf
R7rwi4PVCtOic9KPdZ53uNR2vtxVhuHF6XydSe6aOXhJ1E2dsNz7tXgEHnHDS/yTwQQP2nYfmoD7
SIoHi9SfEQD+I7m1SW7F73PdUACZqQaLhWdLEQ0t0HrtrKEtH0u+IaUy/7lHPy5W3/UNbV/2Mbyo
NxdLoZXDzAQe6ouAa6Rx5++YBY/srW4nWmUhXcp0xdjTZ7yPn20L3B/sBsw8XwKzAEBKZypv+ylu
gpqRnk3YZ3O/EQKhU4CGY7ZGXFlcsHqIpXgH1mJHL4mb/yJJFHg1HoKY10Y+Z7QhRR12yVE6P0+g
J7mM9GLKMhGybnEZmMlO+XuMoZKY1Q1g/5poS6SV5Amc/bFwHEsLXGZRoQETsgv4P+PJzYLnLiwM
7iYeNEs/Qx8f3O+Lc55I8M8QK8oqolVDaBcuu/mX3X2A9CR0SvTyxTj4nU2wPMhbK83E0fyMXAv7
zYtsmJ9Xx9P3xA0nCCHuKTBepm7VbCvGRrG8HvI0baJp5vNEKD3zmUhIzdqxUOunSh41YxFOeo5h
PXalPLKveYI4NwG+KcfBDay7kq0fKN9wbOiuISQaTYTlmc7qMzwKxMZxhXkxMZZYp9hZaHa0SHYf
ejRY4N4dn2mWmzOfCbbuiOSjIVT0H1SZ2fhADPAgSgu5jj4VSVFXyW3BibFWhJTfycXiq+BZ9vE7
rj1Pf3HnzEifKaKGYd/44WhZIVgWU2Mc5gZ4xzUwonzs5kT+W5hXWIYUd2e5ysLl6PhkjDiJL/Y7
0Rka2WwM1NG1AYgkklLke2id9vFbAp0p1paZ15iEOeSKGyV0Gn2KkOyus9C0mNucnDpZHRPXyBIB
mhIhLIXW0UNgyKa851BI0SMvbykegBt56H26QVFNwByZGo1riNcJXE5ANs4mvZo8P+/ObkCzJfv3
aEPwn+aPG2gtyJ3umWje5aH2oUMWdTTJbRPOOmK9VnXblvcnupEERqktYUY3YVGyjn3N/CZPn0vV
lwvd1ebRmoqvDaE7JOLTjVCp9qqcHRU4tn4WkxFI123vqXO6vhmQHhJ0u+O2rU+ZE3pJeemlZo3A
S8QF7Ie+BcrmxPnC8htRqI5mw1PS1meI21z1W5fqKrZZS2GMAx/r5wGEX8jpG15vd8eybt0y1Ir7
/rwPVZLWiq4f5b1zI3Eh4SQpiEdxxMRs4cYLh4T+j8sY1R19apUigB18qQmE5woYgUbqi7Gla34W
ANaX4M2gMVzFXX1/pctU3l5WaSxn9uRMAH6KH4Z8Bq2Oh8xeTMq6A9297piTbcegFvos9NF2re1K
TJCAn5eiu1Bj3y9k4TxRMqWbbjBWRTxhaYxeV+kWhx3ZcfHb8uIiHJaYSEn81+6SsByhIBAKNx8k
2pXjpgNIov6ZhDfEKo2d5/+dwCCeZr+TvyzxBmG/eUCLQggxfUDz9oniT7qhq8KhMMgv/z71ZShx
ked6TaK3buTQuwpkgDMkYjECIM9pw7luKYrnRZkLm3eOxoc7r3eCUyqWt6JfTUPzpwvRiqfRzGy9
FnMy/+IRGtFoFfHDeMH0YpQdhLrdjwWrvtZ4lY6Xx+OINhvDuNS9ZWqhyCtbxkfzheRoXAYQveoD
Qa+Kc+Sg3hxkA91GurZt2RuBTYZanLYIlrSG/dwZQH29Sc3bOKT7IDMpJe5RjoGzFa8MWCAt2mpb
IGv5XMvmenJlOG4U/uvr1dscrV9Nuem3rpjAW5cOwcuYMyAUTOEtW3kpT9CeRyk7LFEeTC6JvaGh
D+OVuIhXKy7p6eFOxZnjmD3XMv3DFJpfIprSYGwgqKhOXXPdWEKSEQaNToAY4BN/GgltEUznyz4Y
qtOs8fvc0yiIYXRgaeEIrNkiAB1SmPO4+kaq78lSOQsO/J5SSQTCxcgk5g0l4MW04v5rFvRZAiT+
HL1Pp4nYz2z/caESr5iPTpkgj/R2ozl5KJ3K9y5v0dRueGKhlSifsd+tQaHcKdUmSjjXSMiZH6kN
oubeXxcN7ZuuyUt2PT/AxLC361AjrM+waXbXYAQXHFMfnoInQCe17V240WOyZR82YG4mna6F7SFP
1FHAD9MyQLmlMeqTqiJSctU9PYYPxsfni3nkW6ykKkVhqUMG2dgrgbcFqfW8PW/ECOdTjfivyZJl
l+ZI+ZurehgxHGczx4pGF9oV659Sz6P8Oe+b4QopenuPrdkNI12MVa5kEAGRfd+wOsQbUegG5aRB
IBH1wC4jiTi2sZo9SC1Uly3zfXIrcCRX1I7/FLfMSu31beL/aTYhMn/69r/Vn/2YUwUxWuERajJk
ihc6QRuecRO5KeXHppDYB8oSr5LASoOwp2ZkJ/J3VGe4gxV/VhmP4Hqp8K70z0uctIWFUkL4+Aub
2gq1ztFbIN+w/NUkNwR/K50KJY0X0jNteh/OlyrUV8K3l5vdYa9V4ndnTz00Gf5L6CJTlDSuSkSz
j456vTYeuSb8wPhRbTY2DDiW4r6tCENSOsFJuDpCN5znEB1aboY8JKqJZesMO4UTsRkSK0k5AVHf
Ba9fIAOKyT54hTlwgsxfAdIiaeVMCsmvPQl8VRFC6AifYmqLHOU2vVzh+L3Gxuq2hO0TrRSrBWR1
SS4EK1WfyDuTjqlWPJLWW8eipylcni9MpQAMC+jyKC7Qc2nYNJORQdeRPl8OM2+3kGLa/p22M0iX
gBkv1r/XeROUPd72FhmZddeE2/diEdho3a54WymqtCKzNP6ttVykttn0EVlkzYX+j3mDnn/0sVXt
Ck9xW/sWFCZcztbUO6PsH3n7WlbR91GLGuYeHzlBdWQ2F9xv1mBWaA3UPq3XbhZKpvWlWDPTLTH7
ygNGUbdH4AxZ592wKEPttL1wTFvGNf0/Wi5VMvgcqSc8CMLKXwCQgO2mu7VUKuC/0pfHyCjUHp1T
XHCVZcTjN1MXgei7umGTbJgBhXnWHsIDy7LZ1jHGoHTlac4yv0uiABmbjorpUeHeV5UGQebzcUAm
pe4ml6nA9YGY8DnItSMoZxUXnps0OjUIizMYV0WrGuk6N2lRQhz/CCUpBk0EWLOSEAozy6LH4dcZ
mbo7+3DTc6pgWwypwgWw9vLnQF7HJ4UmO/q80y/U5vgBvBaROLqG6wcHA5H1yi1uCqpMye7/qg/u
yqGpF9KyJxBl8l6+7uTMrRsvFv2KNpzfuY6SiZUNfrQBqOqLAjIfPPSW5K/kbugNO8tlBE4MjSbt
1TNp0VfAOmhB6E4pzo0vSonWeMGj+Udf6B9YRROkkdJennNHwoDuBKBaU2bNfNNGNL3JoRGtpCO4
8i7sIcuRumjqxEQxczpOc71I1PzuPxag/CO8iNx/U2NfVJf+YJF9VeUHIM/akzxZt2jx8VZpbSAY
RXFtdnG6E4KLuVrWY86PnEsSW078Euv9UywHvdV7ScFXgoPmerljnlLwR939xH65uIj7qDZtdyCc
sH6b75Pro0xoPmOrN16NuAmWIOB1BIgsdnLNfarX8rAy66k6JUhgCxfbOshQYFCZlfpbp/s/lMUw
8c+jxKm9TcQeoBH19337gBWDpEPpdZKAfDCY3ApBcrgOVgGPUVcooJFcIfSIajECLYP6myT3w4Qe
a3cGD4NbO4hUyE8fMued8TJf/kh9N40hkd/wBFKjYQsAPqcnAQPlYutoVLJInelHFFlTF0hnJ3iV
WYfBpxQdT+rUbi8llpM+m+q7ovjucMt8QJf5gjG8e4rigT0ng0ZucU5a4Wj3Cf7hxsU97olfC44E
YumUT5RqCsJ1h2up6C2dmNylweZOXjIIoL+Ip/Pcy0LvO6Omr95/WJKHjiIuqffM7UuhKeIDdhNG
ZGBvKTD+wYZJ9LwjRVASD1WVYqI5+KIlMBW8TB1N8FQneEd70IVKjst4Dg57EyQaf/yAfKbRVgFX
0N4l10dU8M7Cb3uYfr0FEpMQ2mJA847oOkC6kdyggO0IUacw+qSelMTwkkDEA0SWBtgh+6TCQaJY
Rv4Fr2+XZ4JhKz/GylzpcerUCU4so1C1ACCwylhvlxkpvsg1XbJArEgknAmvrACk/wIgz5B51Sb4
lKh2ky7ywoHTNIySz4KkpLJhMSQMgAxeiQLmIcIcs9skUOpp6nQi/N1GJvG8a6xF9+abWMRmRjS/
NcC16PjYX9T42HHqmxnOOlSl13DWNELXyYyAfAEBAtMcU8hVLD08Ry0lHCyEm62o7OgZDmovwE3J
qvIE/xcLJydmv/GkXC7FCcabT4QtriH+Tc77Jv3yW57gGpXODRFW8NhrmhgDek+LcFXeQCj5A0nZ
L6ZHuUCJxDQ4XqLii0KYL59pthWgrkvoQnKOuRq3dbXWLtkFLtgJVOlegpNdQZHuMTco50rARSCl
0j/Kwz0QCQSO7ymoiBNFDVt7FZpZ08gDB9EyYJUCUbE+V9R7a+gTryGKkbFyUnUedEDL4KOQW1ar
oBGFZuzMSF+QOWy3EyFA1c4OuvZ3aYRlTruY8oHbKKlEPUyRbI1uc9a/UPaKGcn+/lxbN6bXJaxg
KLx+l90hDq9WtFUzm/l+WMIGdNrbKbN9yl+gj1JujRBKtWvkzk3zOoIMlnvuaNNV5NBuz7Q7cAiz
mngMiOY49gpxcKOJcT1tOzWdAiZO7b0af9dwNpsVH3QXMZU0EvDykie/cwLdaXel0GLhcvrClO5D
s2QCl3oQfYkVY6BAlpqOmkbDGTGpAjc+nOxiKa2R9+MoLb2CZmqC9wkWGSDNp4wkdloegqwtzLpF
BtBoXppu6P35GBSW1GsCzFYYtm19XTDnBeZogs4wvPOOw5nsvnweiG4B2jr31/JRqHbm1Xw8NH5K
XM54gCtv+lO4EsmSPa2ll5L6s23QeLjDBk9Wi6LxQXQZ1lZyAXth6K1Ywe9C0i/gVLqB5RMNEDsa
QZFLER88lafxwns3smXeisGV4cFKQGILj0u2Tl2fDrUqQBlV42eGRERWoVPgvxTVGHXHWrJQQRDc
hPCrDuTTTyWlZaxnCT2Dwb9yWWnRHOXUvpyTEbRRJDf8itF+VO9lMNWtvCmxfWwIBy1rXcSppwlm
pdbfpGLZiJe+wkUF12VKLWF9Q4oLe0cI0SFW7E4DkZfTJet5qRBmjykAmNjlrg5JpHCqx9L+sFRj
vS7asiz13G1BDqT1DKjKwfcPfxGVrd/3/i3SQlJ/CLIPbQfd8ruXfb0woDw1gdyJeILoRYNQh3QG
wHm4mdq9Bzy3Ia9gVi2Gg/gRkncjmCm4qUl2mvE3Kz69KNAEawM7SdePxnVb4r0tOswheUa+AJJi
BZhsd6v7p39v3hbyC5eLzCuVn7nWLNtz4v+jXR3DHy6n4E/24HXY9do6tlhI1MGtYhBNVBTsFFAQ
YGoCJH2Ivp2QHahz4UOvazbSm9j7Jr25j+9EtQ3QDLIQ+Vw403VrMj6945ikOE3A1ueADVCWKNYc
iw2ZKz6S2krqR6AiWsjvwXuDIjWOg75zI7gHyECKWNxRfs3VB6y0smd+ssvMl1b5E5RWN9tleK8m
lvGfBI7E2Zh6B3jVEfIkgQeplZBupGvyNMOKUl7qCnC1MDv2XofHYog1lUijR4ZYSRUH/i/Nc8vV
wroHh1wFsZOGtTxE4eScxV8KDqNiuciK9Y+63Ne0jQtjj0UOcsqcgy9mvGULLSBax1VF8gkjv6U6
ofitfXaVIrfmRhSRHcNOXVucuOrSJRlvquOE/tHr4oGXkjJ6micNXEZRh8rYG99c+cEkzEGc12Lx
PLq5wu34DrG9mixa7p2VYPBkFMH7MewnG52Ff69yLnBH1GLWdbulWVutWq3CjezkRiuEQ3l4jVXo
QS9uI8kjp64k9JF075AhqcMufGd40qXuPW8FFpRGbw9Tk+QvCBwSaNVSO90oRaBM+csURXi9yAnS
4p/8Bxc3djbPH8g5ClAX74ewNwQDMT8obIxgzIOLfdRoVcrb4tu0j0FV2nq1E7NbgLwUqFpMDP6+
T8+hlPOCp0hMuB6GXQQlkomvWOQiCA3UW6GDSgflcZbgW/iidYVeO5VRkW3HLe31+itq2Z/B5mEX
spXUd6c0RSISKrI9Nrcar+7YcUVko4ZA7XKF2lxZNpR/OjUB9308JyXxGYgWmB8EUBJbj09wb0fd
ZB53ZD6t76cqtl9GibVJUwYuklepYWwZHEliRmhEZms1WesBaJ4SBCHEx/xt0Zu+TgeDsxMgTQSq
qVzyGDhi8FVB3SyBDvi7ZizVHrdfnYVEL8FBtg9JmHjqa3QBz01SHfCgEHafK9qSSJBJLmQadNDj
5n2v1w8YcNWb+wLA0MGm+cSo91hu4I86PJ1gPMEXAwv9SmBBJI9O1g/KGqzMfljKSue9ajKXY8Ob
B4WdU3JWLSTWNjoP2zJr8gW/LlxoCOEDZHZ6120qorvP5yVIwFolD9+dhtehJM5CuFI9/rcvz46F
Ojag2WmhXLxDr/0PZzyTCAssFIeFGnHVn2BWmf3vE8ia3nWrOR/TGqwtqgbq+4WJE0Mb8ntDwoT0
k22xF68oxS+6wkts/HyKBBNjNIupOWIsKdDzckT70QA3CN419Zb7OQMxnaFtGRMtP9ner02kpJiS
pHz927toeBmvQhrY96+qwcSn6S3PGsE7a6ONNIyPBCiFxhyq9H+jRVuKAnZEGI0Jqn5ZvuZxUOBH
l+RtileX9y+zI1wSVojKY6Sxk2pV0R8FZg6i3CPKoJpMGnmZeS280GZ3rqtBqfMwZSXfaSyMlusx
zU7gDRzGLOIKAUIzrF6Voi7EMwEuUu9JzersLXpLAUOttyonDUHyRuNRBEWSM5Zc5aE0rrx54fis
Ks2Uc1qXyVjbdWIR9grpgZZdeXZlwNmInlpYNak/eVvtR0eLDrjrOfosZH29li54TPlaVoucZksn
wOOyFf97+8ri3k+AoykTjoOAEPVc6XTX6pDeZ2vyDSLmSdfmLYA27IeBfA5iphCc73unwfGI01Xh
A9YQIRKDlOVVra02Ma/xcQGqKcUyuqsPj89lrYdKI/QnRAmPItQci0q0N9A2KgAcBsAsGWGtnOeP
xneHG1O07+WViqkqNBm6vPmOzbVG6xH11MSJ/OGCaCjr6law406+cx1ouAuXynAFmkWJGSLUWpbn
9VixRepJZR3Y9Ni4UT+x0kYGBIrmw0q89ZvdfYrOeYHBpQ1ojdi6AsLdMNE7nHKCesp/xHTeWr5D
lew6hS4KyXOiWxehLcBm2Pw3H7Rpu4NDAz6icRCq0E51wfNpejLQBvQUqj7bUmZJtaGa64dAabY4
wG1mbiK0rCe1vUzeS5JRev4Mo1Dcfhk1HmRAxFX/JDCjNLbw9dqfohzbfmvbHnSwdIgEFjDvs3Z+
gY5U4HBUZvxPMyjAaeuUK8CQEU0uekhiW7Z0nss0865VU7aFvYyBXBTBvoSnf1lnTnfYGrGWaJLR
ojb8KemxTCGOQvO+eJqBd7dX+f4S3RJAQfe2EpLC5ORvk1pzOsEoTg1CiDXh0lbubOkLblbIjXaa
OQIH952qIq3zr+lLRAaWlYqH5kpjiFiGDZ3oAB3rxSFWTM06gKd+NluTr6Bb4s5YVyTdybjtGg9q
O53iyIds6j/e9ayjKV8gS0XOuzxDdtFnUjAVrA1hJCAMJixK93+H4v0gfG3bm0TMCtagcibTrpbi
dpFfutosE7OoudD0hMCIxQWiM+XfmBWMfRMw5a3Gjt/0QkKHX+BtAi9U9ozE9WXiEE5Ev9ZBJ6+c
tWrVyyiaKwvBLinoCEL8rktgbA4JJyb/ih20zMnlT2H8p4mW6IJcifJ7g44iJoBa5pNhVKti8zCC
QKxossfsHvOUO20aCTub6vGCi8SL6iuZnv6153mQ5gYngM8rH2XfsH/O+WpXkYW0HSQ8bnIJiYQY
ce6jnOdEeiCtkMXgcpBoya8jpnKjf40zu9M2MFVqpYQ2oaQ8rlXyVj8xqrC42mqbdWszlXCVRCb/
c5ZQKr9Tj4nkX270+CT8kRieS7SOjZLK6Hxx+MG2g9Jncf0OdxqNX2Y+79f1qe/vQuGUU4p+TJzh
JMu8uBzVQLqIo9qlA4AU2Zp2hm4n5zznyKRbN5S9MgMsDvP5Agu/aG3B3T7/uq2fA9wQJErUgFet
Iogye5DLaSq62t6ZtrOPhcPtiWGKcp0WnTIdh/4vzI1yTiho1THzx4WRaA/LJJq+mzF3u+jYofyq
g+DGHzexsqw7UKv3bkoQU5Cn0b1sG1qIV9Q1gsk0st2e1IMooIpb34mvrnLLsig1wp0Iujn4ULfn
oj6UzjuYvKPwKh/EFPOzYqAqWQiUpxbbWISLAwAm1vKe9U4Iz8HG5H6Wknd0Fvcl1B1iIB8BRe/B
tbGUA/d0AdvPEwZiAHaNcMmNZz5hz4EcvWA6WvFOPpNgGwAGAAJmqItLXpCZnoZXCIpOWXynI1oP
b6NdfO3xim3Ilccg3XS9IEmwi0Q9Gat5ohIL+pgdc8hjzAxMXvW4I+Y9Isv7tyhqt6SjdLQAqiZn
z3fpV7Q38A425CMNfi0QbZdbL/to7BEx6sgAZN6LN8nDfZVwuV1kZM5pId3CsoDfTxXSxZys9qOj
hwdf+7sLy0XaOnkDmDViPSlSpbOar11lv7ekgzpm+Imk5Uo1L8Lwyk9FDWW7CQ3qB+9LwDcZNSvX
4WTGEYaymXFcXUJP3pB2fATl8vUm4sd/A5v2UvTNe6aAqfo4S4OGyM8SPlb15QQsXm1ZQCNK1OEd
R8zyyD0iKD+GEUbiQ7vGDHhHRFrN/ybxh5hpEt69Qk6GccHrto9Nq85PrlrWoV3xyj9Ga3IhKAjO
Rn+U2+9Jw3RSdefUfm/0mUwoB452e2X7RISkPk0WCjhqs30h8BLZf45bEGxvPohPYXGSd6uScUMj
ZW47uvyKUfiEomKpPruvbZ+ZeMgIEcLrqTWhgtW+yaE0KBHOY1bcBQcnQasMwx1vVgThrIK/SMmh
NPHHnTVU9W0bgMxw1b5npT0S22J8gcXTgT32yyCb/joB/gT65YiPhS6Er9P5p/Pv4VGVe7VhPMQP
PYK8cdM/17MKq2XDLIvMpEUcv82dclUcKeUMMamzSGSr9zUhmhSWVFqPGZKpialyGqNtcezl5/7m
JA8tZwSddqzTkLNp4iffgzyKu6Ge+gd028/ERpNq/7gqdtws/f2MglrxvdUP3Jvzo/YgoPCJNqv8
jTXZ7BkEoQcu9aX2ljGxzMkwiTw/wAMNHzhgqiSs+qgChMMCTdNhDce8bCHSafaAhlEdt79HK8Gf
PF5sN2WO5NfeQc3gRn/JxJloG9BWPsjJkYNpWEFGmoLkc7PUGtP3RIA8c4S4oInqAyWj7KThz9XX
FZ3suWxL4AwC+p0auhVNNzv2kPtH8PmqA06Ls98rqC9Kr6iYeOG3hjtZ8ZNpLRisvW+6FpHLQ6hp
B0in6wKh3FPEXmVToo7/w4V8ELiizjFgkfy4fOSFSPSTnODu6ni7kcRHDXDXakp0GLJhA+jso09k
5+Uwmjh9i9W9CUHrML+rDXE5/yKJl9yndcBQb7HrSBcqpN7oJstqKB3Mvs8IQmof62GXUnllTXOc
iiV8t0hgOubdzkdjqNvF4NEq2mvhpqd55NG5N6JBZqzXWuzaWcE0r0FN1fseUxfdYqYA9+Xc/AqF
6OjfSl9VtgBfF3SLir0LgPHnn6CA2sE5hBSdgzMIDArz0TPgT0wBrC1qhsTbBHe+MzyiciRwZqlS
0djolhUoe5veIFsafTxXQWz8BxU0+JNdz/OOlHrQUjOhz9OutOmY9h45R6uc81W5OBs9MuGmwYZ3
PDtxXGoHouX3cBqEya3DEHCOjGTsrjLa9dfXD3G3Uu/12aVHORCIekf7RGxfAqCuu+I5aT9/u1q6
Dfx0XnTXZIxX4pPG28CtsCf//ED4w1v/RpKHRO+cNQ6we2hBbVb7tbeuzgJZ5BHt3UW0frWeX/DL
mDkvKsUzR9EbxtO7dqrpQlzrN7g8aSbF3DqthMHOs6Dgcr0MdiaxerWT/+tJh5hPgEUMva4hXDal
7ip37O/4kVAADeKZNH62Nn5xhM25taVfjDxXQs1u9RnXFiKGt8yEcaalf846XlpFBAP4xrD8BGmn
TGjWYv/tgQWfXB6uzKT3adbE91Wmb5ZST2DQKjtxn1X0CF0XvTcUvhSgApcFAH1dRz7HXIw6UCKs
ZoKxhl3xdhE9Cyvi80/IT7qeWbQE8J/gGffr/eSEsutOsZjGO4lsa4+Cg1gA6JeonaWfj/PVRyYp
dbbnFB/Xmw6L5B3IjZxfbWMLYti5vRHnR1DQ5dnXbsPdTesFE98tyQ51GZ77GO3Z9W4tFgBa5/7e
kkNAlJu/EPchr36XCzcn9FZCZkMSbRKMdgdMJBy5m6L/ZGnIyAwh4T26t/nbTaPe15G4Ldq9N0S2
9wDI5WsQU6vM88YBBP75eTx88x3fFY4gvWMnwWgo6XD461X6OmEXzXAodYqZpKwak/w/uOjPBg9q
wx5XxClfBySsYl1O8l/iH7gFTXlqTYDN5nHUvN+hdFndYduijpR6eYXqQPvFiLhd/NZI1Jo/ZFRU
AVDxxHdL8toYKv74Jtg4Y21TSpqaCw1MxAuZeDbw2L+9bBSaSamzMxz/dcsi403xzmfrA0POw+mm
Ocq3BIjtTzDsFQ4W+BiF5eAPvWVowGChtaehBZvJu4j4Qzaro5itLnnT8FHkjgm9OsN9dTZiv87f
AuDk/YpkC0wAXZ7NKGvQmoUnB38KtFF7bRfZ54Vyegi9s3ZQQLMmXmMHIP4nfh8y8Qufmpvun0g7
ysJXDjQorgx4QVZHssQfP8rD5KOndwd5PJpqLYKvLlgPHUudXu4sZYVQcfCRI5ePB2HEdlCLUb9L
NeR6qMeYJsy+b/CBPEuQKUQlFfM8gHO/PLQYpLWgiqrmisjkwnPOx1AaQCqZrEzP4YHEqXc+yJ/Z
v62dczqREODxXFQ+0OHj4zbOr3T2lL5NhtMuFtK3WVQr0E24KDHAxkalIoaphSm7gag+8aOaHrMP
/rYw/Hj9A+CeWMb7wbwLcvqS10F7cfvTx6snm/pfswYRpFFdNdXj1/QUoTC9d5wTGdC4saZbrhUg
h98zAQRYEd5jk5HCZ/oEbTJoNF7Z4zTLdZkqt2glh1us04dS2003PSiYonRmOT2VW21xIyoks5Db
1L5gC8/g5Gb075vp
`protect end_protected
