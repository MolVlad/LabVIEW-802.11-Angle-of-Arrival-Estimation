`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
M+mra5JQ2D3ac0itHRwGS5+PlH2+FajJaLG0gxKhiJp3nrc0xkm25HnDCVrL0ixHh7vW2LJ3bEOC
yZDe9E6BQw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TXzc5w6/FdVxkIqkwy8EoUYisyWwhVYxPD4KhhtWY0Y5wK0dQvbQ+0xJj1AnQnaCHWMtsC9eeAtU
Y5YTGOUKazeqeikhJrDq/ozoFuRcvu3GO8VmDO8kbu2faI8fKGJqAc5txqDS6J9aOWy/cYRRounZ
ubldhP94KzuOW3dfMik=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o9l9rdGQrh0ABfcImQKMcOiLTT6u2PbjeroAzHkGIR2z398S3xAgzz6o8OpGXtBbPXKMOFl4DNdp
K0a6ZQiNYcHiA+DGHKVbicwg18akcYYdxJmiJFQkC4JE9y7brBdWUFSsSLcuY7pzPhOjQ0yM4TfB
8P4WWg06ZwWkN5vwFByIzW56Et+Izk8eEtZZGEzNG/3jX4MU9gz/uvSQzJM23Y6+H+2eUjjN8ktb
f7Lmy/D7tKZszfPr8H25Qr9L8sp1hlA0ICRhs0Lo/oAWOdYakXAdESC3wF6mgWavInI4leQ5ngJM
0zJ+5N/+iGb8+IGqqmH7/nZy2wSelqWCM4beVw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h2AqkNF6D5bgCl38SMNMPg+xqIaOoG53K9bw9Vux8PwnKdr0iN0y+DK4e0ptxfnCmn8mHSpIxYQg
cLEGTw130SVUqE5gASCJufIo8peSjb7aECZsLD65pqTofc+5V+PyJb18j1515iE2EhHc4YHqndEP
3LCrdE1xQ4Bta78g0vfwTys/dxOJiYw9Ta00XDOc+wh90zq1bDm74nWvMEjHihbXgUD/Kih2SCYg
aYVNKdGYDWjFQrRCO1lWRW187f1Ft7sX+O266tWzZCBQ53RG4S/E4+u9Acuol7yQhYHsTOyXv/DE
mbFmRnjn5hUXDNrOs4QhU+K/Q8kDURbjx+C67g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E8ZK41ejIg+6X7saBqjTv2+1NTnF7a62Yx2D/D3vkubIHRan92O0WUQeH7BmT4iOHSAu+Y1JXHDq
dFSI1VSDhKn3SiSyiIkkKYiJ7YYkbwG0fpz3ict4jTdri/mPUV5vTZMPjpAXfnTuV3Fi6d1rBAVa
b6oDEKPZCX7odh1X2z/eHWEhj3c0er2nRzIdIMDIfs41nHPqgefp8vTWCFyUUsv1zlI/srO1nOSk
uKydwNfubbcpFrjNBHD188DlPp/HfzfwD7OBeKigFQ8EuUm5M4m+Dvs2zFXOyttJGjyQl8MNBpKt
9Frw+BvTh5uySzFXX0GqGlsNMw0BkvVPgq87Ag==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kRfis3qig7VYzP52YVL2CDqOSImORBNxm0ARwN1VGEHqA7XlO+GEfBAW5piyoTiFQ0M/LCOS8uzo
iBrTsG4kk0mK9cqVe8dup1DeqnbcHVrbmZzojlp1L6ok54qUThXnEi7DGMCgwgje6XUx412gxj9h
c7h7/BQ7yh67Rptq5CE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DAj6RDIXHwEpVjBtlBHOojV/j1VEISzSruAf88+O+qyY+YZSygTfA+rDLtNqP7khBX6gY48wH6qk
QQWp7TXJuDSkJFKaoPJOK+TvhaSz7pnQL8E4cuyHQRGBnDu6un9Mi35xv77En06Guz1LHztj5ZJd
gSrHd9wyIYK0fkF7+0l5L8CZ8PapvXf5+QivB+wQIlvSL3MgOTEkkrI8ALnP4CPATe+QPpttgoma
Q3isjALfKhQ6Mbz0ejzdCJuAJspO8HQ8JnosieJJkLPg3PC1hCkWlTrME2TUwUrls6oN7Td1nWzh
8m4Z+beIMbumQvfihjQZNVV1XWHl5tphd226aw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71392)
`protect data_block
7OUZ2OXBmoBmScF0z9HQAmALS71cR9wrZwI7AR5Fm+euzp8/3fXla6Jjk8BOh6meimhTg1Y+A6UO
pdy2wL4cVg+M1Yqppx0sOhr24QgSmDHaNtWCwwU2ndHwq//7aDY55ibFDkMfIU2AzX2DXzG28S3x
8BdsAUdy/ZDicCm75YvsRfn7a3JhkSVYq9D9fkoFd0RSvvpzIE2Gu2eGZm1hT8wGQo+/Y8TKqiLS
03E0ijDF9eiKXDd3sFzbaybqGKh0rTvu69W46+qKnAmfbaoxZIkD/J+P5qDMXmrzh3QDVMFdtLSK
w8URILQb+Arso/xsrOi/UZCNheH2bqpXe0qwFWSOyx5j2k67IIdIp8e8Kpq/7NwhoTFPykKUMJAh
Dohm39UjKuuwYVsHHVenlEWhLspQL4Ae/NWP2d8dP2Q+f7OGLXVTkQISbxYHo0F4fxPJh6sQsEOR
4kmV+VqFN8BmZWfhTKDaUMVxJINcT599rTqkunm5EmVBY4wANajDIyOxhqkQopH2gdZ5DY2eBY2K
7ae6i6fRBkjAy8H8VJl2QBQVNR6aFI72uAHwip7DGNlNR7gouftMKKEi3ZSg4t/LN8/jFA7bwCXL
wV+X+xtzxDlKKqQ61oH8zcbbaQ9T40DLtNHHxsLnOkPSJGDx3jT47271BT11hHSUx1lSr5elCnCs
vXETuhMulOeL3UiDUwalpLHfe58YH8gnNv9tZchXlPD9bcyiqHk5sfjLJXhhWXnZPJukCyt7ekYa
SIyTh3pnnhpsINKX8VzQdMUjXtF3+jzHXWhRu2CcJts/m2Tg97UgimSbQCOxlaIq7XXNBI1kdCkG
oKBdV3Gb3Zhwq82ezsdmCyqhdy4SgnaDr5ytKtUMkl2obJal8oATamj29B+XLpstcs+dyFbbAc8F
qg3BskeVuTCj1mv6LGBLjODx5dQVB5mGQBVlkjPwiBSkWhJ0EHqNMi90zLFitfOtj54qoQcm2HsT
j36JkfZ5rqhAuZNHUqlHucIPca264reeu61FsdypOA3kFEV+jHZ2j0CfxXYmwBZK2dxw+2kuxY2w
FpzW+z/qVntGnHeeaZ2FPrU1WZIx5wsybY+ZoTQJyEgXBU+yb2tZ3lUCd0F833KAc7l9le24gmIS
ljehbXVn9ZxTXDnDQA9HLjM+3dwgvFUih6ud9KFpijlPBNO+rqFZV43xIwFnUTpSnN2jjQYWav1c
902mkuoxEXUTg4fB8DMpvC2dkKgOg9C8Qr2JEs+3ttRLTSEZz7Zt2KY5hHQnec4YOndVgvK8Dmy/
RQep0b1hfWDqU2w1pzzT3yUah/8fv7onEItLXFMoyyz5zYVlwm//GMDRir4ZNVrVjLS4nbTIff+u
ooiNtpukOtvqKIrdvkXpiNAsDUwYm0mxcUGXI9hO323CIkFFpIoBrUEQ8H+L7s+TE7GsbhO4AqCS
/8/4jlauFVjozge6hzCgybLrOslcKbzlppAvHsKVDAdSe6AVkfZA94Vjt5NPoeK0iQVBS96gOviS
HwIh+IlNYHe5w7HzuvwZPTa1+ggQlf6HMXq+LZZCkF5/q+xjgyLNMMh2Dr4p669ubCrXTxBn0oFy
j7fW07hMh2M7z2Eh7QQLlTaywUQaiEo+nFGLI5NDg8WNpY6xv45sG4jvdJ6ZPk/HM/v2JnihSS8a
3Y5D+NE4nMgmcN7pdF8BvaJcj1cwpNd+9cnBvzrxM+8HKPae3ga8j3bT/+o8JkZVJJ1caBl/uosv
kijEpGqwGulDsn8iJW1nC8FcY6Qzvj/kkuDXxv5XM6d1EE2VpVxKNiSq3m3ZmbyrSl3KxaYn90xq
/16BK8StYtZKf7v6ZdFK+Wha5pBhFFCz/8Cplpx9lsaXp2DJ0iY000//qtLn02aSdHZITx6EI8+N
w+2JlSUPM26Zo/ZxQM3i7Wgfvy5wgMQPW23wev05A19GWKAupQdnVXNgKgJyUdKuKaUDquhyTqOG
kkjAnsXeAz2MoT5hFYEtfCuDyMqP8S4LVuPCZ00oTIEN24lCc89ooS7CyUE3HZoq1dvvevKgQu6U
/xZe1C4KRufl3z1eRgVbysDsLW8FvHVMWWWyxvAKRGQj18BQmrYGlkVcIl9os2roIJB39K58dbvC
hmwnVPEKX5xnOifBz47ValG5vLuoxWlNkusexR0MS1EwO2AjZ8XRnS9bFeIFkCoWw6o+nvIHEQJd
AcC+Ajn5RX79gBn+d9x5Ic+7Wyh8dbTIELjlPA7J/zelQWm2m7i1cDWaxg4j0O301c8UXRDivbQU
so6TsXzgbapXUcR/ANOk1FdPnmVTVbYZdhE1zZ1REumzICLUCv0gqnkzl+6PGlDD65F/QXsVmvbq
njQe2WpBBW7B/23ABVVJdan6uIVACfBQUp1+UsDKe1LJQnFTuC6W87uNLHkUSsqj4MRZnjEW8asK
iQVOe1B1UfNbu6yZsFHvy2I5MvEU74ChHAnXHMsKVc1YB0t6gFLG6nlQGEpoMPYV9eEuMeaCSWE7
r4zzrZr0JF+t1owqwhHqrytWQreoSJrcXDc4HGtuB45gXntxitkNcEyEDF2r2T6TtZd+ES0RpQPk
vYR11A903rZdXg0Cl4jw1OvoaZ2V52WDtWmLcuUaR9uiZKe+yBcnz1zEcEdElYcbV4qeaD9LTk7M
LRQVJbHlBwSRbhg9Gli2oBx+F1VWb3XJDFZ0OWR6ioabvGRdJqarFcZoQFwtCpQuJ8kqfUonMEd7
9ElVm+QBXEsuOkGYYj53udpBEZhprTCvIhGDydB+fZ6Y/xSRk3zaeAFiB+dKndpvjdwl+w30J4UT
UhrYHFf7us0DuGayq4/lSgHcH1bRoYo1iBkTyKUf7ssgOaLgajo1b34QtYBm3DRaEdf/cKVR8A7g
aLBWJfEcee+ue9G0g/nhUZZVrOsRFh9k0Z5fAfys7krEW/VXhA0njSqUY0XPtjHkeyTktMWpYJ+J
1n55z0K44u/w2GBJ39M49vANYYwK1h1WDyG54fSKxXGMAzQW3NGjuv9T2DbrRKatoWNbaMtdSnjR
sPzmjg0kH/9ezFLR5e1WmSjBgu9cDb4mRCwSl2cErcOLg6/eHGU/m5+0PJrf5j/JNXKTAKyaW5vP
yb5mE+5DETriJGXfiV9fUlnojIuIzGAKTqrrfU417MCccHyRYmHLTPNG+lQTqy5zEBjgKLW5Kp7H
zA6/wkOWetfi49FVZE+iDEfrQxJl/ZFg/HL72Ivc/geZcPuqHgymA+y+C0f+NLXdkvAOhwzAX7dc
yLTrNMeoveCoij47PxAL1aqHFwaV/sxqs7FNVrlqDBrq7gXn75AGiKcdtAwkAGeUjxKP3mmncuK5
zlI6AQOCvNoUGFFJn1wyA7K2gBwDv/ZEid3nRMkSNwS87yoJR4/+/rf+huB5MTw1DIsls6jFwv9r
hW11uJpxzsJHLTTjAO83UhRLjzH8RyXkFDkp6TZ0vlPNVWWw4JaQuSQOrgUidOVwrAQDQc21JAbS
tg72v4X33YDDRm4MVQelueQAz6WekrUXJS4yVDToSVS/j9S31Y2saZEunNfK5+J2u/Jd10stb7Fi
V2lfVvD0+qEKMzm2PGhuDPugltLoxNEbjIBWAFxdVbTmUgAMd9xZTzU9dqTHPYoNJMIa2TPA7qxX
B0ebJ3+csvi7myoHUoEaK+HWf57+6MBwz9or4955mvsLTju0zJqB5V0L0LOj5S+aIdBNLS9wrDpt
dsYqEIT2ATM4G5+4Z1QimdOf5vzdXe45iJ6q/uVKUUQkh9Mtx0MBcqpxtLk0DrgkxYYbkWtTjXlo
adD4dJuMjAU/mi9OhsORFyoltlcHfg4vZW3/mywTs2KxcdGNMCzNrauQWaOeZdHWWLuxn3gJbjlc
i+Z6vLDOXbNy9urlHW8MJG/w2QNihyDIDXMq+1Anir0VuRvOYAl9UJUQmeVslNYjINawMuu3zxXc
RPhlatunFdIU6mOsZaqFtZMLQo0PncZ9uez3z2kmPwlelNRkVcQChV0TKLw7HfmGpr9nxIWq7ox1
NnH6b8IeXhlMWAWiWuIR0voWZg3j1W+jiVqZfRans+jbodgz8+TMS/QC6q/MQduBDBNcTvJF25fr
5WPZh4A+XTCtThYhHL/TwV3YnZMf6q/GdLTsHKXqrQ7nu5XINPe0I8qdh8SKkgyhxMYArIQbHf80
JHl8OzltH8+EP8EhPlwF9OHsumF8Cl+4OeAYDD9PeXzBsV7lYsCCB2oXIzIMrGMjEEUrcRMhv4DI
hIVKffFPyd1O2pQ08wtY9Ow2xnyyhTPj7wmGKEcE6saFbnbZNdEVu+4CpFV4WJuBW2lONnAWVIbl
dGfcEf8OkV5VVxMOO7UJefGhCFT7JtBqd769NJePUdFC2IHi9A+A+cyEuh5U8TJ2p9cWlLyeOKQK
VhJ7wE9GnHowd5pLRw7EunxqRJ7kyhWmBR56or4g4cWeNIj7cL+QqnbZ4KEXskvf/LsUJNM96/jq
tYgw3tAV5y2EmxA3FPATVzuSkX8jlyj/37oCZd827VnyiR9mprKDQURnyt+FEYuHJVx4PyDxvYVK
1QWKYwmbuk0m0/SRtktfb3ZgIZ417Pez521Wf7xopn9fRPd99GG2jHfiObs9RByAutQKTREJuEip
27rAPqaRq0396pq6IBAzw/a7rcYEX8Vav9kLLBzz7iL817LeIzjrhlRGluEmKmLRElf7hQMDLi+M
+Q3kXifIw0m86lGCYE3br11NaleF405Fz2WNFC0A33AKjGE1LD2qmekOVvSWkfuCKyxqRLgBScNw
BZtA96q2wNkTbDFPGS3l33Z0SoCp8YS7H/5riFORUeOmdPwb6plZQ1iwMw7uHWBzw4eTDY26XjOd
vdKZhignc7hnDxBq95od8vprXhPiVHn/v0y+M8EbZL2Z7jAKIMutT24LPED8s1tFu/gcbKjEWovJ
Ft1cyR41d5S9MTVgTFifwSMAeddzCQY3uP4RijxMRgQx5PJGTtPbGr17gdqIUIxGwyD5jZKX4m7f
fjH+NdDARbpI8CELmCH51FVaeq12NxXop6prMBlauMiilqcMfZrx40mDvbBIiuH8uBfien7YcXlo
pNNjyepljQYGOGrpYW6KxYru7eCJjf3ozoRAKsV0VoNk+cHUtWP7rSHn86whQxCvG1X/rFnoQ4VV
T9xaXsYP9Bojm/u4ZIpwgDk4QyDhopXvQIXcQDwtawIp5HLqtdKWOHhBPPSO4+nYL0azCARUe9oR
AhGe/kZJvgT8dC+Lmr2+NUu6PO3yZLrz4wDV4UZtSa1uY15XcXaiAohFQEUgGBYhovd9MpAENO+u
S7Or++ZEVoT66zjmdlWEhkFzQgEUxYxz6ovrCuvxXo+VCAOrgi2/LsuIhLjkUkBzfcY97x8LwA3c
IA7Sy6LfKyUcSHhMv2EV4EQrcQ40TfW/O4VVolpB2kG6C3l4MQH5fWQ/eYHJF1XW/eDgC0pnbd7Q
WJDO5taGHkUUm9FjUCGIilyTa6oKsqnaJOvYOfYKHwAQ8gocAgMcaa8Rei7brW/Z5BwxmXzth/1y
Mm1jKyNFn/48czLUyDvz7wnGNFlFdYh9j3CTCecpyaQ1JnJZ93RMF131VXoXOUIgFD1QTLOB4ugY
tk1+jOAmx4FzzdcMY8J+HJhFX8MPf8Sj10pGYO1SyLEfgqsIwxPnrCLQ19C7I/gNV4uIFJFKQzNA
jJhPhm/3SUtv1pP/RA8WSPD6ZErd0OXz96jW5hse0QWovVJLLu/SEpb9V8juXNKEHbrcTuiCfmaj
j3DSQH8x97oY6bU/CImjQFNONKWjEPNoH1zaelRXF+Cbdvf36iGgfJDEJNWwEkQgWjlxonz7rWVT
nNceBp+wp4Rajy7fUJjmUt7xMzTp2tiIjwjb5Rrd30X/GuUDMW0twrTqS9YlYJMYjHt19h5+Qcsp
ebCDDcpElsA37QdOmEzagDHPI+qHXOPLRluuU+D/W7l0dP+MxXvKfIFGogF7aS18pGt3utRgFUxd
PGh0IwxWaxXiEtOd5Hr/eO6hlCNIPWwKEdrxK1NVeEC6jahzonWWNyjuU3zCKyJD9Gz7abjdDDVg
eUec6NTSBC9eJJ/46FsDR0Ezru6ssxsCquyk2tzVqcNH15kMkLPtl5a4SPoE7Nhx5o70B9MouOaB
v2SDYXN9j/1X9liWKMoTMaWg5aARujnTgHGMR4e2G5mX80VRg6h5N79zqs9m+q+XUuPagH5M3sHP
rR4jIiQ4DkHUHOmlSxVhpy7k4lirLEI79X6+qVITadd0Iz+fVEJ6Z8bH2D+uxyqk5cQfldsVpcRe
lvOXS36xcI0wfzvjlR0e1sMu5HKo3PBiOqDFE94tmxquMytgBu0JW/8vcygICxoGF+dukuI/rLQP
jV1Q3WbRvVjz55cG7FGDBOJ78nKWh5frJ1NI9nmYoFEdpC3qsPfbWnGpeXts4MvlUwSi5vVpvRRB
5sbpCqf5DqXv/KliyTAP+Z7x3+BAFUAhBKKolQnv/XsbR+f0DL8NEj7MqHFDK5w8Ovlu+2bkm2P9
OmjICkPMCD3AHGBUJVbnmgbbnveu7BF+LJMGoRCtdVTP/uarbLOtmAkl960sAl+fVz4QhYbV2ewi
G7aeHrtBq36I4yGIlDQWTNaoE+cWrLdCL+M80C4LMBsZTgnRTyjXr1MtPHDcOuYJYgD6O7gVcgFa
ZkEK7ZNTgBlQCYNlsAi1oirUeRj6pPjXZ1vz37p6gXadP0e7p6wngEEtFjTdzxkcYpxcYMPhOYho
PwmrcFko/VrPnADb5vZKfsabe7o4waqEuNYnz3nOr2DvaBNGqUVu7btGWtr6/y56XTkbBdMYwLuS
05HICvq3kl46MtW28gz8fHT1v7IwCefBLLVSlgdkkKLXfwA6qzaZrXoumKowiXIpki/N0nRRJna1
EkhEd0T608Zp5B/dTQmXAl37tdAUCzDjZ01AwiIBSa2lPz32asKW9p9ndlu3dSB4dEAW5JJbL8bJ
VF0cUA1BwoWZtpg+nHkiBqbWsPSYbAPrxBkqNz/nvYIf65DE60ko4MpMugE4zXoh81CvbsamDJKH
B02hs3pw5ymdbFvISCjTQMqYgyQxOT804t/UXS+xRK1kpUu5olnmMR+7Tj0N4P3Gq0Q947QWBxQb
Rhy7/ZRi4e8AayKvRGhaSAZkYHWFWGogGf6+SxPhSfWnB4o9mQsI5P0P2qfJoKDuNYavJjFgFinq
oKjQCpoB+b7jchUQ3+y3g4Wvj6SvcxKeotri0ith4rf1m5udACKgr5VbU+VrpNzZU44d7ANq/ub/
N3agGGnSNRQXHD+9Crw09z1E3CRuxW6fgWjb8VE0SsHF+HwqV4/5l6dQNcMlQw4llK/s9v8YoUVr
wwyrLBZC5cjiUEIQRD7GVKmOfp8J8L6EQrUdkYPpCEpzBMZPlY3uMw/JMnE8vyuLAJbaqE1rYDdQ
mfAKLGwiqzdS1rsO91Ay1uosPJYSYgL92+dTAMkvSFoeAPbwiP0fBFfzQQi/ihkfVn8KYYSviEYQ
4YdduKQn03100TYsq39hMzmf45WJTPZf6v5uWWt1jRopa+AbEN2JovM/7HcaQCZx7apnCpFoXVpd
wIpHu/2GUNHNu/Rp2Yb8hO3QhtirNVvIEfheAhusvsTaZjkJE6Sx8Idpf/kyDtzE5deq0qxhT7u7
3uIpN7PE+O0glZG6lBFdI0pB18yp4r7JBJxU1zQNOd7Pr0soGYkg539TqANH9lWc4O2fnbqOvimh
nYvlyLPfJG4q8Be2Bty2n1xIgI3euFfIeTTgCH7i+7WgoRVoDLC3DhiabTfC4PMABlJEoefTYvam
Z9yYLLlVl4YORCxsCebCiwIjE3Nax1AT7IxHzPm6OJGbWNM38w7QHcw2vWVc/9B6R9WRoDpo2jgu
GJhleabJPRrkPasNd22y0Mzxa1T2noiKHEJP+oiSS3+AdNJQkte63iw3a0bb8dtrZwRLU2Yv1O9P
LAnjYgFu4YivspkBZ1fM0r4nGocSRnvz0ApG1FXS1Qh1opDrsaaDOf51W973qzljmEm9quGPzhz1
4ArcrlWHs/EGFxADVE4GVaHHxr56xqprVATgxchvljfFllNVwoVJ3z8s6vsck6i2lA5dyqkP4+cu
GcYiwIVQb/rvbmbgBpMKHGS61AJ7Ib6KsIjT+h1WOJ2edzaAKS87tpi1/kKz3F9Ie0M2C7edT6bl
5Ts4jvI2pJQkSHUJizjmn9DAoN93/bmb+5G4Om053qSAodyZdrrZEncXawm7COFVL7Rgg8F17ctp
1pe2OEF0793a8LzST6j23B8NsTzjZfTsj/0RNT1L8OYTo219FgbFUYNh8k/7wXe/weNcI3Iwm0GH
TyhudV31DEWgZWRvYVrsNmyDJDY5ZZgw8DdvNnrFFUy7Amji7uuEVcWwGT8kgU/DFH7lEkEitR3U
eluG3x2rf80EMAGh891Xc7WEZ/6p2vnzirRajv5FoUzgBNH7JPFKnRCQU7y1a3us86NY0uRiMjYQ
1lEa6do6wYnud5paZ7wtQ6JU0IFtzi3x2I4z0HX/I+uNpXdC4aak/nYRjNKZNvESF/CWVU4Q9oyr
niVsRfD6ucyF/IU/M3EuFgW7+nGLlNI8VuiKGbf/urTM+HVHtVfw3SFl+rdiktaa+UhJ7WBx3XGi
E0IFnz4HumvUOlwz2kTy03lnIhFG6rd0nJbXxd3miVfmI2uoKawBqv7c37D0P2GFlozSJfu5R5MU
HqIB+Qw4fpMK1yQgBO8Izb+V+xi7mh5mSsEQ38XaJ/XeDK51kN9IfVca5I7JAbH8n8crS28j6tuB
H73Ye+Noxi7+skEOhKVfLJFNtWLljFKBDR6N14lbX7EqrHoieN60AhY3Q9b5juvxSC6kz4UTW0SB
8iZMVC9GYWKKvruwTh2Ci1Z2VPr63R6dF4D7wqyXSlBpi1CeixAzwgbbxE8wJNEWBAhOhPyO1AM4
Sxe1B10lZARZeRCPvVWq4FNZ9yVQN+g9nwpA0P8LBypp4CPff0ugiiWeGIs0KN1I7mFxQTaX+52y
Jss8Ha28zLPOlvKK4xPwL0DzTL6ToiMAn12gCXQBdtIxhZ/vLflOsoyvGT0J3hCH8v3exjz4Mfp2
TgHpDrPfLpAGRVz5La4zEHg7fQEUdSTcHCB9+yo9VyhLDM/12t819o+EkSzDh+Fox1Udw+wcEzw4
tvsA9n1Aab1mNgZDvPrOqzBRXFP/bJmMWzD/YPzTj0xXghMdQFc7qN3+W281KtHkD9N+nVCwHRfI
5n8Jx21Zod5nAQ0EnPwzz75Qk7IiHYxokA3PX91cNYRAN9SG1sU0gtpnXkeXjXROXWghdqhkTr8h
SPptUqIHBCI9P7k2f9fUuhcZ3xzpEq0FPZkDbsDRJVhdvM2/xL15z4Kg2mumR0i38SR0Z3CbOgxS
FSHOfYhGItDrzso4evqzrni0WgZNIQqJOPLadk/weG56vb90Bg3CP1gF35Lw9Fn+zWdFr7ergfap
CCFumIJ3/XCeOhq/J/Q+Xy5nt/oUvqTi10pt3lzAPScr5KEdQ/naBtMGBJDvi0Ro3xvaMpE/iD1l
w2z6wH2XJN0HFQF9LgMUa7r4/zttciSh5twEfirQjI+UY1VwF5mxiJO5ZZKG3OG5YIAhXBTuWVMi
wWzOJLwgSw/xvwsZcVfj+j704RENw+mK672EFVeFvifESrtXwh7+TVsRuopAnOxaK4rtPxi2QEQh
hj/6+WtArjd9Q8HcfWaunQIX650Oa2LgQ6kGzHEveauXdNu4eZxcAUbZQbm1pxuyNLgXattksdea
9N6SUnxXzLS9qFcdUby9bg8LvnMDb8erxBT7d7MXZzNKaa+xeOpyE4Gk4LWekzljnMPkbfG0gIqC
ymvBT0IBmY/k+mkd+AM6WdfnjhicVXivIbK/BO493Dl1ymdbLRmEvaVVedCApWDWxcl0v3c6SwrF
4bXVqaMpFaQFh9g7RufzULbQZFKvxd07PshAJmzvHYNkEfZvJwfyMXdNSblaimQlljW5bFNPfBr9
PfTYgO6Np+c5QIw19KVOkfwdYw6fhy/F2UWiGfFpguwROptCFkKhwptF4jKuSEK9x+QtAXCfBmSv
htENbgAe5lD6i/A/J63p8rFuMK1XVUD7vx5WgG2rUovZF8dehWtLYPwu4jgAuV92XEbXR5CKlBOL
PJYR7CUBfCH5urfest6QtFninRnNwalxB+0q1o7hKwBvNGlTYi+p+lIde3geZCyxTbXfYVkvGn3d
yc3CV9KWiwaOTJ7ptsw884dogGXWUNkfbIDxuDpN6zrcld9U9k+p3Z3qo5eGabVUn4tg7KMPOij4
1dKbbKyNfnZ+vENfREy+8g1Jd/qufTIY8+7f/F2z8y9sZgu5rpRClUh5JD9WyDsigoFcEqImbX0u
1Rme2Rm5zhrxKKIO/pWw+bFYpt+kSnhaDdjM531AJUiJtrR2WxEp04E+LfOLJ4O9RTdglIkoNeL5
thGLp2JDr2sUnd4nt/yBLEdm641KVXACMEZdGwotfUwvdKy1/nFD5+iMAeCcQymn36edCZEPhP+K
9FShQCdvPUgJoWCDPNUtk2f5C7FlM3uEwcqBs5VHTdS729/yVSbFYcljSV0zncgy5OdXnjnX8wl6
Q8K5vlQKTtKziHXqeseBfH7zXcm4BHqBBEiJxJIbNQzvK3Q7ZmZCciP/L0ZneCISe5CScPkJtYie
anzLgzUUlxD9903M8nXNVdVQ+SRrd4Hv+fuShW5BO+XdSWCvnVs+gA9uGxU3pPuAbKaLty83Qurh
fngWxeJMDvhQYmlZMeQKpl6FMmzoyeWH+fwCi23uBJ26Gq6nJPGYDkLDJSSpxB5oi06Ly7vxIgUd
sU6as3Ab7ZsLgsGw1sFUPC2Jz2lfDgfprcNIWx6UcNZ1c26yWrqae/8BfYPNTvVayRug4Xh9t0Dz
Ul3p+hg1jZprjPiDEsHIfbZAJq6qVSdtriJhxSrspcreRPuVeAe8SPhZZtZmgMcR7pJfaKlAZYvs
6imukHjpfdqUwjzwztj1+pOMuawmSRSo34KZu4jNGchIhhKAVw0QyOMqmcfmKjgqku6U2bslCjY6
Gpi9aHppb3wSW2GxaSN4uwXrj4wVh3ME1Ohiki1ng7YxCYIvQ240aAMF//iFZpr6moaL5sd2abZQ
BclDahEdxSS5HKkmpFAE0LiFoLpd8kH48SLx65aKYpkiLXG99Qx5Nzaa3VM35PvQQfkVS5G6g/AS
iJIGrO0/Cn5yJP78VnlcvFVzGiZANXdPkwWue/JTEeKBM7VJ2Ahwtc3JWtWTu5niGcYqftDHbt84
n1ZSvxpj0xoJli/O4SMEzmc4EWx07SJuUxGI9cK1nBi0AH8kNhH2aYrmdncsgGca3eUcMdrkn6No
RQB4tYs5B5QA/etEDg4zJs1zZVnoeYOM7mxUehPfgFOdW8QEOb5zuKPpgHKJ8MBMOM7FNN1trcZJ
W5mgg71c9e+M+bHnYhsmc2Rfk9YKd1rUAs2EXLYLeqExyM0ftAW9uKuyKYuB5oJoPujv7ZQvQXMP
yfuevnIgtS79BLfEVI5Np5FaHTiZgiKoCrpdlJgQ7xXsVf6pQMnqqV9eK9AD3ORVg43fPTiZ10AW
N42Yo1ye8bTATgtWPGnmtM3dK2asuxp93mEPEvmfCUjLBisMKQ3kZapGjXIUIgbA5wjQSQP3PbvB
RizWdoX0gddMISXwXflDV6RffTmcAjE96YObOvW9oin1Xbxlo0ZNUjsvblElvuNxMCDp693LHJ8i
m/5YxZRXx2dSzU9rqxpodkwJC/iNP5pcag9qILDJKYFHHhAVUIoFKuMIsKx+sLm5Kqgf0QZYZTUe
n/JXvMhc/0RJ6cdQkc0C4tl8ehhhkMjS4/TNgUZetrRzF9ARWSUrMFMxpbX31i8bXyyhomr3WRjx
5UKJljhP8bmZci6mmmTa5WdYTeQ9p0b3/HNewnxI0OKPDI8S4CXKIPilbeZ9bBDQ9Sziq6vKVGQQ
ooQVR/IYM3WZ6Dd4mLFwsgTB1KPA/riAaOmAg64IHYti5OLkeKASYR8e3bwYehranQ75aoAUvHhT
/DIkWgvzA8AYy7Hoees4WXYQQP/iOVzS1a5fz9SSp1UDOuBhTpr1geeCPMz3//tZvz9w0qZwvPPj
FKomt+mxNrCFsd2ygMusD9vDB8yW1OX5on2GxaDb0pTjzTP6gBTwOxnPsum8vTwzeimL3ZIH88lJ
6nrIxjr4cfuRExWdCS7+ekrtbWHx9FcJKz6R7D/Je+naaQFCavJa8B6atqrG3Ah+e9c4ZM9/kcmy
FJ5nn41UcaWHGHh7ahLmgdFGD+q2UIayFc4YO957X8y4ghWrWN+EPNvMrmolZ2EBBwKtdplSw2Og
B1QAoNLpv8iPFqJ5soGVuSLwkXTY/G1+vuaj6/RKv1sp9SnIvDORIS3+KGwBNAKVWNdr2s1uRIzE
L1eWhqeSTSdHmXtrbI7H/+0VsQz+8guZuxLQA0h8ljk2fRElcsg+y4sj/XNPEV6SRzhmHvg28WVP
Ph2yJ7DxI0pl89LQd0K5DpmxoHVDSwzZcUhA270kjs3SShR5XKfrse5p/L/Xs/11TBELS3/dGq61
ZN4b3H35L5E03dcvQy0E9lDfKm89zrlyl0Vo5LCmCErPZbEHyboHDZ/btOdqCwqGxHGOacVSSseQ
mrvh0iF1pdYfEupWLk4h7gPKa+AB0PrSLRTI6U/ay+CN6ebnmHIHvjYX3GmW3yWBYUfAkHK5jheI
OH+l21BaCDHhz53y8encVb+1lyxLk77mC3LRprUTLLty77SUa8eLdowZHeOQ2xijCPXyeBhRRc1k
CaKlMJzuelZ6GwXJuYcriv37dr8PPP6TlyYneNdPcMPtdzNWnXJvIuUMn/VoRwLxVenRVm+/3U6z
wNsP+fsL1RcQY+nSWeAjtYFsUzlKFmUt6PBaS28u+rXqz/RtC/F1RVw6/cdN8fPdkRKwmag19SBF
zQuQib9gM/uOThRKRkDtNHLFUTKcxphUdUizbJ5aMKIaMTk0jsrNGuYZdosHuWcKhZEdZ7GZ/+xm
x8kmzmQOmdLyQT1HPwrzIaEZr/7pM5NZtr5e6uAO/02N2JxjnNAR1Y+KRXKscp4NZJgYQDQrARCU
NyOmm8zpn+1mu2BR0UhaxmIQKww6yoEUchQnXeE7hkttucgLoCQZhRoiiXnT6RDDuDLRaKqA6xHU
PCkEO2JWoljVov/Fpo3PK7v7Zop8BFUuSc0bRlB0j7Aa1CzaZzAMvfCwgRmHSr07wxwfzL4GRSjF
xq8OIZjVhm6gKGV891feph371tA9jGLRzThFsvG0j0VvdONv5Smvy4tNXeZzyJm+VljyX6deN2Og
QoOY8J+f8tn8H2oRZVP+Vygxvz5W/MnaOBtqxJ+o9fpw7l9jeIPk6A5jfmBN0mb1r9MR1bIdrAvo
enHO05LUAFTncz8Lqroiri09h0xVwDDAodJlUSnzCohjld89pFRaR2xlqXWNETWFhS3oBImCC35R
18ZLSD54JnJvh0q+RyIxEzvpsnYfbjCuLkVpJ+4gqi0sVwnLD/airlFc3vULeHIj0SFEWxNW6RdB
3IfH21irwHXoKoDOs2JEtl9lu5tfI8sqIo19w7i4Kovh0a+4myj8i9hDUZD17lH+Zsbeb0RFmunD
78Uz3S4Y8dRC4BS5AcsDGMusw7DZtqYzVXTyQqA5AH0YOYi8hugzwifvppU7n2rdTcdMtJo8hHFh
pAq2HLBKokVsDeFFZXr3ZgBB+sVhyN2fdHrYSZiZ8izdA8EP6qxixTLc7sz+jHWfrC36Ui4AZwWu
cgK8jcYCEPVGFWjbmDD4uosgQeCkNhhIYGC+X4KujBBA7cSYWUkHomCqafq/5Dt+LQTBRYEmL7eK
nwy09r6yJFGuhF3qcxcBlSn50zY966G2wOJFABW5Rt/9X7aG62xT1cHbBvr2ki3giMevuuzdsrnT
x8YKeKTpmOEjM3wRdGOfnSblrihR4DKrewI0X7W8o2MTDyMmRCtJhpONFNhGNsuCG4SPxYJ8mI/Y
s1m1CIdxZONJxffZZAPUnl6Iagbaz5p09ad51zGguzI7ExVMZtj3A3dMof4lC/3n1BsPYU4a/gPp
4E0i3izl1L/4fHRWF7mqs3uvkzvgwu2n1V8PW5q+pH0HrWYT38g7vExwivVumO1y4d3qYEzZUuRH
j5lg2kSI2Gt1ZerDB54OR8cqU4pafaZ7K6NHF05tmJXX/GVP2PW/5jpV5mbZsYwjRMD7sA4i2R6x
204g0DaBLj+xDZHYsBUmU6HnZ1Eoo0KhHMW9c4rEwxNE7W6raJjT8ccBZXs49iHwxD+BqIAwYRVP
7MnVcLunVlRFN/6gIpMhXLcAPCg0DKF0kvVG2DfsDa4WZf2zF3WjZ9tW+Dh9ZJ+pj/HDA4kBpD+Q
OTBV8AUrXV/S3fwiYOJ9mQvw5mqXJnEGmpPYc1mYUFBVIeTbEXQMJj/h9hLGD94hWW8wldMWMsJI
A1BuqPpHDyIBAjnfwfMiam6yOQW9+CyFZvpWWOGNdqY7K5u+1sMVOQ37FUmyllgJSL55MxhD9JGJ
v/z1axzHuJAxi79JMmiIM/KWIIS3cufz2bp3np9WInGlwFfs7PUhtNYgm2TShh+ENzBpZILpMrxP
CBz6nCEefO00PhEoaO/z7h/SkZFsU3lnbS8OZULLeWKVz7jyFvMFMVedRP3VAgIxB3DWjK6ADV+r
tnU/uPmVwQhdHTXwFdMAS2EaxjNFqy9/EL8RENYuYNjs5mBs3tO6h/yLxV4BWcvWLzpG/2+WbA4q
UB50ebfY/WkCSvOlmCV+b9F6Wfi7xyglOexSK5AxH8FC77EmG9c5KK23uJM7dFA6i1YJYNIH8Kwu
6syGvxq9twblwqqu4a9maCIJmxJne3tRLl6EOT2qyvC7Cf2BdzEHA3InwIiFZ+gSca/VJ5pcfhCA
kEHZlbfn0BaiFF6lE9qRGAKbc2mB8XdanNnUpk2up9AINIR2Zn/u0AZhHQ5eNOFnCLs6Jnds+k6t
wlY0ljjfqwpwgmIlT8WEJ/+dooByUvR2vKBW8aYZxdeP9ha9gYKsByX0rCcvOEFxJy2UviZBanvu
EBDrbmZSrgJCd2OG6eQhDEXx9DMyUfLPKa0AOFGjBOSA572IxOUzUlQ3QL7skesDN2uv5VV8+rv4
C2czHV5bXXGtx19quPMXCJ5Fy7WZji+IJdFm5EKKkB76JAlCbIRS8QWIn0NNzMRPV1AvRnFeS7Xa
FJNHUVQILSSO8McuTU9lXGJ5vyS+pJcYaW5c64LjENJh6xCEsL/OYCfb0i8L05FxknJLrUG+Qxn4
c2nZDdwCg7elWldSygx7yrIn/cng7PSHZJYlcadM3naoWSziC3OqPb3gl3c9KMxT1f+ELC43UsPp
W9RFydX5m8RvWEt9B1EWrrDb1PLap+lvY1sboI3eYarJ1gdAaRr3loke1RLeFDoW/8Z30t43TItB
udBl3M47a8VXGcOClRwK3VbIMifwIE0xjQbSohONS08upaHxr63YEWW4IG6r3c67FmH2UAvLba34
1p58dLPmQ5aqlFV6s2Ju13UjjMtfgWu4A+/Umr4tw2zc4LcKWXwmVU3Pk0XUYUxPNqm/UmiU2sGa
AxkFmp0Xwt7v2l5oza7CXGZBFIhlF2pcJzdz3Grwr87NYOF1mfPMc8SjZRIMKmvLB+2vfeyCo/hO
vrTx9vrsxJMCzdXut3qcRzj1wwTwq+6m77CeoJdTG8Gw4swgTyDO+fXQpkOwUh1mY6h61DhFwLyn
MuRoGSYyD3DXocsiXIOn8psf1LE4Ora3PE4WlRnEROht/KM/J50qsgs+LmWAROjK7VmKlQ6LFjmy
ueXhYW4faC2ZKnEKAVvUFM1EuR7ZroQVjs4M/2cUF86fk24+uHTvonVzkDJ1Om6FxXzWRebdAKCG
JcpaUVWR6pLwcNxyEqK6s+b+150XwtvcQr+kq9g8BnS/jlfR9YfuRtwESn5Fyt/bqQHf3uUf4MZr
9mK4z8fzFGVv5ri36FN4IAyooSwOVfl9D+/2/+qHpwTlSHtaJL55MrJ7KRsBtmaOg+6a3J0AlBvI
1RpdVDQpfs4ylSSZvqmjeq+dfHrYxBj7eO3btCyF8tbYjfv+Edl8EfK+2M3au4Livvz0niu3fjYY
j9Py8B1jGm+SnmTWs6tk8HHR1fBdCM5IJAjEY/ivlU2akHzN0peS8t+sekpQamFivdZ50jTYCNPk
h6pKLN7Or27OQFinVfIa3u2bCLopp/nOVEoF54CxZc6le1FEh5LSAfeqs4GUzhu/cFKLhURCg3Ur
99Qdjd3Qc8mxuiHvu1588wMRI2E61Hd+J+CrvcYMGo1Gc/Hf+cc7jwASOpTjYYCWIUtH6rIsPISJ
uGDirhorRnSxmaVb1+YmL63+QUOyZ8TcjmjXRMqYMGREqKoF6Cmro4BZY6M7mkIfln4jZ2+i8MFh
Vr+jrw7rPeoqPcGcPsOL/EaXQy4OvxxMSAVoEwTusx6Imsx+3bbWhQyrPMMuutfHebykkinHtXiO
4wkysAD6oFWOI7lgNFo9ZVgUbFHselKpZOMstSFRfYNQ4Lz+ytGX8Ojd9szxXCfkvsgAXkENSmFb
EWLUBIyI3/6/qMObye1FZAdCZgtZVvPJzSrnY/2MoqXfuM/aL+ZFLj0oc9MZhyV2tm9Thnf02JC1
+0mXqTvlCcgTozhENUJi13SDJoIPpy3q3+vidMGz/r2wdcuBag9DMso4vZ9ZCHN7deF3xyKdtP+B
C63kGAu8biz24TX4mf1K2xPXy3fm8N9AwVkCdPT5eV0NJAdIU/muR01j/apHzRzAu8siEkP2yr2C
0OSHbL2sEHQuWtsgOaqMLPeQNLiGaxdzoI8QS2qB4aTgrhtIr5tEKiGlbVZyKUCeeeVFl2zvPkSR
DmC3h4Aq0V836bfDJ1S1usIEW4A8fPwT/hrDhijvLKbkPd29OOTwZNJ1jpiorwPF6gwaAW7y0BCJ
sf4aqAAImIELo/mq9ojfuAgngT23GhYiIIB0nF3/4P9t9gMaxE33PgUkpVoCIcbR0G8OOpPDPZzS
yIu7p1RfbUMQG1f6lUEIoSAmT0gGxV60kiU8HAr9RIJDFGF+5YmcQ/wnjG0p78unbUvFEAsjGCOH
vNixzl5qYBy35nmyD/44k84jxERcOSSSoC/8IzBRcpqM9IYl+46R6+yfcionqM7Pd1ie0qaj9bem
F0v3iaSPsfGgB7WfrFE0lnLtNpjFKyFIhA6nWYY64JmdqiGLiQxnD/I+gSohRTm+eIiN41qYhz6b
8xJtYSyzGZ+YWAV8VRGHX2FeLNZ/QB/3r9n+Xl02PNhc0x1WNQEp3y5uOTjCV2MxiUyW9HRzyfFM
ngOAR4dZPtNjJC/qvAAZxXucpFaxoC4gcoH0nEAzYgU0pJChq3nipcROr5ZMhD04+V5a2oQ/V9uK
hAKIZk5SzLUOiQy/UXNnjiPZfQMLRdP/n7tpADGqzsiWNmX+4drjvO794k0fPUsbiwRYb/9Sbwo+
rbwbNsuITXUX5bfuk6AKTQZnaamCDger2zhEP7yIXa6IHetvuDW80WgGvvaN2Qx+GUrSMHOgTVJ1
1PhF8MeiEMIdj1X2gH7oc8XG96XUFnjf2v/adqpLfBD7ab+DnftEdT+70V4ZMv94aoAfREPKEFVJ
MdSGZrhMYKrboEiRfVY7c0LwgZvKksk3ccj4z/wg3JkYqZ14D/XLG7QuuA4OEOS8BMcOBkbHqZSF
n3DWUBJgApAMxKmqgp+wMjvixNHai86+1b2CtKCvfdpULzh5KY8q0KeM1wcBuF4VzBcoCgMw4fu+
6oDUuSkWOvbjkAi70b78KA6CsQbCnQUbracY6YzP7UkiDVmg53dyfTYcCBzhp9s9+cQtPXsaD0Zs
eEUcJayFYnOE4v8nCcAQW4KnvDIe+MaSFI/WZGibPq8J0LbaqAS5ERIEUZ0W/SLLgi+/terjTF02
JIAOkOK1DIsdQORohYWtHK7G8brpCb0M/qSWPRqQnz3QNgCnlvNgKhZW/ki+5TAUHEK9+3JS7FqY
0g613hcaQKKmO8nAVTh+dt1DumCRV2XJSFixujjjcUvrwrQF6h9feUUc9lCAYSpTfo7yfmAOegpX
zwXy4KDhss4mLEzM0GurXcmTqU8HyEXuh+vpW2nc3ZHUauO1bBFjYYj9ao7LEYSOnQ+H0IU6tg0U
iPtPGvTtts3L5+LjZRt7zmTboJ/Tg4OLKzFSQ2N5b5Bo8IlYDx0xPm0KDSZBXTXrBajmb3hVXDz4
4ysP60yEZUGhYhrfgMhPNP/n+iwBMWUriF1maV+Fsqx2UhSDzu1DrC3IKuNttRqi4fLdhVX7+VMM
Th7w7dshg2r0IkoY1aHfEyLm+csfTUQba2abgQ/08ckRbdr1CjIjHjzWtTFVyAuPE0rIHsenqnrp
G2UbQSGGSoRZfi903FJL8rEDgiyN+aLGggsrUjiZTLGghi+VXZ5PMd6rkZp3LHJ8LvfrjbtF/hgg
O3NArVXYC0WDS3DOwUpqBohBdhKazQdJncxqBeyOdAyCmOzb/P9vFAmMUIa9pR+CXkVTs29zbmw2
JJOq1H/jUTkF98QcVGcnqP79FB0IrdlYp1fddS3Laxsm0VflnZG4uQ55vbQKQWWNKy1iIutZfeap
NLRDDpE9Sa0dv/V+N2O6Na43Wag9YYnk/ezQMtjrZMEff3E52p6HX7WZwMNhgSz9QFwsJ2K3cMo1
d8BA/piDxpeqs4fyCBve1n/0n8IFXJPLOIWs7gBwn7JEMsy9H6cU0Qh90z/1XgF7V5kJuWRhVVvp
rBj25OOTUNP/cpvB28SL3w6Fn6oUdeW2tgMsbHyFdwWug5oKrgYJXMDYsO/3IcNTHOXpVzViKJDe
IEw2E1tUR0XVuLrFDi5RH/NmMLAXkxTLLamQ7AIqktLy2c5eZzflOjcYFWZ5spIOVozhEeONWvzX
J6YJQs9MiCyw4sDpGZeyVBpcMnP+sG/KUMSWveFug8lPdOqU0B+UPRKob6GHsq1eWo1maNZykuhn
oMDiTY05jwS64Rfi3smw3l2q9wfSKbvMrWPbwa9y7+Hl8OC7HZEE2rBFvxvfdLrgI/SztoM8boPE
7lr0hD25YEwtGC2fCdFMV/5EKaD1l9Qfl1Q2JPqvXnzTWa4Q+1SehMz1OisV1KP+sUD/CWeKTWNr
M9uOkem5XUI8jIkF0S/vnk2Xww6/G5QJMUrbBzA8OV5EctEg/yKrdJV4WfQFHlowAKQVqRKNDnOm
1mDIBF3jVuxQ2pwyjSYGyMWcEmdY62aNRfj92hyBNjWJVmCR46+I0PYlVPyrFF1qi7niLo6H0N37
eWwdGLumtsoAuLHhssylall+zNkfs4/v8fJQwrQi59b2ysa8tVk+eqvSnVQZPuylOtECQ1XV1Ue7
jO16Wna616gONDqp5PzZUThef+khTVEfkx/lUa4yP704njsoCnA7a+tolGfk2ViKmfXCEa50BQAr
N7RmFBMfGIzFltOy/ArdCRQq3dTagz81cigS6S6x1Q4qYbA+3Z5AeiomkOMH/l8FSc2r6zrdDFh4
ZabaiYvtzh2K/GZSlE3yguKD+WgN1MtDDAtGTazMh3zZ+wXMaZK5ZjGSRLJpZonF/jQ+QspuM2u9
AXN1N4Hlp8IfgEd9OBpv03ufGEpRmQT4+unZ7wyjDv/3s+/+u1CCML0kG+jwXxg9PRAviqweFltB
Q6xe/zb3AlHxmReErq/z46PKUWwEWrBBP5S3MwfWDP5V22dOfBTZyYO3mXLdYMkXinaS6MkWhIk8
h0GHhgnnUVnR23Ab7iHHNsA0AMd9n7Ary4BJJDfhk1oAeA+nWa3wDI0oUyq5bgsMTxg750azmExE
dzPl8hNl7nKNC/nWyRpEpfLMlMD/X0yyf0HFA8M3E8nv8+noKTRKrG0ObCAdVnhHXywsxSsXcxXA
FfJNCQS2gUrVF5wvJVvEC5rA7u89gwWoixfYmH1lGOJfMEzwBk0ahIK6VPPtLm2akNiDxlRb3/ZV
brO6aaSLyaZgXTMBSZ33z+kHWhpKkliMoC2pOs1Lkode3gvgkVRTeoKfaCgU1BnucNlyor8KHjzu
06f/fYkbS6X531oFBA90KWpcke3dUjYamCKk4Xl3N3C7/CiVuu9K0+Fsxalj6gApLGSH+s6C2zqI
tcIJfkJByX0o9SzX7vCkkX24eQqBgNpuh16G6KG5ZZrDOXrUUPgKVgpy5HY3Eo0QRpSV95wBcpfn
uZlA5FBvEINijL5zEn4Kc4lG0jUnje/VDOxfZtNNiF1bRhRz6BsHYMpFJduP2PJWxBQ1kmEg0Eci
QFCiRgGnQnkBVQxLMbgk8ytTynlJkHjspyjjSjQckdagyQ7IiIZYoEOqPraNB5TUWYOs8wBEpOTL
qNVcR9GUu7J7VzHOxQK9c7D8MirflCF3LkUGqQu1+5b6YFulj7HKnWP5w6vi9l3lUB74jVBEVILe
bJF9o4tbWZZtboFuHADtXo12SPAHIPS1ddnw4eJ9DvNY1OeMrq/6BuXwovQW4VTzTLwFCDFleHVB
7f8pdCQLfAhMNJRjbAdsA+92BQCzT/qvRaiE5ODPhoOPcqPPaMvvZf1AvioWoF2gOSo8Nh0KFv/T
SybRcKabyE8cHy27w0NRGfW99m5awuiNVhCZArNEp6ivaa1nrFf/Fl1S/ijI6uliOpqN+CZf6U2v
bA0p7gfKwcGdQgTdkUzpdd0tdfXRb2sylyfqFChJCVOt9BiBkVCkva2HsWOWOat8VUyuCwfPSLUu
xlZoD/JLk2ExJ3yCu8YttANQI5XIIgiEvfVhxTnKTQhImOI2Rmng0Fn3PF2w3lIYrdi9Vef5Ujbv
6XL+25K7VVEaMlTVXlVOjh14Y8IDNqWBNi/wFWcluEgGSCNP25MHaDJqisUNu1/7W5kZN7UKkDGX
tbb7ZclTRcp/PLLpVFo1N5+RCx50c1Jy1vUYAu9FOKFTVcpFdfL/BXEaqtk0ovH5Qorj3TDSXyC3
hydefhVKXRK7onxakSMDs6iOYI2hrN2O0l39V1PQYJwS40wfDY1Yr4raLolGBdCWJxC99pxvfE3G
hXKQxcF44ZTPTYcN9I2OsWTeGfFZS+NjkiU3+BezRRtv70t0wrERqFZkYaFd1B25ZYH1siTQh6+H
EwZERSdXjaCL6tDAxrZBeMauQ837wXj3UatP/uuWdxplqMv8Z0l7iybHvqyEwsTGC+JkvSjEdKv1
04Nmjn9j2yC9erDBFdP+9xw4Smv0STC6pSgwqqMzJ7RoKsowwoLFnz55EMJ0OE9hVA8LoXqfmHTj
l/bBY0H3T/6kT44GwgqsI/EYK3s8wXnFwNPS9758HNlBQqJ5/0oYFEU6j6KPh5vZhscUi3hE75Jy
ssY+GcSsx49Uprp/QfmmYCuC9Y/Q7wJli6hbR5uwUSoBQ/aYglG9+0I/dpi72g/BHQ1BwzzYwYrF
jHCjdQGMpUoiGkTRWH0G+UeAV0O05kadmrI4fV2nVmjGsUseoMzm4wZ5IzgtYsFJKelkUB+7DZfM
djFLARt/IT9Nr9152jFrbSn2WAwq22lXSGYNrG4ZVZkw31PN85h3mi5WytHkpWCz92juoxBnE3ih
GXlKUcF7kTR1S+kW2PbykjiBmcj5GKrM0NoSBN/kNRyYL7pduUcaR1Z7OH8sd2b/JZiNfui+vmiO
FjEWTec5IWdBM3LMYciZYX99P2rZSY2badbUlLXHOZhqMD6Myy4kzeY+jG41Leou3TnHAx1GBisc
d8HZXwyrpqXNK6yayWIHih+yPUlQwyMVMB9ENeoslRA2vY+/MtjDTthQnI9lGcgsD/KYhVAdFr9B
uPh8+loP53mke5jPTR/oj4RBTdBKBlUZ7wDcy+QLxfxW9/4AjFpAIQERGoj5TUKJteBwAMBRI/m6
arnKPK5KB8BzC43n7C58EBde4eA3uDrss0MnxPlkWc4BSFitCq2kxPfI5s5aHIZKCth5W6TRdPQX
EDCmLp9jl7Xza3u4wXlOMKXaPdjoc3UlXJV8b1hkHpM37I0RJcVrFNmSjZxFziAuweVku2+L4/2o
cUJjq8AP5ztj2aK3ax1QEF3jniaHKJWlr1yEIvXgghr1cnZtD+SbMOJ9bpetC/EItBrJ7rawp7x+
MLmwm23mIWy721E2RPe3vmDSlPO6L2Bx2FmAzpw80fDmyaX0LcHq61c8xEu6KfnMSnYmL00KaR6h
5zT8IGCpeR1AFeVPS+vP8XvzFrJSO3ERx0yLo5lcro+oOhj9/j+/u1Xb2igNRvpgarrQ4Ez4bPlo
pVGjuFWH3AUoaNAwqGCwT/fmkVnbnJJYILpl/+dVfY6vG+Yj5jc0dCgn8wTqRq0pbJc4pwp8U+BH
FPB7vWPu2HxMJJINwu9qEjBqOhcC/2WgtGf//kgRAxFNCngxpFtVJrH2v29c9vAbx5JDh+oxG4wQ
SYjjWwTJy6af3yFETB1fiL+CafB407Mx40ZoY0/lGTY6lagzTYLYJoCQN7FIdKtwxGDW7VWiSaYH
BQUpQDRI7OD6qQODklZh+TXIRXukMXU6CuzPgURSZG0IvFu9sY2ZmSWcxmeXD55oQuFg7YNvY2Ad
WJAJnQ0TE0Y5Jeh3AXM3C8WGDrwl+H5mu0cQm3Kvmc4NCBQzgPwyRl5HwfbgamAOl8qBdo/LquBq
E8li/93/1o7uljZ2IODcfDETDPnLoIUNZgAMZ0GshQHb6CgwrnwiOgQly4QI5kXxD5ph9x+SEmCC
I0EF/4gUVVaNPXFG3eimWRL5nKlsOgSE8xjQMPMM/AJZYcgY8NHZVWiW1OtzeYFG/aAKSpFKl5xd
8g3YGll/pJwiosADGvdVjZevB9WpVC+rjU632lZr0NcfPn6XwTtpgXbFTJUOMwlqnmSJDAacnJXK
ag22iHuUHzlzwf7zoVDAs0EaI7yO43R7UCVXx+eUrvZFj2ap7+jGnd4bemyCnwRhEG0iOSXFD76T
v+1ggCvsjZu3R82EVOQ9rbHS/PXPTQAwe6ojdoxOXv6Fv29W+Enr623SjorjiR1n42gDBhGYRjyY
trzgnDB5Ozy2Lh5C6PoZ1BIMt+EgptRqSqLjt4Xp6ZLWkCM6xWDc/5yY9jzob1RyV/SSkk3ezu1M
VGPZHqoAVTFwM8K8U59ZChRqyOjPInGIruOyX2/cOt6uqwXP/6iEYW4lplpEQRzwEzfRo54AzQMS
hXD7UjY3lvxT/hn+XmWDTxmJHKuRiGq0J0Z0zlXbosz/Whz3+saiXOnhj84K0PKJeW4gX8+FZTrT
5q6HVqXCj6wTASPf4UV7LMjYP+B3ggoLN4cjgyt2EUhtYd1wN6aMYW526g06O2z42pnG/biYLeu1
Sk+Bvb1F7WsalkhMEUd5dUPNKLSQv40q3DUBo0W90ZsvzMq98oYv0PRFN2WEwMAFb5N9maX4droK
O2K4XK6FGnPH5rTTM+ENUxPOH8KcRgjpSEK+1a7ugv8+OjlT2Bg1+nhCRK9D8ZaVkstrhoJ4h7F4
8jwTuZJu8jc/WInocnNVQjzVXYQ4g7i8seMJknBo6xsv441BVIfG/Ws8vBrFUug/K7NhIxR1i7bs
fEB1FVaV2gPYDb+SXqha/oUsbH3bbl0E5NM1Zo4uaY0g4aPFkN6eksFD+BRS5fbAnTnI1xyXHK2b
r/YVHVzG1wRgNz7pMSzj1ieUBI03x09Mas7xppL4azcN2EaSm3hcrvxtvlPl+eT+zVuVrYtoRP9S
R+BW69hmvqLyHdSmcgY6/DdLieXC9DtzTJcw5Vj9rWP9imG0/tN0HKh/fGAFUEfwAjMBK+huAeLR
6KSeIo0O/2LBh0OjXvdQIhPx1Fi5Qgk+ULsirkUMtunj9Ox6Ge9kQR2dMJE9rdPGQtGEvBoO4z4l
Y7spzYX4ns1tkKm9IzmOEfotT41C8nVusuzBscaQGhtho34qUs/SD5OSQYSjGe1LsmkCvq+s9eJl
C/VKu6G7qfKGj+ulsdwEaXJIjOhQYZfzalqat4wRKQgTEpGeKIqLDTmCakXEXQpHZXFgVrP01GE9
Xb+sIEiUzaFOr/qksmfcKewKH2uB2b1reSWDWfg7VT03CKNQn5jfXabporV6ukS+6ynMe77YwWLj
XdG7/9BmN0S71rwaZg5YFQxJqUx0nCwNJ8gL2w1IBopMNkuDM28akOURMvXUpAX5stUHJBEoJo02
OGcrbY6yKDQtv9H+xJ/sfYfM1yGyct1Z+xfnoeQ2dFEuKVe9SOh8nSoKbA8BuyExJWQvHjruxwmh
psWQkCNkEC0SgE20G2bmPjTMZdkR1ORayAmfQ649MXSnnfNCD8IUKkk8mBiDvyJM+hbYS30xs1Ha
48M+7AFy2IgLKHA/dw9RXGx0SEAfPRcwVUw/dtehn0/g6YywV1Qw5v5l5riYFZhrGLqzg7uc8XcY
VmwnNSKBySl5TJ+XJ6PLgs6ICib/lqMczaDmPIhZcQT3MrvOk3D/2PdLgW3wTi0qbpG9wkZjQlRW
Lc/uonEQd9ZJY7d24ColKD1cHo6rmQaa5BDrNKFBB3dk5fyOyPtoTzbiBicbYtDeem+OLhICmshW
d/2ab3dU2MtTkA1AoZqpw6Og0gs90H+Nbw35j3ol64GGxwLU16OYOIVzM5aoo/z8xWhthGXDUc/l
DaRZPcxzWdrCarFhMPCMyb0P16QM8E099Gy2g6Fx7V1rT4eK/9mTER7CMObbUgg75VbSL0FDcwRO
vf/bosdeBR9vZJKLG1rwRHSqKBugfD/aehOR7D88g3U5Zvoq5tJGdSIafDmFeYsDqN6Uci+x3QPd
3NumMl3bXptD/Pl1rA0q66fGCTZZHjp6suDJNSJIbPJtO9HqpkrQsuBnbKJ7FxV49wBv5/kCMqSY
B9SbjHWKnH/8iDERYPeT6LM+H+oRXXTzp/sKGH9asTJ1w707mSTXOoadxm8Wwn/jFgLCdH9fjpaq
PN0x6q3SIUCX7fhZUU4O8umLC4xWVM8k/lxloKEEXDxgpF4QrwK4Xip9wbeHxsOrKFSm+/iRVY3/
1uqxA7JhEiYaNieJLi5ZgHk56gAueK0RZr9NHtK47/JCeFVXBXyoCHAeaz5O919J9j2XfXrepAwZ
R74uqTZcavInQSpdc8Wg4IrTYbw9CxBSq9f9/kEI1xPWU8AQnCtgG80a4WazOrIibgKndoTXqNtF
aA0MjW3Maw8mq+IPg6/OmXW2VQrqE6UI8nFQdP8Q1BlzPol+0kN6YJmUrxv5Ipirm3S0BCpTQivl
tyzgWcC9oFAI3sOR/tT79H7DbLiEu+8lTFqoonOGrm6bY3co+sbAQTxHvBhdHjOOISNnltZQTaPv
yL+L3YtGHmkIwh0+fDpm3rVTXKkYw0F8n9weQWfoelSAMg+hUICxqMb39gj4texMVgm4e9tHBFBQ
0Ff9JbN7LwqWtrpFBMY6M1Pp7UOf7sniLWF/nMPeXLNkMNuoAl2O/gzsB8180VZajTeUCpagtprO
UExjDuFzMRHYCWzXrSydNWnl4XKE0j4p9rv+rmjGSxnqo2QottQfD4aA82FJ/I8i0gJuqZHt8u0N
BdHh13lwQkU4/AnjbyoryD5eR6lrARynX6Qa7eh73BhvkzclOOvwFHgkqxdtaiuJxmccRQvyKopg
NWrHXj987qVXRu9TqP4RuNgOf375iTONjD+nSeac7JuftP715FKdlykdv1sB4lZ2jVgJvXQwcJsd
Lphqg+H5pelgkhYcmcTlcdhPf472Q3sbin9gj9ffiKgpuGemDaXjZ49sK4g42Rfd1kPZeghx6ABo
QvRGM+wDFGPqyWZSXexGsEy4vne/zVF7N98nLdIMNjsb+PKsF//k3TeHX3DTkYXIpuV7DLMcklha
mDnnzj8Kw8+GX1P9UOLNSBQLIrmZAnySSzg/VZ0mrk/tHbhzBrEhCRJCKVaLpmQu+o8H7WlcpHfN
NqcEtJQ2snuLAw7DQDzbYOje1Mh2uxk7Vhu4bFbX3nWiy/+U4owvowh6Kr3UAmli1N3uT+7P3Kh6
GIEQ90ds0wEz02o2qbdnZODmibrcs6cvC5Oq9zx1tSPu3Kjk9cOkF8Fq89YQNWGGOSurtBW9l3Zs
+1fnTR8pZ3xHqOKn0H9HGZineSOAqFbGFg2yCxA0w9mZzFLCPGJ2dEH4JtlLWB4l37N0CXk0MlXE
6FCxkUN4jm8sZsfvi6G/DudzReUD9CwYajMX7gpBabW0rvIZVyGG8EI9z0cV7dE4JSPks49zpjTx
c7rDNjPAlzSWu44GFaBKkz61a9HQV6sQac3/5ZdferN6vRrwAW3XA32qIKtUxWSyZdjBfk9ZHhjG
aS6wdp7h/IhTjXPWIqmZVsI1LAOGkfzXyv5+SNtptc5yaTxzJu/KlutCr6//7pZRxsyTYO1V4yrC
rL9ldHVDWBJ5te4vfNoFeR5QTfAzZ9r5JKFxUoD+1FwOuFBwoTsMmR+evxatEaAeD5Zv50UsWp9J
Pa/21ZNpHUBmMMTOevvN3hsBwt3V1F7AzRS+RfZ+VsYDFypsSWiR7rGkHEHh3C0FZzBB4W0+0HU0
m+3OCexwGX+CQaCMqKBcJoy2bwjZtH9z3/4Arh0sW+mmFieLjvcJ7GUMVp7BLC+Ev2zeu8pRIk9C
bt/T8X6rW6/py+b1Wo7L05yLuN7o1U9gCwsFN0prT/9sKVDctYvTG+GPT7MCUVApZZe4tsITnyJ6
6Ujrvf3CBN06OGfI7VxUFvq9PzLqCKd8HJH1WH1sHu0oHj2bhJ9ERTr6/N7fNEKIv4NH33HiC7Ws
vDroyBBHfUHLto4b228yiV7IXy8NVHn79018KhUKyEsQsF6ka8ouBFShTMvA3TFqWNfmyLeRJRlU
w4qcFVFjRKKIeYUZYu7DlrQA19T9kzUhMMagrSOKPLlHgZCmN0YKzUx83UD+1chP68GaSBsa5KHA
tDwtJl++hZdv9TTX275PJkAdAH23zBqEKxdyy4bAU+pWPvPvQXST8if1nfO7Vn+/zK7uhpZIJPiX
2bLs2l1jFZVkmSzkZ5hYx1ag8/eIfSUPQIIGUusal0nUWJUGN22GGmYAKdMJ6uM/ZHn2eIMK3WVK
Iv1gBXXTDJ8qNtGIRpeBzQnUv+3wHJG7DuKYU5nyzRqH1BEC3WBxuP+DEWlftqssQdUnQXuvRbTk
XmV6L9Cpg8lcKBKNTnE43sSwPMjaw+nIj37iBhS++cGg+9Sy3yv+3TXpPqs+8e8uIUdXKJf3VkOb
mds2k88ee8ZyHgjEzN6NGrMpbL/ibeGh5dYJmJdkpDhmehbIjob1Ars9VV09ZQOTYl8KDK97+0dV
WU00J75jJfSvj7x8uua8k7qiK4pqm7f+VgeWPjbuU84fhrUjKc+YleD7ivp6imGCSftivdE1G0W4
RUEGrojFLrwPsSLtXxAgFmFkEEgCQ9S0IfAbMNmD7N/pgc+MgF00AThoq84a5SSoXfGoSdGgFsFr
810iQoSAcTVnSKZy6ReCcbvBql2PB1L/ElR7AaYHEv2D73aH6O4sZUZc2jERFalYN6qPHB8a9MSV
rZ8A/ThrfFw8mA1pZGe0Wzy9z0+5eyWcZTAcpeyz4HFIWEq+g9KOKuB3n9IVjKWdYmCO+gMrXRm/
LKFUqhcW1He1N5ThMIQN1k72dElrpssrovVItUtc/NJ0aKnyLQJ3dOUhBHCVbi67YpvHPk0PsM9p
Jf3Y+8nze9OjARAwhhFdnc3Eu6zMukVDFG95bbudSqFKZa0Yr8kodlWIn1UK3edK+4EJ0xpeZm6F
xqHNZP9kPjY1kZYyU1XGZGbrAlxFXYGOMUYtm+/rbz9h7NlnBaXPoauAd236/cKqaUpk9fhP+Gil
IPPP/xYhg3u2zLoHJJgZItFAV0mtViEbZz286niD/4Vh7WX9VJ4Yjg5a8AgGOLBgJrXx0EiAiMsW
eXn3fxIkw/2YxhvdsLEYWf0wovD4ynMgfuo32jFxUWxRZrJ1Lh/IAzTLTNpCZRzpFU5zbKasWJ+T
Nfl+RBN+zkCDMxTiQT1Ms2TufNY7IQahyIuGfpYdEmBNmxqHmGiGivcZz4zlV3yIR2VXTClAUHa6
0a1IK+cEnxuCqKgJNfaCmVll9AWn6ruzp4bap/sblVgPh+gHlaCY5JAKAR/IWUFW43QpiPqrEpQp
zGHapd6kHJI9WgTgpkBGZLEz3I2yGPvFClkXM+iRpV2u6kHX3slTOfJbx6c0r0sa3n3dBlh95jJl
g0bL7gPN18D37UtdUt2+OCWHkxXucZpLZTey/NbkW6IVcsTPdxBi4inclTSMsOVCWH53HubMZ8GB
ahj8aJ00e4mujAxsAKcD0FWlqxKGKbVs/C6IYNE0jNUX5f//Jk7b9WcxuN3+DFNmH/mh6oGbiHuq
XfX59/V09/DJTaaFy2stArDTSjZaseGomVzFAziPyDczw0MIMFUNmbQapp8JEzAqQ8fijYBmMWut
Rgs1hOfhZ0nRfcWEaFt2W8prHrb5l0IiCwYteWyCsZdVslzTcEoMmZwR8JNt+INQxPsYHZ5H2uZU
5/x9dCQdTHOerPo6iUuHTI6Qp6NaujNF5Sxuv2EyMDpVrcucacvILJPzvsqTxXxBnChLKMV00bDa
+Gl7rv1NoP5VRNDp8rrBiom/5ZDgDvJq1fn+uKDFf2NGLn05K0rnBbkXXRMbOs7ltRWdpoQV1ia0
YUYgk6pmcOqk1iMTi27eSeKzptzkcq8NJAZx57WnLU2cxxLtHmQZ8Es4sSwBU4ApBddPAVDBp6jl
d1gAkXNzhzmyO0rhmgljWS+52krHOU8wLClO8hdJ41lyn8E38iOP9HqeqIqWH1FeSBoP7tBDpGKp
rbiNuE4AMwXMEwAgoIiz6BHPHNXK4RMDIYgqyk34dJdPYAnZkSd14qK4qdVbRdpJPl4WSFDgPKoE
om1uFGahYlSNfs8j228jxe5IaCxeuenEjNJzlOWCxS9Qjhoq6C5KK4PIPBihrKIT4C6+2HcWxrBr
hrW7B08UFIv9bO2XbFQc0r2T1bFruSFSjbyRPmRs1nMso1r1AdMhs1mLRO2kbMgZP8H1z4NW04tq
nklGUZdXK99p6KdCny/qZ3QVfkHPqFmltxsmfeJQvuTLt0EMJN6MAwbr311+5yXa5eUO9QynqmXj
TpZzOnpoYU+ut7rbB65vCtKlPhvBCN337EJwr/Fc5V6imbqvXZSr0oWipVcDU5qslYscKwQA1CN0
CBPOFBZo0gKzXvf0VCKvvu/3L40Rr8920pzvRUTqy7xsnRYnRLbIilF9zn8StLipbJvxM4iOzHF+
ahr78n73IkcHg8hMHO/ppbvkpV8yiNwBqHXmTaLGq85r6rUu+WrC3IV8jaV1B4TWmmU9HNYKHK61
uy1U4DI6NCvPL+btUqR9HO0BXe2hcHMw/6q+DS/1LroYev8VxOTUCc8wjI4ukZcKv/6NnnNv12u9
fQji6DNYF6yjpMuELb5MeXWN2DpZ5tUW8Sd8m/I4SrJdBslANpn3/gyQWU52cHDC55Q5u0kDs/sE
MYTm0Y/TSNsUou4c4ymcRhnQk4d3B3rp7HZVTBLrJ5rdBvOFcR7XQjnX4yyKi+8cNKKN3VW2a7tl
SU/Dluii23pOUtCcOQpewaKRRvc2Qr8qbtPWCL6/kvn6uaTtsJOwd4XPguYU6Hwmr7uEv+pPqB6/
bBNB7ijbcyxqtB2/QR51ZJ2lWa/hz2gU2KobuZ6zxW/yw3brujhRT7Db9kZdPRHa24AkQqI7Qhv8
jF/k8n/ZBPYjkKQa2B5vWdnSRGa6SHk9P7BjfGkKpP09XAHzS4vby3QgDFjro2cevBTw4Rm+MDf8
qB+lLxspz5+RguWLCkbRl8DrOsycU9YNBaZLWlezmz1hJ5hrBKQTo0dboxpc9F3p4Y1GlULDMdcd
QOCPMucVHQ/ymwPK6hoqVmIXfzolT8Uy+yg4wWmOCVFTwB3Fm8cil9NoeDbosmOEU82ShPt5cVQG
4KiWYiLmFsblus0Jb5YEKASOp6m0CgztQwRGMrph6TAKtqs6NMJUeUblFfVGnUCHYY1CxHNVOOLR
ucUrxi+HB37SvuXNoPzZ9AgQ1quJ1RKWajbjzpI9epiByFbaolz1Xf0/0ICvT9uIX3kBZoMZqTiO
86FmhV076Axe1XMPZ6QCyfxjeYql9R6oL+TIcSiX7u8TGK1pVDzYZkZQJEyATusDoKtJjYkXSNfS
1ylL6BXjnuE3hd32s43dusXznMSyoqglfq3LT1k0+hyOoDTz9VNzG8AW2UvgBFfFzrZ+Ukw7XTiD
bP/LuFS3546/Yt44OMQUdLS5MBDCCAaDthVtSBwm+rxAYXe7I+L0mz29qUHCm8fDMELb8X4z+tU6
Imp5SJ+Ov74I0KA6QNp9uHuA2QoIOKZIQhiir2uaa3984yPKVQHNwOrqZD9FSS8DLCYQ5GxSS9Sn
TuhNNfAO0PpzrBYqlzjdWfNzBjC7aiRgj88+kK8+UpbYPfbC4ohK2H0Z9tX6aD7HCEMbcjTRpXdv
jg5AixVb+TtdSIMp3t5C/wYyo9B7/FYuNYFO/9t4QYrk7vO1yDM8yhfZzZSHI23lDnlZbDEpxaGo
C3GLcZuT1H4M9gJcvBX8QYMEu5PEew3hEwyGs2xnNAKrEhW+ieN0S6/5GFWk6zA0uuAvXW3G/qqT
TcH+wP9Fa7NviagIb9HNNcEN0lq/GskyGIuQMVlPI1sUffJuR30FTQxw9OdNHmJeHhKxrpzMGP6U
idtDhWmlYKATiCtwFFnwjvi/pqhG5vys3B8MhmJBu5jnhTXKxioAfF1uhAQ2MfXCUKlYNAXkqjOH
amy9Usi8fhNr/CVlygabSF042HR+6DvySqojAv9sAwh4LUC9xOQMJr1N/NiEuy+XXfkS8K/1WxRq
UeNe3/pZyGLshmp4cnK34/xhMWHqR6PE19eRN2nOoOB5VMZU+DEOkDJGf1978it7HPwIyOwvnDLT
EenAtY4hmwerzlqJclRve83FOUyykmG+b3YVxlUhucl4urTxCwBMJ/r7b87ah+iPJhHuc+DY15PK
DXA3nhYy20tR3YffYTkNJYVMojBL97bMm6VUZiCsUaXr0clVMiwkt1poVLnUpmSCLLQ601MT1ldA
Qn1UlnMgAPbUCbWLdjF1tCaPlgfF5Lo2FOJ35lF5vdACSzgb5nZcaVKDaN6DaHkbp1PEXA4fVC8+
xIRPGIXm82o76iVw851hGpc0bU3GHk9RMsA/Fe3c0jZaSd5gEYicc2u0qrKeFWoUEOXMKMHLhREi
yxka25Eb5E4P1BhIjv0wAjcs1NR0HznSNL0FPn6TlTG9dnCXjYA36/j2vAcSUYSJG6T+flDjsILi
Iv+Lp7zt4KofWLqH4NlHP0uXqs76Ry6VKpNaLvjet/lgBGDE9ZTK2hqysHi7DdWru+SBXfKiy81A
1RxoRGT1sjhJfPi88u/t+sgCxWvwZ4vhSQwy37dwvrmyAStMG4uvNeAGseUhlGyThCJm1o2hR4YQ
bjoGHgl6x8JBwICDh6/FCSInkAQ3BBecRvQbEXLqLSHRaLKBKFxe7c1/HVhPuPglTJbic+h4CsWR
Y7JVWFmLy8SqvVL9iVczW0lchfEz8n6hgvZZcuLV49M5PscBNfuBnTlGqAWqLQa/etScTfLuk1XB
opBEX6CdcTnT7osr9DvNIvfFTNXPC1oJaTWb4pxaR70IDUh9qsC3DneQ6RoRpOAQcFcw97Pzc58R
jKhZSc2N/tw7Xv4C3odlKvuSsOJ9Ofdia2Zi3zzt2wWA2APQqOHNFdGUQFtUB7lSHUkxf6/5XWK9
SiPWMBH/LAzGN8jxd/vASHgY+31OPXg5iT0cZeNxWKZjLzbxDlphIBgo8EADgF/36BdlIZQnnHcO
Ky3+nhAPX4hYFwqF28oth/4OHAi23qeer6NxRoz8AUnDhyeIaBDR3GCrH7yGc+zpg9/OuFTZhCQm
Qr9Kjtoy8vh0SEQ7+S+82ZyYGnmoy0377LxUYl4euF70PhaB+3H+UslLCS/2lxsWMhETTDS+8pJF
ZrlRFuwfbJEvEyWmCLen/+6oHOdIISsMw2t/S/Ql5C3UoUf6HUTnjvLY5qekBXRZIUdGOhYRYSUY
MHvGOs8GEGPhyqlQKfosu6BrzTXl8WzGwt7jPAqEsYVHdNMiNnjLrf3fas3jWoc8MbSpy3Np8IY0
ge3YVfO5LoJEL2nUhjAfMnaSu3JO4sxV/k9VtTRhlkCia4tQz7LgEJ5r/AqD/sKFRqKw1MJOnvaR
1J8WLOhkxXjPqycTdV6Rz+Rx30tOSuJSKLEzh8VbUDXE9kVqwrHkikfAd59/Nybz0e2OnnfwGELF
dM2LVtOjeZsxEtweC7PPNFUKsHTL49zRpDAhymLbiqDlv9bJjjGgy/pJY4SXlI1mmWMYUcuX1DGF
dDvsTIbdwQYFK91jaIBbSpH2IaJuWlsPzbMChVhN5x6vuobD0ryoztwjkN8LGQiNjKmqrQe57141
YWQ238TQp3ytmBhMEYItC2DFDkbgYePNTmwD/6j63dvJVoxnFzPkn8dTBatAjWmLhgor29b1L5Fv
y2ayNYFw84QohrIUMPYVlMP3gIVVreF3Kee5af8b3Sgp9wmi1k/32s2PEazCEiYG/lk4zdxAOVbj
BjVPXHj+QbFCl5kg6b+YTSGXoH9p+4Pre+OgLZr9gcLb1fJbE8IXO4H95yx73Xmv7wZT7k5YkTGF
j9dmjcWraXu33R/1JD+n6mo3J+uwwRJclTCCMIM3ikwrEiLaZYc6b5hzzENnU/iywdOMJmjXANqt
iXDEhIjq1ihdJ9AyMO/GM6Ppn5wtna/Bkh3FE+mwBj9/Vj4ixtqZusp3y5LKH7oCoFw3wSxCOaut
D5YdY0jRPBu9ahwZbH811iR7E7kuRnyWjqvIrTaonJ5TomA5HVVgWO5Q4OEz1LQUSLs7ClfSk86j
TDgXGiTtttccEIL/jBKa5bBaQJJMCL/8Ro4mI9FrmPC/y0zgpAaNxjPAszv2OtxPS9bEj22UIwL/
YHVQ5r/u/K0Slkgaym9rRrpccnmWLgR+abjzTkvVJDqCAM/5/QI6bO4DtBgSqTANSh4oVu4H7m5T
uAgrXuBfmgeMMDYfpZ+pCH9vg4vdd/Sg2QGgSvpZSu73aiPQfrTwGgqppmQ4cvjAJRmGWpSGCpWk
sHAumcNIhZQRvd/06K7CBgFmCq1TaqsLpeKvdRxqhvL5gNW+7HZV5SoAUWVemie+OM6tBGx53EKn
DMssnXvNUphLYxx/WByQFgtCEIvIav3L+Itk4AyuU2seQIFod1Th+n2QNeal//ezd0wFuaHdr9BO
KEInNFtLVDBQLarvztONIKolsQGoSQ5CLx3cKevvo4Z/pBuU1UzQomvjJDlq548RNCwqCAnGLVf7
eP/EwdOUNJetVgaIGpKgfcvuXCuytNS4AAExlfhslFBvFY9uwJ5EUIVQ8iP2K0pEJPHbCRYrddXW
lN85rIgzURd8/YZ4Ej5MOlGei2YCFG1JJIKgJnKxKPNzAheYHXJcOU4IIqA/FqVCjM0O+ti9ATXq
OHR8nUKAZllRHqMMlVzAF02O4g55f3wr1sL8QZRLdu/f2MBmVaSeffymlMWQeCbHzb9GqHN21q06
n/bOY+RHQJSHNOEbsNlYNG9g4m0mLy/zSU+EEWqIPLpDsUyNqzZJdpMd802Nz4FnmgQhoGUYP6nB
pnHwyC9lg3pAWOjVLdL2cW0nQV8IjyFPIuXy0djoMiiFaElq9eNlHezLlbaFDjvyLHGNKMpJkhTs
+60W8zsSg1oLdAURQmUlwVl+hSnjMmgqsTkYvyk1JuTM7wqAZ8u6bWeOQC/wGj3HO2DcGIjhn9QF
8S0jzWSZjRaG9eEH43iQ5fuZMvDtXDACEfhT8bgfAu9ln6gP4dCioxj9Wrli78P1rczJL+l1sX5+
d2l5ZfUG9Oyyk0cNKAej59RDNPh16kebUhYj3fV9XcTHiC9mDEUbk+M+RSZz1PkXLXQzGD/s3V8T
WH5CAjfPdQ8DpYxStvpIjwSmUBujoIeBf6pTccAFa5tIbVtzIShmiRId7IF4vVnLDsG1yumhntxQ
vyOebjxKQl93QLg0pDNkvckpY5mah/GEKbLLmgvU1CXHyKAYut18lQbDs1krsZpOk0ZHFaARMTcc
l6QrBb1ACSqSUUBm7JcVNg1sa9kvGLL3z+JeeTkW3BzymXlIKjeTS8b20A8pUDm5N5X3UvtxZ6uJ
FVUaCErUtzMM9ZIPaaFtkVQPCrS0Bv8dC0dncNKh5g+An/ZtP47+ObS74MgIkUj2L6+VgIBhmYp9
wyInx1Bzf7OhW8KnOKRTTHcTqBWNWRXVQKu58v0fhNrtrUCPbD+MbLU8OwSRQqQg9ybkgc2bkxb1
QuajFKPVeUa+71gui2dOqfvwgj8PyLv0X3aTi/ttqCBVTrV879JFgYEGpA0WjElmdJ/jov6umJ4a
rcP0v6KfTgh29ddymPlHTNYEsjW811ahnFASnmxHkpfxFc7vukDlaA5eeTQbC0TD4e12JMZfvbmA
d9XoVb3FedBLD33dRGX6iHVswnvnuTgIfFpC0TwEF8iyU8mRvJFCxVGwKdCJHRYGpcsF9ee1waoj
YpttQc3i2Gb+lVn93pgyFdg+f+6qKESe4Jyw1b18udpPa/WtKcqETyenBw94iHaZjr7+On4k6U4G
nhqPIRGBuZcAptNILlHTMA8+/1HDqH2KYLPg85iZltZIrv32LPZkGI4Ylajpa5vXmS7mimjvoDbR
n1rT/rnVftSa5halh3ZXkvlNAuOwupy1duZN/7T5yzhNlTkI/tpC80glyIVjnznrp3EL7hO3BRVw
7tidOaa7MsFLi1OJ5uj8i6sA2Dn19Rabjd9zuHWLY/OZpMUq2XsU3A1Ah2Hoi8ZmIetuv96w0pEy
JqW0QoFYQTGdVyuXvllDVT3ep4X/Ird+OaeCN2gwI9zbSvNkzcX4BHnMarh3lJ4leVdti2VMt2pC
BacZmtZQDff+ZCCrIvOyjjMk3docGUxFJ29DKmn4tALui9K2Q22clnI8NqXJdEBUh8u8B8mfNcvd
f1hIKjQ/bHHtBvt6Bg0DN3SrrjSg8//ric8woTQCMpbrgVz8HwOPQtfPPRDYExSf0OWpXqorlboC
hIpTIOTnSrKGqWm2Xkj4IrMOPkY9dszVZOhz7G4bRzc5EXVew+5QitGWtX7Mueptgemohh4jRwyY
Du9Hd0oSQf95wlLuke9L+57jlaUBrFDFyWJqVn1rg00Trzzyog+nVpT9EiHVJY4T70r30/3xSNyd
2ZL9pTzvoh8p1GZdfmgiCLgpS6gvLQ84QCHHnUqsezzyE3PNPvF6aM9ypxhf+eZteshl4HmMfpR5
LtTxRdd9wNNxNhpeCDQ3TvqfPWjxHeO7IpmpqVmHVGy65xME0ejf6IueZeGk7+Df0KBSgWgxIqpy
kAHvEcJNP7Mht0ArQsldJEwh3z6XrLW+vokSCZRJbam2y01qHqqk/XVkIzGvB0x8DorWX8NdnC5S
7+tM2Dif38w5JRzlXj5YYcP+9XoSNokgq0EKgP/v1wH6WypaAkkxOwsMs0t2m/LTXr7gqpOLqVbt
ooyqmMO6wSIpz0O2MUpdjl8YGdZpOACaoEaI0m8e77uhvj3mPuwfhZu+9gC6p1pe9v2jwhisH1wo
ogLUjiIscUOkKJRUSR6J/l62pWq5bSjQxiYZ+lzPOtfNBdAIFpH5P4DRQIzAELh+rf+K/wmwSNTr
0W5eUKveg8eNttaFJOtYeGYK5eVYqcbRPWsekYCxUJ+0UME52wF17gi8/wX56qB7BfwT6XYHQCmR
uNSgc0d3SFvAqmvuQMoprNWMoTWV55TyT9uKDQg72uzENnCGrOfhpJ5Wy+ZzUXkY7mBmKBcKo2i2
u6BCmsb82lvdoUdwMehIKxCJn8nke0cYcYSYokErF5mxP6+7g4+8hnO97QsuPFEfhnrl6NKyvftx
ve8kd4sZOTOTUfr5zcnSthvKgmsd9mNu3ARwBTgMNi7JFaJH2AVROOuQJdr3W7+t4opUcFCpmgbd
KI/hJrkN+yx7PEGyYhWiO3mLlA7d/4aE8aXDn13tQMmPJtjSVOak2DKdf8zIv751WCATakRITW21
2n2Dh4knVuHBkYvdenjdO9VDRAewvOmnWm4oiqU40JrNas5t674jxs73xicTb75AMk5E3GEX2U45
eGleeyVadBpxadk5+5Jk5tVOPGLxXml4kso5QujbaLX5spNlUGKxURxniQUwXHgKV4pPV8HcMYdZ
KCDPoUXOjOTy1jWi3EElsAF+Z65+uNUyKUet9fKr3k60MAWqLQN24mzRGYr3N9hpRs6bg3zC3ryx
OsLyDDaTUy8Fl8ShivrLwfYzoMU0xLX4yCc+P+ALUimqbOoKnDrUY4JSU5RRBGl3kOtdYr/WbJ16
aEyOb5N/8UqQu9ZkF+/PxWdmBQsPx1kVucZQYFd+PMWO5qAUQvsWuZ6dO3Snz1C8dcdmr9/Jxb7L
OM9T92uIdjfWqtKtBIT1NuDAGCVqHCREmoNXHSGwJ0HVEPS2Xue4/EYWMLXWIPV6hmsSrsvZw8rk
7Sc4ZAFL93HDfgWoSheh6frnNDAzKTkAGMUrxxDssK9QoTIZBY9yswsYyeoJcpG4jWPWsacUmcoi
zG1gafF7KJbpRU6L8wKKGa1wTJAlCQyi0Iqi8/lg/0g//cPFawzoUzVQ10hjGhkp3Pr/R1ZVMod/
idJK/AJe0V+cP/y0RGC27Wks0Cb2VvnxR7jlvkOkc+fpaygZXABhO/AKRIE+D+DjZAJpyPntYKil
yTe2nlROLBJEmK3mcoZAdpDtipImjP3hwmMakEONLSgmhOPZT5tix0tunMHq6XUGW6j0T2bIMwOj
78WwyLNvTyWdVOSv5j2rOBLdJlfUmQEEvumKx737UYTDFtcqwdZ4Q1LP71VlhFbnu3W0epydHqD/
y7KGq69H+KQgmgp9H1adTFGWNlV3JeNRCHa/VG+ayCLmC6U1on0nYK5EDIvNmGzzjY0lKIyR6nEL
6sRyw7CBHie69279Jj9NdJq+bZEE+IE1uG87Sk1fteZRRbth1+Er/+5q7D782HQjXB27BbFtFc8/
2mVwFTvufu2Mes8g0xT1WxU1PxfZfe9Psj3ODhMI8YK0q97xJoOy6Pi07DHNa3CJ/ZHNo80LZuJ6
wgHKvQj5FTKliLEhnjRWQzI9ELKpwKVRhGyXtQ7oleGjCI/aB6XTlRcu+xSQByrEp1oKRCES4Qiy
C64B1da20unjTplhRUTL5RXQ0TLURW78xWH3nGRrkxGPKfwQ1Mm0+iyYYIxd+7Y2LlP838cSP3A0
9/47wYkT8m829eGosDIiXLNXityoaoPcftSMJhT4ChQ5Fltzk3Y+BojVgtIUf6yYxOG2i5voh4yA
CCqoYOSfrXN4O3tj9TQMW9lHyQZagyGwWx4rUr+0AZJYvRvXX4ywMdZfbVvzTAT3CC0T4ZS8SdvM
3+/Rm+YrMFwmmTYnZBa2PvgWvvIXM5QLS7K7K5r5kyV5ZnRVFg2TbAqZ3d3FwAyC10luAZtlMgAh
6WAvmzM2sTK9bYxs5SSeA4HdIG6d4IORqNbU8mLhjfSZab3806Rikj6qF+lTW6QOGpHmKlb2b5My
I4hKJ8TJbKmscHLxM4YRaVDacggatqSvIB3M0ptc2VSJfXOTvY7pgQ7JXuZ4rFQyacakRgIx+be4
GJUQycrcgqg4tBWsFXyT3KxMbLPZMb30a78Awp1sBpGdT3FRU7evQOsxt7gqo0Y6nN8DgotzPwvj
sHxZ82bLqhEBEXPlJY6Bc/p0EZxshsVEalvfLzN7rNOLfsYjfp6u9TneSauYH/dyjwXHd2KT+0Oy
VfXTZEH1hywtlFS2bqmSXUEAQZ1UN5g3HG8O2NcoUH2gdkL472/GMyq4NwVUTgweQS4lG0ToLxhq
0gOd6odc5lhqx6r+Owby6BOCKgoBmEpSdEKJn2Lbp5/VwURJIc9XRNKZfMIzczm0e+Q2sFQkCk11
ixJGzkk43TSVPdRZBEUbWB50XK8vw6vRpy4Awq3fPoGbwyemh23q1mDI3Jw8g+KVKGHWgJfJniAv
FL3EarRkCPiTHucrhFc3yRqxEUwUD6CSGQIG+THRZ+46fuDSd5XIbLGJlRZXVP3WbTIj9Iyb4HiN
RfXCSj7oOTGvct618uNu8hFGJbZ8+C8mcc18na/Eh0Ix+MN56O+D8auQhheCDgAREz3FguWeV+7a
UANhjsiqy9TcYEdehMEoW9IlMdV1SEhSa/mLeg94GX7nmd7gHSkVZZe8yT/nNdwbE7dHXkY6ZJN2
IIfgxg5y0IsQTC26Yv4zdMySl3+xy3aF3hgboEE3alQJr1gHy0iOPMlNZVVeoigEDF8e1V9nv4lA
6iXijIdxh5HdM2mpNtClDYkxBveDcAbfNnN3KlMaJGWreWY++yfKEEIUrKb/j3q/X88PqHSghmEb
MGDTrrVciaBFiAU1sSXMqb2TZWOsMB/6606hFWguR0gekVxAJF1S925GT3MpuDlvECU4383A7VHy
8SR8M8Zf6ns26AgH8YWx0BxotCFR32LGvfgw4Kt2pTpoZFLmb+1s4CHlombKYWIzB95f2nTAIQx0
B4ggMF/TWl32ml8wOShpam6szJK2JmyXQW5ZjxmkYkdtfbTS7r+n7RTTlw6hc5Nz6q1BmI74Cwb7
Q1bvWkpxFAjvAB/6VpUULMrk65YLJsCltv5DrayqiSp6XA/AA/waC0plneUL7QozuNKRVkCrw9J8
33BpuuYE6MQThXKK+amhnzkP1gAg0RaXJ1qp0aqZcNSW6pLLD6wkwO1eOLjvA988MKY63ABMFnAA
6FtqPqyPl2DUXHQMMYUWbg8HCAXuGVeFHHaLzP6bwAnTC16/zGrtpq7+Fe+SH75e8tRrpn5pSRmB
6RJd/3NPxuzFE/rkqwgtoga76xa6pbmH0tAfRbJom9YWdTvbNnmuUfSPNGucATPqNfk9vlLlHePO
RMBzrIFSh4rHnlxAXBbNEkTBpb27L5XDA3UEcqLSI+VENJPjQ+u3tKocSxtrdaz42c/ZobQ3/w2o
2jbQP++FNwlalz7NTOKfVjKNTO1xsQtVmNwaL+Tt2c+QaYFBNVcChIED1HnUfmdsbhjhl0SyWVDg
7cLJ564npE/e21jVN7DscO4IdNUueDp2A7SLxgPalqGUWhIVM9Oq/xuUZszEfiIqOvRumAiR3Nof
LcU1tJmKqlQABWItgyoJiNXjCPbAazEcunPcyzvWJAFMvEXmySqnig4oIYpPgHP+CLI8dxOubKX9
mKs9SdInr9adG/U4I+rIcgF3ZQBIIz+9v9DbQVGGjQT9dKJAfXfyD9ioQEztxrOdEKPcFf3Xqbim
l2P3QaK33qgZOE3dmdA6rvmvIdg5f8caBn1kAc1kLeTtdLbC+i+pBDgZZjJXpG6h4yy0IzoINPQg
wn8GgHDOItQoDleD+pZcruCfskJN8sQcMG6L1x86jTxnOZ2kpnkUV/pHeqdjF9IVqfYT4J2rwWiH
MH0kvPeBP0Ej3M/bJI3rus77HAI6r32zOCY8c2KRNe6YiqFtx4A6xgz7764D5XIJR+hy7WWtSw9u
9ihyEakraYmIusY2LymmNNe7oZKw7XbpzjRhSIJnBOOC7SYLeIOOcBiZW+TJAvhzLD0LGm4m+hlf
IBrQzM3rTc7ylDX+AomqQ3umCSRwDflNwTlZ+J7hzBX8Q01DAHQMUUE3oaxO+sr5VY+aMNWoYNkg
7t8/gXbu70/Grtgp/JTrinY/gVYGA+/g94SPJshEWyPMGcJY5pg0+Cc9HLg/jmGdd5uvc1e8iQc4
kCy7O3zTW7+yzqwhOdD/a9oeCvB0Osou36Gyw90ibw1+gvcvIN2TLabgvrTuKx/NsXdboR7V2QbZ
MKDqLRRlqinBAxuHxr864y5DSpX767/7MkMIXo8TKzvQjWeLofp7N5LSgPOR7ahEhdXuBEXKL+bW
qpBYb1+B6ayPTuu68/tG2raBgxPzgJZcymHV3rsE1dOT221pStf//eLTriWCGtIxR447SVcJiRTy
RJUnsXgAjSqWaWDUqTsMau3bsbTCcpJYwnYR5+Khg6qJBPvCK77DR4PU1yyu23+ado8kl0Fo0mgF
vPAvdxI09BbfjxWRxUOvA2j5BDEKwh9vj4zyN/GzawJqe3VpZnElN8jA44dpkkceW9Ejt3itPCdZ
QrB2vIvr9igTJEAAi1euWB5wDKsLZgZPsxfQ53i4kzmE264XkuOsIKAuvinyYm2ATaiScRbtfJLo
HX1GfMFibZSPMy3i2zPOCV4GOzt5REin1QwuwApRkNuV/g7y3SAx+vWwCqi4dU+M9x6YPsSncG97
TIug3lre72iNr6PlTvIoENjnowLppGeNLvLV0ww1L0gd4EZH0l2QH8zci/+QF/3VA30bUolGXWJX
aTwtwrxHhdiMI31G72zWoYNub26OoPFneLkmI+DAck/fH9pB5nQkzrz8sIxk+D5YkPTkGls1KnJw
mbyAgCLsVMMNp6JMke44ODT1xhg0Wr3T/ZcR2Z7vlCjDh9jV06rhFltHsT+72SXcTbZ6mN9Jm2lO
W8BOxiinm5cUPzzwd05MkNQ1Vl9oxYbPFHq9m8EA7htGcEYeZ0GTZAf6bWMRMz6/L3jyleEYZXBi
GuxBoE5zFf6DiFrOdOgrLMv2v0mP3+cJvWQIKso0rrgnVOVJIZISrOfTFNaD2XZ+kAMbM9KfFWx2
LJEudjZKOnevN8JNvKYYBUhBx5TcCihudL724A5bWekzDnSc0+hQEjKCwrMjc3yvY0ePMpVDeatu
OELmKFAtwYytEMgP8Cor1ehPgD6ucjlmV7hGFNGpiVqOr04PrvX4tqdfuOg+fmgTFqj9ClqZ6gTy
VmykYlwWmGc9v5CoAW2voFw1ERS5EqHviZTnBXlW45sFFopoBqFHYUZu6wbO8ke+P2e2zK77QbBc
Os/EoH4TPv85u7pDdICkN2yIhuYXpyEzvCPiF0QZp6RwbijsTG8FzPPrxRfIVvfK2C8INrQfiNFM
/xdQhZnPhgVh/bNr8pWWlDoPnJBLb7cmBkT7Kq++YneOH4vk5lJxQOS03ArqjDpHaIPOQzIeiFZn
qsFEHyxi6tS8PaKQ4ZVypr3IsegylHCz+0uM/lUQCmeCovCxWD0Q5IMk45xPKwyzVP/MZuGqTuuQ
KKq4wsxkbH+69GC2FG8j3bxnMu3C/KOk0wnqQck4wNDydoxjV5JAt3CFBa4k3Vs/MT+3zrLaBrvW
lkjlLexj1NyAhPmKz+wBVOD2EtvcBsbAL35fMhWBRGibLJU7HY4CqY1LOLSo4vcG8xzHMfTThBzk
j1xF0MfAY1LwZndN2w4NGSNO4l5Y04R01/2MkNo9IkBiI1giMzFGkufLmwEmfMDwUnY5KQaKO8OH
/1Ax8UlYAooMEBm3acjPRMKl0DdMt7z2ZP6POviY3I9n4tAFRjTidFxDSvAjseIUUDXSm1wpjksR
xENjc20S2oerxyijXI1tII9/fIIVgyBnvXlUr1f6FjgErF6A/GjDIyaR98tOXofazr6grSI7cEKP
h0GQXXwiXMb3iV8m8h1NA9LOJj7AHuvz7Tyz4xEnIE0c/UkLAeM7akGrs7EThqDi9OLxnGWt/ESl
RRPKb4dWA3I2dkSLlrFaJukIShurSkY6LTsXZL5vp7YVuw0QwNpDYGvT4A7LBqFGGpf+OMNA0R8F
ZRwNBwq/7Y/Iq+sSAH1V38rttXZSkNSrI2/t40h5Q8etk4q4FNWn6pL67c34Ts6d9h9MWp51/fJX
A0BNopptv1FOCQssAldOkZxWe/nvdy+fWclHC9SAXfFuIRm2VbvCHauhqqn6duP5WX4y5Q4Eide8
fWK8c1b5T4fMz0yNacYt7kEC7zVH5UN/uhKM6FO4Pb1jPQCJAdeTMVNSoeH7ifjowCbxYh9mPrgz
oenCQjvQACz8/taGt2B/UOEXovVBpZ4AnynpYGWfKrjuXQOInB5N6Wp0GQP/5Il6ijya81q8+PRv
Mc/ckJZ01RzEyIDwjB9R1kU3DziNpp+ZTp+Oywr+dirHo5V3n7e9HeHXVRJji6d8ZWE9etZ6+V5R
fD9TSBWcZaahnBK02nAJ2djPQjAy6B8g/74lTE7l+8t9tTLZe6iim6qXd0nH0onIjnEq3egOagZw
9ezYdo4lD2f+PaTtQnrVPAse06Tb6lXT82jvOvApHUbZqSHMHPtXlyeEoIMHkGEMu/zDsv9lorFD
FEs2jFK6V50VARBeTTNh91Wr3WyOrRr7xlByQFaanzrT5iG0jM9XrsF7sp+TDADRxHbdk2c2NzdX
q/sXzzcOgl+3TSYX2o35Sjvs3vRIhcsx7v9Ztdft/aGYkhq+Kw5SHcJ9OdkJKXcWrSTjpd/88q2h
A83L5N9SPmsUzPd7b4GURO+UkTXaK8TSc7dq+r+ranve79eJU43sbuPo34pICWGhaUXlLvnh6B+F
OjuarnLiEf4YSPL5I2mKmSGtBMVkprFnVPzpUquvpxAsh+HNQ/De8xZfplUuXFC/w3LqXEz3FWcx
F9r/01Ni810BuOPqd1P+XzQrx9j7EgmLWc2FDVqgC9CZHhhqdN4M+3ppa52n5QX/Fx/AR8LSSs0Q
8odrmg0kmxgsfDXEqaMIpvCHycoAgyeOxGen95pKNMol5a1+mqL4yc/UmPyoSilb1lmkB6eLBtQE
1w0Hm2BXLdY8QOwJ6UDe6ZetgMQbXBn/ep5fBRXnd5VimaibcqCa8volpvNTsaBPQZwoYQ9CgkP3
rwHxEFksEtmTE0fUX6ScARxaRrN/yPjhH3akXS2/QLr09zXvtXePbTKrfaPGHzHJJDKUhzOqwNaI
DEvO7QvDPz8v7g+CrhCr0YOBNUJaLQFFdhLIuspdafpyJooNgkGLnTB1JwFraCX502o+off3UFHA
FE0uuN9/lHSUPIF3AYPbd4EhB+U5irmu8Pu1LSQJKzClVrEs9jwzxHggMSNcYrE+y+r/wlVMTXgi
8HUiJry8dG922Fubn1MfHnSLJmdiU3cnh2374v2xdyW1DpclaHC7gZU3aAgzSyDhKGtYa/QDocoG
seVsmfPpyTGXA3ZGCP6WLZvUceI2RHGnQqitCXHnps/+PN1U66CEESLlV9HwE+JNa1mQ+b3b/u03
jE7kc98veKQkHrwSViimgh3cmvm8/8pnbunvwFeVvtWvwF0zrFKx/INPPHEpxwjLfbNalWymFGdu
y1TSvhvk/gsgG7RgCQolQvkauJNLFX/QpSKIrRsw2o25zhXg/UvnSI3AJ6/6YDruTEchs43EoGF2
LW/bHj0kUZDG6IhekVEtZbjJDcKUU1yDe5cLcgyjSQfCdCqpHntIGxk8/RkzURrzPTaYMqCwIHTI
OzjiaTezpbg8BrGvF4Nuk/viJ3rxfKWn9vuVnd93cA8s8iPHo8VJb0lWSHaholZCBeoDs1wwUgHA
lwTHlLt51llnFLdeL4OZRytvjT4+Q11HqSpV4YvOc4VfZHoY7Lf1cW2JCYx8gt9+fvrypa13xLNc
v0MdIOIlsr/3Elr3oZTDr0qYvulh7hNOYUeUC9cuA1ZQDYmh6TnzotGaiR4maJx8GtNTe4xZ/bDW
OgLMTH1jA1BPFKSTn7qn2xDkBwTPAddKoURYpiTZvkCk2ehIINRPEgrI82nBEVsx/pZhUak1bEYs
rswiCrqvXvKO2wR9wZxlNHsw2seV9s1cV9GQCe+/JgpCR+kj8FaoR2L9nHthg7AKD511YbLMV1zV
xW4t+slj4O1sA/ktFUMVy/Ur+ooeDOh9eV4X55zQ8q/KfBy7ekE1RgO0wFJ/QBz2U07JlFrY30IH
s9oeLyMjAataZXOhKxK8HsmxvbYT4GnUFruyoc98ptf0aDO4dMX+EDKtgDD7qZYUGtTUCQeL0KL6
KJEb5837kNqb+UP6T3dfPsdyWJ1MQT1GX3f7FuqHDIShWstLNlt3znQrc18sT4Vc+3g2NA1Afywb
iPwYvDG6HCSvlytCQx3PGF8aK5JsugbO8CY+G0RdyT75U99Nc7Qa+71OnMJww3kzgqOHpxjiCPBn
wLC09DI1xaxWehQtRasLZ+3uq4NNSoNtE7rxLaZmKmsrsd0x+gOV0mzR+FU8ifvFbGeSfNsaNlje
iBqpBVLxERKZbKxqZeLD4AJ6FmGwQDwjxhd8oYKkf8DxP3pIo6qyiC+VMP0kurA9po5wJCtIbHIM
W0KzkDeZndGEs1L33mPMYwa0x4i0K/9M7feg3jAqdPkElAB+CcpJvMPX+Om1bON2fniBQBdWCYb6
DZ6sV/TGLGlHmIhC8iIzHREGHLwH5FI/qEZKopFc0MfRPclTa69xYdXbGHCP4oizoXiB9cQzkF9i
4hEPYuKTu1AiPe42ZcgDV/sIE5QAgVs030v4q0UE95Az5iOh0/vcoKQNPSHhm5caS2eqSnZF5CnQ
rz8nRVLUXYaYQtzXUz/q4a1JYdeXdqTAldXWW0y8pEKEzPcRtKbHQPRsJPWI3kAR851DjWaAzp0m
QSD/LbpLVvd4crfu9Eut24vHTuDsJzRO6Tivzi1+FHfI/OLtK8Xvb78OIiZKOy4ZmaBfwnAf9HIh
rpAzJr4w2Zw2JucCrV++3ybhKlN0emdiUf6C7wADHdGihpRppafhFVE4RwH+yB4WcbKeloUV2g5T
uIZiTYoJRKJ7mzlWcg2D1r2V+cUvo4xG2e4yKWuEiybM1xke+iuqReB1YX7i2rdt+NPBNv7jZwxl
oSurKEpE8x36zJ5P2zo19oLq+xc2aENKeTgZs6mz8c3ixtLzlIicnJsWWRiOC2th8VSU7SjSC0Mq
RZedDdW+0uMXJ3T7wO/LfmDJDfIWBfkadqnQ2nl32tf0nErRRimdy70JsiN5gIuckFLfJlXlhOK2
KwiJKa2xvQGBPowC8E4UBvdYV/AnGxvYd5qOtN1mlGU+bkDbZOUF2Eu0ymYIDOWV+u6UPtXk4pX+
kGxqRSIF+hZVS82lAe+0yPzefhduXNOWhA39giOu2ozNm2DOumKEZMa9EitXzOcWRxTcVvUA7asn
ergXR3/15QS7Y1ZONLfOrN1+scSAZEndXhmUDZpaavNXmQRrbIEoVreO/0Zfphys8rHCyczpKQaw
uRP3NPD3GwzU9fTpGT9Uh8wz0S9Hc72oE3RTHf/DDZdMtox3TCIeOT99q18gWETz1BaatJFRGkB7
GexP/RsNgzi1J6iyx+Rhpw0LY29PHM6FwRLKFVg5yTmZbSx3a21VXMNHPBgnLTqICTtprsJRtRzS
E6UOEe3qk3ZvTdvIkskBnj+ZiRWDLT2/xccXN16iuQCyGKD+qaRky8D6KQuUVExLc3fuJcwlZ7AH
h6r91bmVDACUN6J2nV6dIQTJKcEo6NKfyO8e7KJJJG2oo0JQQl5BEFvgkADxURD4Yd4Uy7+Z2yhI
qd/k+qXAYbF0LwimdJAP3KsO01o9zD43qlfTTmZiyNbNp6hbNW8NdxOBNjsEGRNJkwodcQyT2Jtp
nGdCwnzePAJutTnjL5+Q5na1aMzPCfpSSTRaeaLJXmdQ8OAcu1vfS11r6iWQLtD4HeUemKNlXNO3
Y2AX6qUFOWJtr6j04xH5yikcZX0jZtaxsZQ1lHDfyDT+vuij+PNZeg4NbnalRlBLgS56frdTHfxR
ftWcLCg43RjDG3vbYbGieyEnDeTlKOvk5lb5TVxN2/7vbv5aHUWvXP914/IiMN3D9wwXcLE5ZILj
uT7kaG0Mn3o/B6rdlq9VGnVo4Sp0wuEB7+jE0XzenE9zsmhr8+3lkiBcFAqBqJhMBsoUqeTILN3x
CXW5jnulkoJOovTl+mClEoIUm7RaTODo4RjlGoSzB8bYAzOqjtrFkZvxLzi1D0qa9sEmEBrBGCoq
AGoqdE5BBNTxgzhLTZ0nlFXZhWfwl26y/gnveTXmh/NdgTz+xw08jS6YbsgZbA8ML7V9mikC+pti
evcC5mDw73M9J/BVAKjk2Z+fQNB1ielFM3+DSYv76fl08zJyMts05SiehKQkW8kPrfhUDpjOrVcs
s7TxfdVpTjZNOl28RsJGvjag53R2FvzBNYZDlqN8wC0z4CrNxouTemZW4CiHUaTBnQNk8RhO2jF2
R9Okrn9RsOk52+r+3jc2MVAPIx5o52lKpR1C/JMehSFZ9ketvJmdjT7EcMvKdSKNj9NsU/goFDZy
RMBmp1DrxNpX8hdIOMjhm0wxbhukpNGALq3DgQ8WFbCInMuYEAo0QKGwiFXU+RXkj2UyvO6DzV+T
rqhFQvf7jCrkfGLv3wZjQxFfvNzw2dSyk1WhwZIfdPjoIMBIKT1ZMYAwUzUbt+YTeA7tmyE0cdw2
chJe1YjjVdjxU6mMq+2Had8+SvhiVW3M8avdJS5fKQ0WOmgJTPg7S8lvCKfdgtqSiFkNP/ERUQv1
Z3qNgzj1lRtA/6+py9mdnsWAJrntZ/xeylphe2BVrvnd4WbQDH0JAliqwlssluhg1yRYGXuJXqmr
EFbjd65HL+2vFtDvwbGrbYXU/bUjCNp9nf0kHpFH2h2C/lj+tsuQIhRM2i2gy8hPXGmpFBRBiRDa
4p3ojzyJJiXgEsqTNXFEv1+2zhiFssi9hjADi1btrIRcWjHVRnD97B/tjFkw2RQ00l6BPnsA6Jzk
TRzpvBmt4eG/Dqurn1dJ1i6mdiNIfuB3Q0J2CZeqILKI552iqDSxu6L7bKlWg3mZbThz9T3lRroN
O/LsEIOY0OSG5yuOrKuXLFPmG1LPDBXkpLfvzuWUYkOht2i4GRT774bDvLLKu8htsOBR8gubNRUS
OUZ5XDr8afVrgveEoHnmtvfZB2IxMEJKs0OrD8FzFDcGM1l4WfZWub/Ru5n4oit+skxJ3r3mr+di
2TRHsfbIRtuoWnPMsWQR8kRmma2LDMB2wqPg5Ju5R9Ex9NdQrgwJ4Jn+v6SK304WTuofjG15BdG4
YTrgF5/iJiJoTgeTm5Pt5kgcl80ubx7g2kNXQfLrbQ1OyAk9pKQgXfM1tmxqAf824LtWv1dDtLqI
OlplYCnFm8EioT24g9rZRSvGei/eKGyT1RLfAlTbZz5y5EgR6IaVJ/PsnlI76kiEVxHQZmhdckEe
aHRvgdUaOxXl3Xgz0xtjfS9bvAHwcOIxRgH6Dr0e09e5XI5j6qzZEFq/03f4+3iNtNXMND08KViu
kaHaGd3liP39ajduIOfX/iHj4kyVD6Z6q8ee1MAlkYbrJIcKdg6hwhBNFpQVSL8Up4RGTX9uNIPm
GqVb33tK13sLy9oX2XSldvu2nH2i1OSogQ342fvmxQkLaYC8CtH8BEAV6/D1lJD9KpBVSRN/gbHl
TUorb4z3XvW9FR3FGiNo2ZwThgokqcbrqiTmkzXRcIYmQfrSgWdJJEUetdFV0d4gGAEFP+6kmdz/
FsNfgb6Il5LpwC9bN0feKBxXUnDqwu1CDD/OYjLvVwTJS+sNxTPMD7+2GNhSAH5IaqCJ0K7k373r
QIL0io5+KFI8wWQLPpXSUYBlrb747Ie2bdTtSGaIzwbwSw4rOKZT941sYjAzOmfZ3f1l17qdKMOR
XvPJKOSeK8nNmvUJUzS38zAdVtobIx5zqTFHO+xrXaELATF86hYLZRarhizviYoiyYROugxXHgiR
VEPl59zNqcW0qTvmJp7rOCc/EoOiG1my9SgOeGikHigxxKC4gjUZHsl37WeMRTRNfWoferK4XDcg
9AVYGCiTYSjK81Wc01SaCSpS3pcW7WnjCHZFPj8qn8UfPLtBuZMRHvnXreZbTGtma/zUmmEpmo7I
o0T89jAD5/oQiXO4ITdldlWb+0v2CrCp/bcDof1bN3deDgZvtjePOKmTquLjR2/hnEvBKAjO92rB
t7vjRrlJ6cPt2uMHiXfkv9dHM0FjsXMuaJTgx2ba4M/NvBOwZe19YTNyIvwIA1RGogel0ZyazwHE
3tgU62j3cNCLh7Jpb/pBjkiK2AoQrbxWt2xBXAvKa0G6IEUV7DrFNhBmH7v+OPTFkxXJ+4S737Eu
Xa+jQ4ejor6sEVBMAH4XLea7E+W2dL6TphIbhR+fyYXZARXAispICBL/sf/jcee9faUfFB//KW5E
nDhPabKBLryHafiNZ0GqqXeX+6aXpWPZbO8umQmOn0iU5YqADkFfRkCXPBsM0pCeRLCwwbFG95Cu
v8VyX+6dFT6T9OhlwdFZWV7l21XoTQW8HE+2c2+N7C2jfBVfMdIM056G2A028gaI0O2RF/7ilA4a
hygaiOgUeXheba06YkmEw7AjunAtFJ1SKCPArElNedItFIz4juAsJ8GzDsIP62SentPfI9yiFpxN
GT9JBcEa8rCAgEuupq7Yd6QQxIvAh4pZcklPw7e3ciEQJy4oE510W6hlzP4RS1BU+OfHbhrkbw3g
9pj0vMgQdOLAQfU4udaZS1YVova2O2DZcbh+0CPBzjl1KMAqNX48NBHGya38vmSMDhqRZUGFZYIP
ZtLhxxAVNPPIgacr9KEd8fe8Vr/xhzGMd2yjlUB0uNjSHG5BLHTqRLQ5KbA2UrnoqsvQJBOt8JmB
PDSRlklNZ+wyQ1Qa4YhPCZXBO94kUEoE9hmjDKmtFhcy0AORapGUlGMfqeJ/9JBMsVMHfxVWDI0y
SeTPPhZAkoVb9Nb7TfDQij8Fyl4jfVFMUJ1xbdCoGZ2z7zITi51HknX5xd2XE4+AXU3mzVVMgNva
KPthnearbDvdVUv/BCqIyTbIQJUk4gi1owesxw2UGgTGqDl8PS1PtKMlhOZrTOnjsIJPp627kgBJ
Dkh+Wb2nw5NoM4GloJGPMp4q6r/Dns4F/JEwtoErPkH4I9gr9vcEc69q8BNS1vbzBOuxj4N/NOmR
aAjQWxIZVE8ukrFtIHviQG+Po5543QoUzYLNV47j7RDC1ULeiLEoMzoGkdvyJzyubjS+H1nPte17
yCxFDYGazxQrhi/WOsismhGmBl8/pxVCLWV2bdE1L3E5j7kYieyJh1KY4W0TT3dpOwy41EXpUUql
SekI3eh+3KT7jmwQeRx5df0Nyb1kMwjSOdLCJElHegaC4O8XmgJX0pWX2aDPZrpLSMCCnn210jd+
KVQsy1VlGbBm5r1Awjtxssd9HJGADiq+q64sAu7lU57HmT3rIcE7JA3RaqpFLRayml6zoRavIm8d
TXS9VeeLPldksBvsRipWXwoP4ltAWn+jUpn8qjZXJ6SysC3QjHC8MIgTxAuxarXOlLCTE29avsH5
33LqfStgaUI4nGC1b8vZyWCViY+wodRW2Z6L5GbBQscMiSGVSB8B4XFkKduBvlgRFXo/AKHdsTHy
W5d9Mp+nMchKiDr3iEy5gT+8NK90NirtulUcea0lSYr/E4BQ8pJaskOErcWTppG9eljvJruRb+zO
ZVysvlEDRkcoRVicJ/cssdbSH1t0U+5gxyFsPiCRqmS12/85zIytfEbxHPmc3Ch2WTQeKGCo7iLF
jC1B08QzmeNK/qMqBOKnnZtqOPCii+hT/Zy5VdhD5Fet5iEum2FLi7XClZAU77aD6awZ0/REgQg/
sK5IwloHNAv7CJW+dKhnz8F7av7jTGk88u2KiUPYIORNMl4hox4W5Ew4hj56lQBqaIST1zobptjg
v5CU7NPlAmfX7i5TRmjG79fR7pQFogYx6bAgHfD0ifsXmi78+N37tY15PVvAAL+/6jNcWX9sn7GA
ttzyhs1ZBa8iatl0mmA3t6tf01gnmxOEh4QkqDay5hIXR2nMLa9j5CxkWGCvG8QhxDbmn+Hde4Nm
sA6Ine4/nw8K8XTrA9UjzcuN8PEwuV/Uz/9ch5MgE+fb2EAYaElGn9RD10Rxi+NBpmATqLzEZmHR
IlcH0Xq+xY7Pwte8fz/SOHCRX6MmvSjpsGdtD4oMRkcCmkulnEalAiUeJn3o8pKr+ZHruLd6EGaI
xOPXpEJ1Ohz9EcZ4oiis0skVRii7hVtc01QczOdWhIyZ03GineooSVMxoU0p1xHJPYUlJD7In7+e
4+Tv8UYc4SjSnZGijX0YLkY6J3z6dufQv6LPtv5cAIrm1fAGIOirRaJAH2w++wmz1wh5qdfVz0/n
1ckb7CfK3dV5GZTwpc8oODI4oHy9jtbFSRIs5MAyUH+US/98UjWwZ8y0N8iGzr4E8CwN600H4ZZY
mPI8XICT+TpnYkulURDfLB5gVro+iWg+JYu6aIfP2NJbBlQBIkn3CuZkBqwxbbeSF0zJBTb8iy7X
J8Ek4EbtIcnsjCcu8GeSVjCCldQerPhXQs12I6cThIDRuroMIQ2Kc8zhVXXtWx5d5xlQNM9MSDqT
jM+f6hYdmdOg0UGAuScCJI8nY4UgpN+8DKRvS29IkDwGMNNUxLNQhS6v5YGllOb+u4XeDnp66Hk2
RBBA3t8IzEEQ3EUebGeYAvOPaUGfViLAgmb4TfSPYe+yzQnVmkzNdK+DSW4TZ3bc4wbpRklGO3sX
L6stKtQ04PfyImjqQmqPycVWlikPRsyqieLOwTq+rbL3x2F2fitZbnqET3fCi0kOubQV/rP/Wq4S
RkfuN3D3BHWUtd7Ikn8rgj93TGtoZZdf+aRGIn0dPuZ3jEWSJcmAADoGy7XqwNCV04SvT/W20Daa
1+fCeQGyJnuV8RUQ3N/oXtfEFLfoNYdsJRXtSNWZf2IUDVW/A0fDMicRGZ6Z4pcIVmm122vVB+6e
GKGIjjOR+VXkD8VqgAynGwwC0tx3nS1g32AGOBl63LSzE8wZJZOg4Ym3G8t9lLI5p14By9IAqCqu
ffFQV2UgFLls0nIueb1hsdZxEZV2Ev++sDrD41DxILGWQgBoleYivq/Sie3gOdEz9arLHsVw8kHp
1Gc+byH2dNs1BVunD+tR3rvbpg6k99nZTqDcmf9bB/iJWKCLDfGfWTHr/wXtNfT/lopigsRl42Fm
HOoGl3hjacv7QLH6YqxIHYBrMEJiGwphhRb+FZAW0+Sa/fcUPXZ3RgWU5gdBCoo5RpRrlBNHpcJo
tIn1pRhSK1IKUKxXNSqKMgcKelHUPTD6xaHTSFG9smI9QbvN7uuVuG5EucGqoNeimRgMaEqw5czQ
A1zNBuTiO6+4AVG2H+ZYq3uAScIF6fPP4UXO0MZqaemi/JHMufxhoF+cn6kQyiAIVlmeHXGEQvr0
g1E1WsB9U4gs4WlHv04ooUUktHUmkPTio1So2bMbPOjVYBBUNkwu6pkTz/pC3kx4Jd09cv7s5F8t
zzThLv/K9Jsj3MZHLttQM3E71sC8jlZyCFe9ldd/UV9sgwelJUaZsZwwyOXfcTalqJgNNy2Me3k7
vikgote8pG8ur3I8tEsSNJ6yJY/nZLI0cTsEybwM903dUMRhnQRmNbmMYT7Nw4eLPOokYap/0nEK
knRD89m/eSuRfuBYEmG0U2Tdx3utnHl0vNAnF5hoQQNDaY4lsTafry3BORVSaMRA0kXitqCujQ7I
ZSgF1/E4dohQhi/7IGAs4TxdwJWZWSIdfrueFjGnaQ5dY84M5G12gl6/SxpGQCqrq5rwHDLhknMg
Nkm4+J5hADf6Y7zZ+yYA21Z2bUt/SJ1NBNPKTaO2pCNw+jFl+fZG14cmvwZGYvaEqq9GG/XMidEL
w8Ajbsb1AVeOCJTUMFB8inYfDSccs6aj3VobLfvtoku0jchlje+hjiBCbKa097T+8Xg+7wUYXXnp
0MNX3sJ8Fs95Rc/5JfJnPqbzxeSoSU4nOYtSAq6QZYPp/91uf4zeqoFpu9u3egHY1gmII1Pq2NLV
7amf4s0vrbMmehlpXPp4zoBvnFz3n9eHeQ2AGQi4jI/staA6E08bayH+kZBrgJsKv37GPttCVmzK
bWwh5Yekk5CF+pBauJDFDiVh/t58xtf4UzLGz6bB0wSvG9i3F0w4bZweOHtNH+6+5Cex9nGLU4Sc
0zdp7T9lCfexjU26yFm//40Ek1M1LdoiRBNXAh3g7zViMYLZSqRFNzxTvWSNe3t+6aXhgZVtcjlc
0ua854R56U4a+JflbB0TZLTfsNcLo4P9ZjsLniAQAFKKCOUzdmyoWqADzxyzGZqiODphx5mMxnYZ
6GrDKFosrRpu69BULQb81rKeXUMdZ+ek5HHZYtwO/uQXJKiuH/ywE/6FgJhFcHZHHFTqkcdukp0r
9Q8ZiwX5vxLczNGUzebcJRlKuQAynTXnvoiKmpZ27KRWjzYjclvxUcLWVO9hPcFtb+zW2uwBiMPn
TNiohJHy5xmfdRKrchiDMCkxvzUxdUMNPYyqfqATI22aWEVvDCsb78vws6bCkutXxsrBy+nWZcDy
sXju4QCOzRiqIk7lvMLoUMxtKLNOZFJcxCBM11SBxUcsT7uDxPtllYacqt0PCSnOPfwM1x/c50Z/
xewlsjoen/mcBigYAKNgdab86joelWGV1n/n+s8sH9ImAdOfF7v4MFE4RvWhS1JGZnGPn0RJzrWf
VcXD0UL6j5msdG/5BBHv1oMqPJQEa8VZD2o3byyxp7DMt8EyCyfGL/6Rwl0cK8nWNeN/xNlk8/SH
FaV0HxEkUkfpRj1mPcPKrMUuVFkrNVGfMyWRva+GHs5voR9NWno3fNjIqkJMjrpNCRLdQaknlMiq
OGVKwlsWVr16a7ZQjcjKzqOA0+x26HSiPLO7cHV/FVvit+TX6oQGWBny4gyGncPPRa3AnQsSRjix
J6V7Il/xMc+S/JnyJ6PmyqkI4IQpStjYxaVu0WQvseF5SvItv67yhxtuDH8PhkYFnVGWRjz3YORR
Hf16jJfP6GW/kNMeRd61es/xXUI22K3gvhSa/yk5RjdV/GgklYKyImKTpNXr5fWz6gMK/Vn8ocF4
MwsKNUiEEphjHN2a+9RKpPc+pOaz5Vt4xLbgfrndhSbOBIfKsWZnct0S9wtQglXIX46s0LIagafp
yrliGP+ySBGs8WAYoIBgCJmDCq2o14vHPuIQ0zS7qA6vn9ssbZrTN1MKgFs7rb4K8qTLWemtg1s6
fRAuj2js8fXtJ3fqygxcX9Snetz3OW0ez5hfQ+J4Tvjy1lA+LW3Wf1eK2kGVRzYnCQ4Mo89NR4Ru
DFkvVk4cIs9MqJq1wdkA+/86VJc4xgB6D/w+SeF7pgd++LcwEVpSf8bRFm4lASDtc1c9ADkqSKJm
103VlXP2wuxRu5+dkj/1bczg9A2Lj5qMD7d1fHWSccVRA9addkx5E6elJW2KC5wc0dC/7mbhewub
TnWC4OEX2sOsDdeaublbkzXc9BBAEsmhiCuRg9YJHAO8PP5UaTuiTVIzsAKJwoNEluc7DN9L+X+w
jKLFTeqSRJtnIDBh/FzZpfqlufOcRspUOJG5o/Fz75RNZmzAdZskV6bo+hN6iHQW3+JzGzIkCL6V
t/wlQ0AgLkjAhsmtQXBgBVWV4eLwhjiY8OSnWPUKFFUtJ4eQkjuczjVoywbszNHgbLtOIQs9MCxo
IfXTxEt1jve8yb8Y9DF0SEnzGeJdqJ+4ZAR28tLUXS7MwQtiuEyA9QKJs9cA+vVKdivlUU/MKS5h
q2S/YeuiQcgNezGKDJEa/lhQw6k4gRf8DZ6Z7f9TH2VckVQQiLa69v9KWKUWYwQdxy2ZUxO2Z09D
dUD5y9Cce0HB+C8Cf2TTIUV00E4o5okM8fTvznbA8rrTayVAfRynBJjORduuJDL9q+C1IZHpjNV5
jYLqfWr12+IkSGmy8/JE+wdOGNOq0afxBJsAgjV7++OAJ7MJZHh1wzj8Pfz7Hz72IQUJmOvoZcfy
NNrIJLBbEePVfdqL4cfoLc1g9K2y+n5v5nxLhESvwgSub+PxyfwMrcQYaIgMKZCLWHCzAuyAGH8m
S52UZkZqOmBYcN+wbTX+gzhpVFf+kP9AuFu1ePqhXGwpNJhSRK7UphE/goZiYJ+hidF/CTQXAA/M
3w96w+xtwH+afxoDX0eCqyDH1cP8bShP8iHeQec5JKjKRsfSYhIfyYUUnN38tuRQb4KQB5SKK3WP
T4GxzFRdk8GeN9R8ALt+/czz7uS385znS5j8un9v7jmNdPu6Gm2qflQMBH5y/589wjtdLbsxQyxM
Wy9jvukHvRLcmP8aD5cVR604rkyiRpC17VTmesCQ6bFCkRD8UoNDOmIBw1GqBjrj9YaUDFdr/ohe
H0zGQI46d1RwJK6oJNRKqG5RtKAryWawy7qtfVMEJ3VnxQ1NkhB6ylakfXPJJqP6JwuYnli8AhHN
28P3o1z4SPSdY8Lk9+nTIeaw0UajeTYEswQJxpXx6r3iAGQqDVLvRGkhEkEpPVv1Xh8bDUOOrnST
e12Oohb2TC+1bMyZSvkKZKsr5I88WyF1WPL0UvReZUYpQ+D/JdlhrJkpp/omfWye8ghOtxHIk/Mu
9My/PBYpq0wdOpZC2oDF401y/+1uNs0DgFxk3nw7t2+qNAkBZUTIapeI5h3X4AfPUx3zGL5TP5Q8
ZPwt9mO616+kVnPa8ObGwnzuBPMm4q8135yu9mkd51OYYbrTfccQCodE4w1nBqAgFC9V4C0EWGVq
Tsc2M1+vF1eHsiai3pxf/soW2ssfA6vtu7WNDbC+jo6aB1WgaZIN46L3MypzZNSdYq74OlkMJWl8
08LBsKsbFDDdQe58N5k5PjUN0s9upIAM0O9HeW0xXYPWJS7RJIF9pHogBuB+jFfI6dtAkXFab97r
H40h6gWvLg1h4JykQFM2sAXJ9zf07kTdp3M+AeNaD2zls+tuFUktsv2x8X8bjyv7Zhn8GSfbF0A5
t9HpSo73ObmMqDTZVaeOvFnfTXsoFdqTbbe6G9AGpQXj9hrdKXcxbkOzgGOkNWeLh0A5CLmIkgwI
kAwNtCSKk6zY5u28kwqdgnsecKSciWLXIO9ZHN9NLuUYaNYQ3H0W8g+Q65oaMVx2RvAdvr/NFmSx
TGQDirVEQLdfHPN6C5/i6RCvrIYdj7JyeRz/qKzh6vFNocnP1GXNcEuqZcssXlCFZU9EVhEi6oFf
px8OMSZLY5//07Z0dGP13h/TU8e9TaeDOwL9buG0PI4icIfRWQYOCekO5ttsXcimD3/FgfbibN3J
6/gNNf5cYhVehixvFCSSeLrhh8+zMzItrfu+znZUmaj0Qri+IIasgQyVT9IEFVjKEiooyZh9ISt+
9ZqF0bsCP8E6j0CiD1jmN7MBXgX70RsJpHbtEZxrd6jzJ9effPBkybtSGwDU+xi4/8f9M197uL2Y
+Z/u7WpC/tdSYBHQ2BxCfhhOqZLzfNa3RAh89J+KMiebsNTCFfUG62fLnSJRvbBCiT7aC2igQN1n
dgUPmCC5S54j7jQ4dv0kAjoyVlIwVHr8qV477WLzvefA0OrBS0XyUDXPReJWokxAuTa3BNGRYEBn
x4mTD8E+PXsysgm7WY4xEkw+Pw5/u4xfrFMPvXu51BJAtjuQwsOLNdX8UHARREQq00eDPWrR3YIu
rotrfw8PPhEYaXYv6dYTi+GSBZrhoVfKrYWa8P2jgyRbs+9T2tb+FwD7miK9Wb9FlRIJy1+OsCsl
ncY+soSblrsGHNHYWyREMNpvCwMY6dLjHxxG1IBiYL1+cSJha8eXNTQ3I3pyWXeP7D4BqJdoTbWN
rpYtpZaEiWZ0AP5xSmGC4gW1x/remTwKziYnYb3z4TIHie4utuOH7l8R/f4b9qn4qJFZgUaIeD6E
iDCriVBTbCxbyuch2r2pG6vRbWjL33xbqgtEVnlPYiOObAByh9NbKiEZdSg1uiNtBg7UjoxFxvv6
xQaQjxeCsSvqTIzj91zWkBajlq7LBDaxaQDhtVidhAcFEXm1lcMRsAINs4YgqmzReO8DRdXYFpMw
c5x1hKNt/IeWkUGq7MjNrouFfGX1a2r4VZU5m7A4HA6ZodhT48pr2KETuEQFYHZP32QSSwIKynOn
1WV+gpa+C0tpNxKNYsBcXZinXpTGzAwv9JAWlPt0tlF3tu3b4Fm6Ju6CmauduohmvvSiozms/0xJ
vrDYEahc3IzTkHeMAQOT9Q9q3tPFYUTNeG0rlVVqumvKocqsPEou+FJ6WFnYV3kaejxZHpGHMTKa
EEvCtLBVwhprYUYbhwkb2NFSf/0o/oEQ9K3+7CjAJYvcMEaCvBfwXZCs+id4k12kO1aOoclG3sFQ
LM6HvfwC0DS0gA5o2m+NiyYZjU9sripfd1xTtvW6RqPTpgHXezpw5F2zcBkrqqQi2C9cqNxTyC2q
aOo5tvX3BBZuq3PlUiuZsEjGbGnMMnbShtj6rfixCp6LTarVaXVSjx85ykCtDj5eDx42NZXg5pws
9W4tSqEaM30ZJlxlFRW0A7A3Phr7S16XxR8iN4oys5AVX05A7SubzmrGRKX8u68yCaSFeYqLFZqL
SzXyizVmyeGY7k/1ofF6gctRL4yt7ueeTgWjn5+iqteSsHd6DRx2TtxgJavpl4EPacQ6lsl3ihiM
ctjfoX2KZ/wj83Pb4ja1ah4+yBvFA07Ce18nMTlfU18RaIaXw+/S1AzWe81tB9yE5+AiIQh2TJXB
t2J7LtouAGM8URRGplmqrCZABC13ZmMolcHHpocb5GoIEA4JUEtsI9LmFkeiQwp8BUkIrkiswdr6
9WBhf73DfH7pUELxVHAlUivP2k1CPbxPccBmZLSk6Sjc3HUekOlpYsWgAvAEgY+3N4QW46b4+CCp
9bIuQQUAcnPV65njDUNVbIVO/+FUWXyOZ4kDTsS+kAdvi6ijQIH3rSvi5uLMNvqSVszJa73IID78
D6rY2MUh3W5vFzgKbfoJ0tPZ/7hK84APUKfp6JOZj3cjlEPRtV32tZ6JfQmCKAFoERl4BedezKhU
7c5iAFQowaTIekWLhqoYqev8R5VLNlFrbkDG+0fbK22LU8m/SEhWw0X8aqFX11GURcnbB66jATDQ
t1d285WMtPHveh0XnCoh6yjD5zg8qkk8SJFnFHLKBMJC7pVErs7J3tf6WGGkoqTiCALvdqC4cXYq
tJlMaspWIKtlZzMKOZ0leTjwUmqn/KbZ2MAhdTWFLAItTKSPUT1zJacx6lshByf23N0GCbrKQEpf
i92izAscK4Qe1VnvRgOulJn45aceYnuXMmzQJM+XCOXHn3VLB+/s+sFD+9xq9hm4MmopPSxZS4sE
/brWvFNNiMK1i56HVP+Ga9wWsD2xBByiBmvf9sprTtStnEFR36GIF3lSzjh9gaXAeZslKFqETqQl
rI8UheBR8ri5SqFkLq4xHzieR4DW2BMBwJHpI9Jw3sGrvbcNLH0LdN2OtiVwJMqj4vCG6cpSSAzq
L3MtJpcp9TW3jtiq0rLybuoJOrg9GUH+uG832xlZvAJ9Bw/p84pwMsZ8zp1A+1WhJmBEkmZRDsIX
c4EamZRcgO4eT+clNwTt+Ya/1F8Rhx9ZAj0bcghP9hM2IocwTRSWdW1JIobgJ9QpNhh8aQyGjELq
/cL8KUveMOG3TqIgFECGU+F+gW15FOLMECkNXjTiTXf98vmVxCqyjqJ+CM2UfQeiVvmaTQEpfE7p
6n9uMzRRBMflbEhFasu7MLMY36KLNvO2HrYHTKNa6+zIsGvTEvkZ3KUb0TQ7dpTr7dR2ZOXYlKAa
gjqggzS6tsfWYjPk2YsxOoqJHkzW0oGaHvogozAzjJopxKPJJpp0u91clCetYRNQp5bFHcnERdeb
BYZqK3C3N8395UALqVyPNIS1KNZj0yE5fWWPKxpvFXQw3449zI4jNPDUd7kTSHyNUjR5jgTokP5x
3Ok7LK1mmp1b7Ax2SKEaXfTD7JGnHr+g6u2bQf+ifeV7Ib384bsRbYMoRYMONlT881Ho+N8WtOwt
tKf+8Zw6ZMRoVTS/Hdg3m+xxCGwSIsj2NR+tNhvOtQL7AB2H+7QeqQWStpznbTvEWNjhWKu+8oHw
YTimct4LMwh9qKOfFD0OUyMGCpR1qfPU5VwS/kO8mEyXQhvuJZlbyNLBuXynHtDaY62a9Zm7Ropu
aHOrzq2bW14kWuOIdYIcQP5ffnCo4rk93eNji7t60KqTZ3+xRH7cvanihevFEy54xGugo3lvmRiW
MJIlAYVbu5edlh3hhE1PKDZizmdKBKaoIbH7itHzuhvV+ZP+6/3z3V9AnHpKAl5wKMFCWH9yIZo5
g+tNte6j3TkEhN5R1jF1zc8k/iCRU+FA5qY5l6qqjDdF6/xOjFtfHktvqTgLaIW98FvrVb0Xwp/O
k5MywOax8dZhVh7ShsFDwN9mIkcwdNFOK3LEhenO9mXwrzlna7T6EdlKwKFNDz48MHGnBBAeRqSj
xq0gJwdtRAgDzFN3t8ygjkG/wpvnTcZCnfe1Z2UagmOQ3Bh9Bt0D4FjjxrDbSkJSemuE14flQIG5
YFUrzDm2EvWagU4bT30jrTuX1UctZ0R9doDQR5KXR6qSah7UPalEWhMjgcjbvOaODZ1YbJzgHTMh
S6GAjtaKeOzGLJQUCwZfrC+a5k4oczYapAHFTHoSWTQqKHV+l4kYcMXPxOGIWQ0jI3KHZWKJ4zR7
q27ZO5bg6tkZUE8fbfEHfe2EgQC5T/1DCfGGzAJkTdCLto2WKQ33kdca+9+L+JSeHyDFSrRsxPWZ
Yx1Wl9cx/SpdAwOPRQ0H0vQISc5QjLF3jTq3OPQxhVhwWbr6tk+wa4+QDUNL0iE1IgJT7XZtquUL
GwFX/vebooOHJytS2M9BAyrjAAleytSBtZ6lVm//YBACkjYVN70UamY21y1FTTRk6HS/53lwLFeo
dDcCv5X1gvVF2G86/7Cj6zHWVM7mQtfPx+g+B8IPCLxwh0EPe58MFYx2GWwNKbQ3ygiCYJn4zH5Q
kz1KlP6XzrqaKgKwZnV8ltPrpoJo0mILONAGW+Dzek2XN7GDSLZQ4dSeTv1Z1ARzcLYbRIAPyB/1
qSKfBUbH7EkqCNZqpGsbkwA3Oq2HlwjUqWotnqrGYKd21FCqv70hHZNsUerAbozvwT2VXnxWt7wi
LMdGqkm6IRcTWMElTX/bjADB9Nm+dFlnLEaZv6DMLXNTWamGL2Kib7MrG+/ESVptwN1JpcHcckGe
neZzvKPlWFl0EwhBqH2VCS2EarXh2Lm9WRFcX7K1C4fgAHWfjxoEbb9FBGJInPThqlBmPmNMR34W
/YnvJJnod9YrrgqLmfNuulXdHF1yrnRnoKazup0OJJQASa876O48S7lPNCGXCcZgDt0eR12cD9Gs
cHLRclWCIlsBx+B2nZrI3VdQwa1Iw8X8+iiADmFPXXdLU1XkiYm+heFVlbil5KfGcl72c97zeLzF
e4yFq75k69Xbi7BZjsOWH0Rh1eOpdp3Fv9uuNCj8bl0REQ+eUXGdmipymCJU9gratDzCDz21Saxc
OWkV0ZE1xG3CjpyiQG+vYiV48bPDEIer/GAKrnrb/q7s1euYUFqDqY/uO4Mu/ji1DBdMSYRRKc8w
CyrBM0CnuBhpPk5zgQx1nWQaZ5OluSiEg+ZbGxUExyn8eS3s7I3aj6KDIX1laaxuUVI/axL8olFJ
xZAjy5lTE29UhsV6tcBTzYSGnXlDr9B+IOgALHeYe6wfDU1ZDJKTIcgv5cgy+EzjKiaBidQpm0qs
ta521hCFJ11BTWQfhvoQq2o4nOURrtAJbR71p6ghq4h0ec9k1s+rSHH6nwhKOyO4gfVCiOpf/l/d
zSi0nhE7aBlZKbcwh2k7HulmAIbDGu9Gckfz0BSFCApvbDO91+nlhSuyZ5XGXwfE1ctzULcGmc7v
zKmUHZ2CUjTjQvSTmgzfBzOOCMxqGyLlAk86qKfOX74U4/OsePvFSxr/b42byYwK1vlzWec95PT6
9+wcB9IkI/d7EIPn/2twWkuI0yO+O1mfYQiuQRk2znb15pAAr4cXIDh0lYdqs5CeGwapmPW/lVAZ
ZnaV6XSR1xvWJN0+HVmPFcCJVI1ELsbdb716qncKZi0uts6j/5XqaALlteYTy60CWDvHpSGV1XBX
Cts5p1lCdydFj1EnRROkjZIzOenc9SBOMskyGwMvwZX0M5nI6eBd4/S9zIhRvU7La+H+cYE0tT2C
Oy9KpoLZBHr4IsjgSD1HDPjXLrkt5iB5NjW1ST8JwL6zmRipiZsZefDHyUEkku0Fd6lWzriTRcL5
VSBAPvK+VQuS0Utp+VWYDFHYgccwp6BEOx7nW7rtoImf/24ctmSiAame+bbCAbLZB8oZYvRBZZrz
ccLGNDLaduA2kp6UaKm4XDJwGSX8rJQ0cFDI0nWHVSB281ypV6KK12f42T8KyLcLnvwcMMfihe+M
T0vxfG3lKdPhzabpSwq4IyYdVl+N22AJJQvXP05SriJqhJgP3CmBqonwahmaHCn0c0hOd6RdFLUI
InzrdE9rb82eus1bpy1Wz3V0ZZW/d+VHsKgPZ0p4wM0cph3Bq74nNTs40rua9kXV2ykycjhjF3Kr
+wVXzp8YrlCkZXv8v5ovCctEkjos3UfpIme3rq/tSJ2F/5Genxn4/kaPcN8eUg61Hgyj2Co6j3XK
sqAwV8DlXlsNbWvyDhFeXkh/dGUPzMe4B9g0jTDUhsx39osUBGrxMsOMG//bAxqcLgOQl74JY9Oh
a4yXn/8dmjNwIlPkbgUfcN965UbvAbvpJwGvby+Kh/rlFXJm7x7iXkIXPecNwh46S7xTX291SJiV
WeZ0oMUBa5zS6ztjhgfCfrO0MHoDx+rqCjs1hSDsrXWu+sGyl7a5+uAeCqThvEx8TDdmS5AifzJi
EKN33J3sgDLZTqG1MniHuXlUBkQmeZUvefC83/j17S5xYvn1QPdI6/xOXog/hykfsCSLKvMjIm2a
OuMZK/lAfIEuN7WSEj0/lVXE+Is6gaR+En8S8fwX472yuKfJA3nIvTeJM4hOu5Mhgcnim7o3DCQV
YuR7cX0640tc1uCafrIuHnpSLTplAIId4v1mbZ14kAP+Xmw2+uDF1yT39q4I3BJzwlyHMoFJsZxI
d2bF8RPW0JbTidtTk0MUiZNfFjJ2QWxMS53zRuddvgi2xhSecdTFcnNfNPxLf/MX0Xos+/j/gGdp
nU6DdM8s7eL3igaNnWbQwYUJKPaO/Hyb44T4bBRukCHoq7V4H5tSII93CQQaAMoHva+Cf0tAqC86
EzEnIUhreT13yNVn+AteqEb3kRoTxxD7C/03SHhrPFt2nx1PNTgxk02mSZID00I+PDcvskskIO67
5ZYhLDk5sANV95rllfD2eKSag1Ka54+0/2in5g1K53/SXQmCEOzOx4FiHtABo2sJ7ufqXGco49m6
y6KA0RioP4aZyCKx0/oPNftMXpA5HjRy8XPegSk9fgp8Qi7LmjBUAw7Z42aXRASEBbed3bpkH36i
6C/Wvz/y3PrfO9GytWcs84LAPYF1Pp/+blZi/7NC63NcBFLSNWBqv/xm1E2SJJAtRieuMarO3n60
iy0khgQJ+EvpDo8qRkJi73H6razz87M/kdZoALwFI3u2AQ+M7N6sAavrPR5VieI/fiQrtRVbWllR
NeSMS0C/Om9KYXAl/N8Zc/yrHUuvKkzmWmyo7/JTHqzV1/GekuiJUISPjwwmNkPQUuJzUFXJHBbO
XxJM/FzSK9g1U5+r8tlyZvOtteSjRtNTH9BGE/zt6YRmmue3wRsofSWb+QuVdPr3byC7sjRC1RVo
CJvLEFAssNJ5ZVUxDACJa/4b61GFUBSlp60g7wT3/LT9DjOOoY0xSXHrmsKelG4PuEbgfKeVKAPY
dV/dBdVjQ6K0c+gF+QBqcduxR6MORE3Wcxzpq4vlFQEUJkROWWGP4ovFutvlmCYCH+sCh09xpDU4
A8ncOP4P3GcKbFE/ChzO+hqVImomorlflHOs848I8CMCrF2DAIAhZRsUYyqL2lNsyx4Gv95ktY8k
PAWL58Xn4ED2g0y+xs6psOxOPuQk2MqlbSTVfr6qzU058IoRXU4wX9GiiB5bv1azgCDuGrmdNvCH
1OJQ6iEIavtnh8oHtCGqJbAwoGBBgalBaV/vt/WZmMkJ10WPHeMHmMX1SkruYYM3GrGBDMCJvrMW
BKsM4Z8mjm7nyBYHPrYzN0ZX+xNgRvKm3JberMl7/5Ml7mcDNbOSUk/KVhZ+rkgIX5ZDeXxdtPir
njYZD6HyQWulywGyNMS+B1mbu2HrVu/sE00QTpU35E8Nlzc0xVHk1ZXd57kSXtBW3aQVL1tHomtk
7tP7nBmU7dW4Fjx9ucHoH2Vg7Iradd/LEmUl5mh7XbTCad23kXZ5Lii0BtsaukAEG3aDXwviD5d3
g3bIe8saobfai324Duv50R/VGq29sK1dAsGRS+5Se1MBM6sITR90Ndr8B75/9GKNE4hJTTSc119U
pDcpOeOJDTnW2nISW0m4Bk2o1/GOAFD9ctzg0V1XB/zlxiRLQxV5hrSU2P5mzdIaIwiTOf+zr2ry
9uo5HVa49xgyJxAz+rCip6O/8MxN2cs9BwXflLlLIhrhrkFQj6RBNrNf5b2AkZSWq4YAl+K+Tjso
6DTEZFmLQzLQ7qgI873j0nlXJ1hlYHPnj2ILsHH5zBELnQFgqu1cvKZmM+FmuCOKgdyawO9tj372
yDxy1yy17zLR6Xtv6D59bQ71b/Uo4xJAH/4aQ8Xsr9Sfj6gSQCqfFratctM8MosXMWEmhQrWPwra
O5f+38Tf1U4BduLTvErxCv0udZ/OdAEge7itC2i2KEzfh4O9HqFc4bup0lZ3Ug8sq6q9/BPrdK5C
sWChgmCrEhXa7pKjFMQ9A4iwNQ0snK3ITKJRU16vFnFaWUNx7F2zqjxWsqa+yUwC5G0YyOTVZIjD
DJpHdfPL7se3qzf0FNJye47Z1LS3SLwYcDfUyCZ7ZHzgibGn2SWPKLEH4q5VKhruK+TXWWY9oXxN
MuJxp4RPQNRdb0e8bYasOrAslPlChY+c9qBfnsT2awVFD2EuLXEEjJRcVNK5E9Z261gFQUjZjKXa
P0nJGRSmB9ntneyh7f//gDZt1c8oWeLqBeacvrJnb8291lQ4InxdnCl/zeWJB5dm+ucRuS/gC8Sd
JglJeUUHrsga/9TnYnHs+FcFDqhatXBpCurPV7ezIL4un6eWU14LgumQlaV55Iz6vRvNpzlEmctB
MxCI5J1ihmf3dyx12KVuCd0IgcdleV1c1keA8j/8rLOT5+VBvS+0zA4ECHwLeG/ylbGgtQR4ktGt
sfFjmMLHfc0ISC5yYQLLOky7/yNFg382ySBcm2prS6wHbGSl0gioMgtw2ZX9LUjuprbowmCuUQHG
uHq229L2yuoNmyXhgT8JwDznDPttg3v4JxAFvu4lg3Bn5aWk+g+MQP4eCRE5H8nHGmDPeCKotvMw
+RILJvqDVmujZAHql9VX1DHlB+T28P3ohPWZugxQasgpSB5SsBOx9qUPi3G8XoMKmliY1c7ed/11
tPdBv8Mb3/c1oX6GCs1S0ruNcYzdqOiCGJOaHXiggnXCSpqIUV32TxYVT1dZn6oM+TAPPU1U02vo
QcYYoMxzpi6iXI4QiLG6LJPxt8py6njo94TyJRr49omDNF6bkgTyUTvDmEc7nQ+7rJTGhP5CKTPQ
HZ0XJ8YtlZUU9tDTWKjORlOQg96jHpR4OizM8bPhVJKjSZ/V+kj6kXoIqb4QUyLUxYUcqvgusgJg
f05BbdGWIULNhAMsl/DihrigD116G13yaVb+uOk+zvIs7xFseFsh+1sqThXw0kcU5DWZe2PDMnNg
FG+gC2d1tJVI6EpUe4VqtMAP/XUQ2HjjG+Ahe3CPJDIYOaeOImq7hYID5aGN+wmIZNfjMYJddmm0
blRU5MmZaDNc2MAfPu2ZjjpnMkCy4a0hCGKTtJ+8ROPavDipWQhr5xbHFWQM5qfjTnAAXwzeJKYs
UsJndztK3/39HA2qYpgymJltseVc/HjIxNu546guvI0Yac8SwPBrFYfCMeQ2jCfZ3WrqEKfTux+D
AqMT+tJ0MVc6RrJtSt/CLhV9yzGuLtexFHl9Z98TA3hEyOn9ZBAdw74zY6FREu0hSTA7GaWU8adl
OwYMcKanV5lXdzpzplsexUqfXuAQcmtXe+uw8sHVzBDyHYSu3grl2sbbnB4qDn2RKxiD+SnzizHY
e/Sl3+L2TcRvf+mXG5s6WGe0sxw1P8BBfivQexcwieJpc/+p/VogsXnwpVGDgjqkLs9cVrJLR54e
KHGXhRJ/8UOBm8s6Dk9+SZiULpKnmCmG+iIMv2ft2L4TfAtWUYPVh57Pyf/LJA+cNoiwLXqR5b/n
5p48pCRgQfSCQJnmKaZpJQxOHZEyosAG9vsiJi8J0AWJpfftuof9jzFbKyNGvTQadQPVpDtwBRax
Gs1kON1aew6BEUxAYcyCvn1eWzxyil8VXrhSWzmqOwWxLKjZqzyyAzboxc+k1iXGEKnpnKzIlU3I
MtY/fG8J5cMyWmB0B+NdYGQcbLkc/S7nkIuU57PHu8DAxc5t252gS7srXckIC79gxZMqlKz37TYl
gfxX74lZuPQd9zNscWjB2Qs2YmsEW9QFuYxPefHS1dJ5KS6Liz6TgnaClkBRlFIswT5Oe1+/1INB
+asIIGO2CqdWLHq3CqImgNFDb1BHCws0vxVptMdahWOmcZidSC1pVP2PgoJNlH4gJwA0rfCjOFKN
4P/CbRomVxgMWnw2NWwSpRMkIETyYIhyI2GLerZfmfWyU28PbV5YhQ4lwIbixm931392QK97qDsW
JRoWnon0VzeT60gXNnvkg7ZVVRHVLRhi7VpBqPIfUE1YEDeKDdLcLUxPqQSjpyCt7EpWidoTmuaQ
KmGxAZ7oyJxXDCt55rUrnyBUn7Qi0b+Ee3BYAdfIMAvM04M1CKlSgMIHdXBnGrAtH+Kw4kzWKEJ3
NWS9KrAd98b6PN+vmExRWR4mbHd8Vw1yJDwSEDW8GFVCDbyuMVmuw0cSj9XlIdL1JUSwQ4bHzUli
2riaOChYC5LgHeEy5O0Q3CSH7eJ03oJo3lSCmuEDIfh5AxSK5aIm9P4RHF6yMoLqiFAlyDecJU8F
fb0AOlQWhCPj8AS/M93IxhjUhxR0HbYhB6UfHjsW4H5WZtmGC2PnHtoudvBQbtASz8uCxu+jGFb4
pw06pBrF+IIGFJwRrV4Z8I8j1c4qr2KYQOwC8kKWzycpqBRZP5ckdTt7dox61kqTm7r3swNyxrmA
LVmFtEw6FQNXiUc7nyav7covf17AA2lNpYr1DOZuEEqGjhC1HXh5TdjHdMcL89OYQj3o/VxukyxD
hWXNt0ED5nKSe/RNUElMSa/Uk2+XSjLn81QUN4XHBanwvKEoVlAmUOd0QEMbGlCHKuEM7SpJia1x
aOcFPuBWOsNSCThCp+tSQJin5XI/7z5yBr+o2duchOuhxhn3HQBJgvYdu4bEnMpvG+O50/b1vrcU
3RAB2aH1+7rDq/rJc4GPELICbazWgpescYDXveTQ8eu8wyNwlHRNGJB3uVc2RpvNclN1aGlbyQCa
Qy0XzIgZQFiegB7ggpyuzzzjHF50pgMbzwmPw0MGzWiib7BGt0M/wS7HOKeGZL4Wvusb+VPjErl1
pPIzCD2hy7+g2tsp3u7qt5tNhDCXtBGD87XrmYEt24TIft81iXwUFj4Oo7TCi3fU4hYz7ks1X+iE
XcgyuSzLbHJ2F5+jnE1K60hrHjIJKjW6Uzz3tRF5NzothvIYhLnHnbrMjYPU2zXNwtu1cXMtluhM
bt4183ErCW644NVNSB31nPU2mj4EfGgqne9L2Vfsannq0usEbE0VG3QBb/YSZv1H8EPpunMIPVKq
nK/UzDmO5qJ8xkmm9te6+td2OxswFTyOtFCZ6aTXuZfMQV8yhn5vMGgErW6ecWtScgZBkg2q7MO+
aJw6/QSi6L6xaIacg4drXtT1lUevzutk6fe5tTixeqIjHK9GBsMGlu7PVNk4tpL3fHygLRR9nboT
h+zheJbTl7+T8cbdKSpvQuRLmMyykrXjys+IRAP0TgUQ580KAZYbzuVSZTbOxw+LNXZUdTrno3A4
mRUsKLIwQwmUhYbwnpMDHZ4/Thfv5lSiuiKoQlXXGOxN8Waz6roqI0ffRx8oXwgkmBMoybBh51tT
cSeo+Vb3D9yMxJ6wCB2pDrGT9022RcPYeiF8fukITdOwajVr/OrHDQBBVy9ECGCtjZmbR2VB6FZ/
Gl2F5Bl5aQYcYz0wOC61uG+/buE1CwcFEtUp24k/8UQy3ljFA3A8h/f97VzQnuCTg2q69Q+kFYT5
8d4m/MnBcBJAwZ+tIyXz18EA4CWAlUk2v9gIiuiHAX4qEU0TJHyG0cQaBAXxcsDUPNQKwkBUwown
vckFiDJBbCP/KEmRKfCcI3xFTR13s9kqtJQKSz4whWN08JZ15vv6X1YCKZhV0WiETNbQrbf61Kko
5RQcAJwBtPccF3ndSdCItHnj+5igTdV9Fii0IbupI/SXFZZn892E0thWLogJz9PVwor88S1L0GFE
QtSEbhIlmqalZUNWSEZu3evs2hr6mWkL/PpiM0JRqO/BpsZCTUtGj2q8xAQ2hy1qFvhV4/mn38TU
pIh+xu58kOyx2ut8pXzd2fPONBAEhJ1VqGsk3kN1BvheBh8pHEtl5F00sHJ9FhVR7VNkCOmR0rCq
yevpl5B5caUjj40l0Q+Tia/nWr241jFQ4S0T+w5tn7mzfgg2AUIu7QScBJqIlbtNJcjcnsBG/VR5
0aEWj2Xpocg5QY8p+0i0VjOjUVHGgOZObBUrBpLYtZskuQbSR16/vbbE14QrnkJ4KB9n64mW4DLF
5EFLbrgJO6yUWkU+6+JPwJRU0EuinTRBorMbzEs0sA8Xav/haI2BalPJa+KEeGUBtNV01n97+pfV
aAs+xzdG/w600uLQeQ/e6x24xCoB5RvKNkdNAN98srq5ZZ/w4wAaGFzMvpTYYQkQD4IQyAPNHbKb
8LHaETiHh2gz8e70QnWo48xBYIR9vkmSwBN1KHJB0x+h4VTQfdoS7eWeqbpblq5tRYkLYH2F2Eff
7ZCgwKZPwpX4u+RO2sAfFd/QJTyAMbIciLfTyI9EOgMERVkxUQq/MCs95eFs98tSbpOBseXwfZai
ZzbZO6gxaTpDB8bDSaNVSMCRbEU6yPBtoPXKrSze6JhvPI7+dHBi4b8iI4goEuK6/ix2Q9c0QDnS
s9Dsho07pp0hTBF8ls0Rv8+XgbIvMjGnBOQE3t8yWwu0JFzalSoUAMxLYmW6vYCNyaZCG7KOMJgO
ZzazVNbKnwwghCVTpWJDR5PmFdQjf4472RrpKktJR+kkz7X3o+jKg8Wxd3EwVwWVcAaLSHHhrQOU
DbfoM3e1cJ5yHgHqTYcYddHdye/0tgv025PtxH2ZKsnNSiWtx99c/ZMrdskN+/sn+BpZ0a0DE0Zu
Ui5Odzu+TaiyHwyyiJaIQVZH3uYXse54V1RC3mCfGUGaopj+4Ug/Kz9tAELE6j/eOolSYr73nEvH
rUAfjdMAxsTo11214Ga1vNPs+ZQxlVucJhne3lsO2xPrBWGYE6GIKNc7o+Vo/C5VNTBeu1qdlIII
zd8l0Mjaz7IVskDZFX3/PupmbJ6/6bohBctzUlo+WVLM2r3rpWHZy40bKNXHhfJbpoPzIF4dtQQr
fIRGAOH1x8CksnVzQ1/a/8WbVFOwBloXcpIEexAZoBn6KJZ7AHwDNEMug6G0OnlQO5YxtFOcbgtt
EMkl/5XRJPTrSwAiUsv6/sFoAW8yOM+WEihkrEIW/idMsyP7k61gtB4wxhPt3cDbcp/hB4BmAjJM
TZykw6uvTSNiASxRKFAx+trwzRKN9zX+p09P7KtN/MHFxK+M9eatc3thuw9u74aIGxliAyGTBGYG
z51uBIonhc8ZlIV6kj+L6aGR6ciTGkfx3nlaonFJLC+urE2IWtxGKQDmOUr7bi2dfxcsUMOdme8y
AXVSx95wsddyn9gob+EhgbXeWsuIO/fD7BQ8ccr75A4ouvGBS5bbv46NqrDAvWRmTR22eN1hBKxb
WYPEldzN/lPE3peWlvm06luE5dhX8ThULI+z5lkreabImeVJ8OHhGpkJcsUpO22JplPX4ZbkZNl+
UvaacPBothuPJeVaxgv6ymSXR+wZb0d8E5bFJHt6C8pVDogH9PxhECAjKogsyQnhfNLhSjRTYeDN
oG9sCZMBMqQ3hPwfeAk00sirM47ZO9WZoX/aXTRN9le5cj3wPwIRX6tkyU3qQLdixdauyGeeTIzV
deOzRK0zKEZJerH8dD2QyglWCb+2MN/1vuiUD8PAoJTkNmYJpxVo+oRdnlx0QRT2r8mY3z3pxFny
Uwx++Wcr4ttGpt1ySwCFG1KZq0Om3kP9IdCrT2+jPvEaD9OKf5Up201j5VyFpUXGeczXNZ0glGQ2
V+mv76yPnLNPxX8qbTmq+nTeicVDqu3n+/EyvoqmouBtPOZJxzSzzvkYXJXh8K0xf1V/PSIGWqsg
KBkcmtKxa5WSfLhrOZ5NTqA+zE10OXONrcnQ0/G9X9Lo8CnMB88aK0ZYOiNiATUx5wMqR3KuMf1F
aloHlpPkdOc5JJfFYRXpElI+23zZaHMpXVZxv/BlfKwHgDs4+oP7R+ee9UhabQtyQMzM0yLKE4dq
M7sBs82bPlmYfWwufN9/j5yy+K0mI8ontP/Ua0d3PI/J8H9QTGlpOOtMifqkokl/c7IuZTVJlVw6
HRujSf87q5pBBO9t97TNQfk5dCwuz9ieNmW6yzU9/uVo59cOvPNqTZSoFdOFE2pDQ03iu4+M1A/m
peMS4lwxpNJ8ZwvSawulQnRK6wEAul6QY2KzlaiuCcl8usmqiEIOARx/b6bcgEotBw0PZSiq0AJz
orNnX7ElNNoOnzSfJ15D4W9Pz0WmDBvb5N2e9TV0jl3BR5RPJRoidN7rXG/6dQsTfR3Ostci8rFP
O+EMuhamWZWN5UPcMoSG7TPiyA0oXC7OiwoOtS24NSP23bD3t20NLyKc1fbQpG0V3xyog3PW2fBi
nTSAmSBQ/d9HSKiWapllLzfFIYevohPXRm1UcBHszyzHGMDZNeFvm83s7ou2HuvUxjAXDOg1C6NC
iNr8k/HXt1EG6HPhm32Qhl/KFLlSqYL1xkstq/9u4PATWPDZi/APMcC3ixUUl90whopjT9CK7Jao
rqWRUubYUTQqk0Gq835/23BGfPMpPaTr8nXRVFICukSfZsklJFg1966wxrd8fT90Ti7pntkcXUo+
cPavdtDLmF23MB/jxrXewPGHq06kVzplXPa3nyD8BmTo+u146EA63fJMAgMFUlrjPq56AP88aq3c
s7b8z1UDRX/2AnP0ks7y+JqINGq+yIyqoDxBggHc/3vkz5Pyw7mO/ZpVE6IMFiert5cd9zrXVYF+
D2QtsCVqfQjDYLfm9+Q7ILoZ4T4bwOK5c5W0Vl/M8FaBaYvn18gGIECwlJKo0fJWpCUnnnvKAxir
oE7RFDEn7/Upf0myicoGFqRbvKhbObxGyOwkXf0ChqJ2Y693a8joMRTgFkv1D15Jvn/chHXqhxuF
Olo0KBlWaKntu3pow47BCzZ1xpQZRZa7t2DD0r3fJX/uCtWU/7p1ExZl79Oh/R2wICsJRunIzYVa
RTetFCMuhltCN1lyLJbp5yTLJQC7eB7/bDEVzEigx0ljVVj/vVLgStHm3GINz4kNBFMlALU3w5dm
iweSase0VhjlN+7ppmHqLCS4ObKZJQFA9n7iht+FSc6tTyzKG9OBP11cNkgOUpuxbD5KRy0o/F0M
tqxIE5WcUoNeKRZEMrDARCkAeLMhmYByeycy3B0YhEdJm7EmKkcPrctLCEjz+Gc0NV3GOT6Xz/Cg
gBLt0GuWXb43+GNSEFHdChWhqWgjAA1bz3/IC1YcV9nxXe3wG5h6yvAZV0ZpUsUMSxix+yShPDzf
UxieaXfwSEPTHNS4pMQ0LSv5zPRZ1ZjGhYuTEmA0B/SiMmsTmbwN1QBp4xKJ3p/sYDzr1aGwP2HT
GIVh9k75aRf98A4BIekdKOMARpFljfpc88cfcAy0XKb9vsaFRwU8zCKaLC9luihHljOFAtB/13TW
nDW2rr1VsvC2KpZjO/RsG5CzUqx1FCqbE8hqhOvDVAGIcaHsH0k59RjmTt8agso4DfYLvvDb2ps/
dT/PJfZt/HLXxxFkpElqiNOgdkTBIYahX05YdY2Plf6mKh53uugN7qjLe+uXfA1zaqmIBVEtFkFA
x3zosrXoxXgTwuWjEUqW4mijaaC007jQWRr6YN1oP8zKdwECuzbnLmx8E7TSh7aQfOp+/61N3EPE
H8zeCo7hR99tMF8l9Gnp/BfPqsV5bHGMhmIt+FJw9eHN3j792s7mm9Jea3g4kQrjAbx1p5bfcJuY
BbFmUOfLaJEudXa9CK+HD7AyFyDPcMMoAiXLHzTcyvqCyqhnH1XCi0kclMNFSkivZL/TSBD7Yeqa
djsC5KSNU/QL/yx3++/YJQ2knFGgbB68fgvj90sOdMAmv6B6LfoGGle8PfNdHTO2VOWM+LPhBk7c
dgW6hqu4l0x4vec8C9Qy+B2Zm0Nx7kh91BmhAs5y1kq3CFvLnqyuZf8H/YP8ZbZOu4S//ZJC1Q+Q
I7XKYGfA3SESWwA2bxJq/xGfZjhTdysADwuSlSmfbU+l1uBqcjYYAZgfi9O/kiye1BMak4aLWVyr
0CVeZQ2pYD61+emPvI5UjwHyO5z/XFTWWG3tffWaCI767/7RN997GJAG57YUw+zGnq7ZqwbL5xti
UYrg/Fvv+eXBrkSZgeyng08UKpgjGu0xhMW3hd/muwCODmuZ6ltvssA/DuR8/FEfLsc65XgJcQ6v
J1KuKrTgq8QEM/aYdckSwRnwVWowy24g49BuiAH/SYyQnYo4SiTntYjVWSa+FKwDwkqv8ZDOy6X9
JcfBhkkGIuqM7/RZSHVnqTP6Pnf/d3x7YgVZUQXOyEh44l/5BNTMxjd82VGuA6uRjMerODSxLRz7
frnlgy9hTzHngiooGLZeisW/V7iNnbAXFJjvW288/TMdA7AtN7sUk3mTlWshFd0fp0P+WiW4cdGi
Nohj+xDTEhb28FzQUpyRlAewpMd0c9zNve34YOFBTKYL4Owz/SS6ixyPpZyftL6cn6G6J/wlmxwx
BZrWA8ELDfIcKgB6fDH5Dn6VtIwPr+HWaJ9W2CkjO+0kzNExHv9P2GjIQxA4/GEftaImVabkAsQc
4Vgp2OkSFI0rdzlD3PIfvgRsDLcFR98u5TIGB/Y7HfF7e9RIm7iG8BVV+6HS+RD8amkkrDbPAY0n
E2Xrqp2RQFKdo4miva702/Bz9DTCi07q4TXutr8ZdvuF/lxBRDmdLjHaQNrYwDXiayCcdg3LINYM
Nn389fVwoSCoQYn+WeLcsMpptDtWAzkNQUf/31Ko6JPfLFjBv8pLKiOjWDUXC3nGEqryyerTuZD7
YVYe6UWf9ntEuEIbkCYEZjhGXJQVwK6U4H2Qq+/wIG+iM3sdOI3ZzRQy6k3n9yAuNo0zoLisj+d8
JtRgOdAu2vZH0aGDZFDwJ3TpcUW+ozRi7KwyEVLJfTR4DuISlo2hSMd5sMbPKAi2WHl9hS8nmdKl
c3Xc+lOt9cTwEd4ufhE4uKHx6gXe1zXDzMk8Fk7k+09bVJY3eDdxJhVgG7CAwFmCQpc01oBH4EoP
TbnEK9S+aKpruHx4kxxlstc8JKXuYaXhdkdh+1QR8sVyzO9+C5JsS5K49EIMUsZkgrJTuYWCCce/
CVw6rOLMjB7TkVEFYacYXv91pZz0qCRoZx63/CVaZphJPYr2zhK3mck77mJLga1xNz5NvXZaY/QZ
e8FhrpUI6abdnyiXZfWeWfwaogGji7ZRl96ObD9FM80VXYKHiBVbyXjedobmWRt+dFfbqSVm5EuY
b+5semQY9INQaRd7UaQTG29b4eVmZJNoWapzJgqKdczWuztAZTooSI3aLqFWZq4k5OsO1pixCfu9
/3tOJ+3NsbrE8aHLDAbva85lCOQFi1T2dRElfOVgISkhEyWULsV9mNGZTOnJ6HV1hiDrqpBxSNkA
vs5Nanw2lMbzvL5LTHKyBIpzek9/bCnZQVt2duNxZCWAuM6ciA1154su/ElKpDhTdqS3NTtmMY3Z
Z7c7M14bW6+vACFOQ2+9o2SV/exEC35WkUchTG3xTbprHebztkLgikeqY6qHrxSlIkBJa7EudsfS
Hn9uDRIsfwNwispam1GDzH8mw9bJuGZZmFjn4sMOl6cBliir3gJGM2exle1+X5QJvTvnkb/C0rRh
Hy/8MTVTCT8AQPDAr9hIdsUZRDtqqO+LFzrzHya9Hpd6SKZZeYuj9anRLOY0iQ+ankNPY/a5LmrW
DPdV0C9bD641wKNnzjvh1pQrsLZu6KC5PLsabh8HgU8b/xQqhcW+vkFUWzoEt2UVheUDOrFZlYAu
r7XwFFHdZMfNPka+oNShtRZlHQ6BZGLc4jqR9vM++yiDszqvVcimxFRwgLqUbzGOu02V0o9Gy/gS
GTKcXFtJChc21/YTyE+HVP55TBbPXamInuXBhCoML1BdNRNRklupomP+1Eibt+uLKf1E40MJTDXU
lR4X/VjmJeteqoAREgoW6xSH3U57uP8L3aAKIIg+cZD1R/5IC44B7B0IgFUUmwzT5Os84CQd8D4i
WmdJLIFdKmj48HNcpuEyxwsS9nZEomC7CN+NpQ05fP9RyGum4WJOzmtR+xe9z9Ar4xn5yXU8Dl+L
SIlwpxJa9Z7MzhXk/OP0YhXxeaJKg7GRrZmAL81EYzt0f21vVf8tzNBbH3JHwecSM2KvbvDh0N2P
O7DLVB2YXWOp6bBro77FzVyhU1l8x7uf+QRLo5IbMkMG3vRECgHS0Y8AKxBzETC0nWk1rfvCl8ZD
fLXflSM3ggblY/ctql1Xg+whTgrgHGRaM9DTPhd42YP/0OS9nQoxZEbiGXo9yTdBzYWsc89B6wDK
f7Q4aep0A4BRIzDx580yCINlSae4WTZy3F2J964eqnINU3aPVkYwUnL+8lsxNmCmV9vEi5U+XU5W
plnl51JGR4pcUImDp342I/G1ccu6QAkBH/hGVNEP6UtXjWJh8BEo3o1jZTI24SnaTuboSVtNKJCv
mlPShIpmr2Ags5h/JjPnWIu+sLdy2Lz9Vi+yRTO1Te6Yyofulr+Cd2sarrgvlkOmBp9f1fu1IL1V
U1IU5hzANWnUk7w5rOQK5UObS6l7Px2tYkHX6vOuI83V4zNljftj86ZWH1JSoYtBm/sSE8UkcUIT
fCkBiDrc/xmLQTs9pyACYDesMz6YValeTPDCjEgad13lsk8VEww/gpdS3G+gcOQel2eSr8IlfyPT
uxG0MjJbPQpixpev1sTzixTlq+7OSToJreR3wkcwqiLBqzX+YdNYVe4xLkZdqCN7NkohtImU0/ch
w7q/P7HpdLOK8Pl6ZITNXirBT8NVgYLRxpjhBOGRRNQlsTnOKgt9uLx2AVviGylBwQo6fEwWn7Fk
5uDLw210e5Xsxghsw++0bnwvDyhJFra7J1XBXX0RcvSEXHVYwNSGm4PW/Efc8rWTMtkvLfIr7v7g
Ve4r+phHSkPktAhPtVOmiXaDxpO8mRCnQVph2wLSlqgBXRD9DcRRmEVUtnm1fUcpXtoWVBQMy6LU
Sg+HogaC2MHgEpR9BQSClbDzC4u7cx+631Mn12LzV3xiQ+rPGEjBVAMZou8H+Vmd189685Ccv2HU
92QSWSLdy8D4dHwnyjQcGnPMDGK/krzO0OVSyy5VJK2W9u3s+uzcX6DSJJyuDOKtz/A7vYEV39Mu
cJAtq3EbvYHFDaVsnb4KoSPSdPerkkvrKYJmDRreH8EqEvcR5EsdP2ai9oAMZzwWi0emvyMr3Ym8
2OTBpJS4IpDGDWlbqYRTG+kEJpMVfL1Cb9GzSjiiUOhruXQ7J5u2RGk5JguwKXud+qMB+6/GgTdQ
3PJA7EAkrnusYNakKvX2ulLxihJ8qgDeQkqNrWaoHk1Dyd/0hb2rg4cM55QDQ0IzKOgndvuD5ngj
Z7jK5C29oWQ0zfxsupqEEE++6ZUiAqcm3WaZhC48TFEjLICNbrkOdlmQhwQdAA/VPjDkaSihS5eY
wtVdpmqPOZFrsyxSzR/xVF55/xOLBKrq1fklyBkh7fdZV6U6aBfp8coRWXSkBClYjNiGHw1MWSFs
rLk+c8NpXuQhjDc4kCJJCl1cIlmUdDU65GN9sqqSDw674nSXQBNUZ0/w659Kv0l9+IoUF6HHWOvm
K2c4XaJw3pvlZMvCLG1Mx7a24UwY501qKawp6J1+t0tr4zJ2BFQWDn3MLdRJxrpOH8lBxYgQPkLR
mlyxZpSZtZnFTrDO9LcoKVy8GNMupBrwF03i7PM6gRvEWGtoUwwUBRzbQDIZ/XmOQtIZrydiaEHG
cipS3MRZqHF9NmyGKknCsUP3X5BMPafrGMJQMeGn57p9rbKsXK96zkcZT/WS6LnG+gkfiSTz05xT
b1gtU3IY0dZxZpOIkqxDYSNiNPOn4eaS/AtOI4ppYb8QtJLx2I7rXWZx55PTsdptUC152kRzq8QY
U1YxhIyDqJXZy5TedQAiOk5j56nql1YaD4PKjePRaQLt6AJ09NDzHN2NP7u73ldD+7NrkkWNbnu+
vWijs+WJbAkIgqGibToZj/oqTYGgCpGmGATn5p8OeG8tLHjwel4gyr1kaiZbaiU1Hpbv0EVRb/XP
BT+SmEctEigRkjfU+l+wrFuEf5nXM6k9abIc38eByYsPfBuclxJD2W+Aycv/Kjrc5Rpee6faushr
+wfH/t9WlspBHQGEPpq9xlvKArr5cSoUjOozRUXoFsG6RXed4SebyLSBSJ0llnVcTERsnDP0Jf4h
cEFaW/wTSo3mn+JkrgeRl7rM2ke/xPllsMRuYkLeddKdcix8R4QC50Ls1b8m2RwhXpSgOFCo123v
BopF0SR3GFmWPL8KdHak6Wm612MFY2xDSsuzjUrThdGlUCUIP7TZ0XQt4tSaBgCMI/TjyBA6e7tc
UQlwvTmd06TIUJV0QXOLlKlKhtaNALYMfqS8VcmhsEt/Gwj5yg04Bm/mGWeZWcHRiUa3DXew9Emy
k9r4ygZNuMBudRpNI6zLjsGjQfutuzo4bvp035bI3LQmvE+10D3x98p1TsbqNcDeXbL8n8j0Gj4M
M+PSsNr9USocN6BXXhHYGb9VLyWU4GJj1mFDTL67Ga/dK59J71acbWXTYWine02xZM88szenQIEp
EZUOMq5quCYZENT8SQ49J5pylskAerC0uBBcAx78GrUZeqqydwLW54aiyLWFmwBxouoB+Yyef9fg
3kxi4JaVbLJ3T86R+tlj6nLH2DCVn8xCNyyB0z/jfMPzBA/hMB2AgGCxweGrGHHT9+rj8Rz39bf4
aaf4uuQjKAF/Hyr4xZt9hsnBlJSCUmaBYyI9Lvcr82LP+3lRrZ9f+YjDJmU6H+kDI5rY+JNtimG/
1LdeT7hPXb13CIhWHshjDhYW1433I3mDXWxQ5tKRjgU2UA7mcE2Q5hf5VHsVJrw0uddgF3UbY/hG
AkoJJZprbkcqjwkLqeAxIB38WTStz9QTMXnhX1IufB6yMVOFSuaGP6G8/dpfnpNbV4v1CbaXuLlt
j5xB4n4Brs/1lUVexSEgyDB3HrmhpGtuajUBw9kOrPRLAiOgh6JwYRiErdcOgDG5WpeKZtqui24l
X+PqIQ2Nj/ABP5sIH7mPtGjJc4mieBu7is7Gcj25IUy+Wn+VmBBlgFQE3WqI8a+4mR3uLm97a2lI
QyUTpzNxC+iRvYlNQj41ErSqKlLfV/VuD12ENZxH0CMQFDt5uT4LO0cwJId7bP8bIHSQALuRRkQG
nHWk8ArF2/hfpk8kb8qBZvH0yq8EJUYvJnLUAbBwM2PQqKzrPnch4t4hbDi5gl1Q+icShC+EdI5R
ofZdsuqhV1OaXzIvwJB3PkOCjy61yrhxCx/VQ/jlzos6W/XWGcsV8C43REOvNr5TGpMwCaLDLT+o
lqgULVytbOTiomf/SE5YP/clGoNt/07eDBf6jA9E9LJ6vQ1cKhzdLyK/ipRNaOxZFhtUwZgaEGp2
IZ2U0oStHUtcnWGuaOssZCJmo/iCFoaibe7F1bc9R/L4fFPrueRi8fEniXBo4H+/R01EEezdojTv
yQygflekiRLajtaLvI+JXVbc5c9z9AiU51fSmnG/whZ+Ov3ncGe53XFeqzM0ur1jun/BYdbNwCND
WA87boNMfyLgFpuG2HFK/oNzPzf9vYsDVeGTuBg1wyirEuoiU22aZrvRGvDHhEgOFAhrKMVAOovY
5jbl3YWff8VVfRX/cHyd5hqIYFnZF4WRKxFTwuhIkSNootZXwIywNFdVKY+ie6ydNSEqYMH2W+oD
QMV3fumr0LKVpZjmOegJZh6lkZsUvyv6xeO8KdIrDwuuKmGL2WtO8Efq15XjZ6iO0eabzbUotZF2
YoKAjGQXRM6a/zRxbkurttkg3JXgthAaXIcbissLhLOh68dl2apoEy1Fasem7rgh13qjKjplG5bY
O3LAbSnHTnHG9wRmhY9ryhbL8wEX5VYghEaTqe89iVj0ZxyO/jX86F5zVHxyqwR4ufUIJXccBtrk
NklHTzPWBANbXa4xZ85GKDmnhOfwGfG4co5wsb2RUMlrSHKQpD/5LxDAwHix/59XYtpi9zqkezGG
zG2ETewh9Ghuha88fNRV8WjHjHTM4X7tAyIGUWCcULIBqHbtjLj6TU/g5RjoD86LmgZXLQh48BiQ
runShpRJZ89r6o3cJtWQnBaK5nhhf6vwMCZzQfLoiF1gz8sNtZGpEU23GxYXkf8HB98NrOcAut/E
D8jzhof7TJ1gHWcrzHXMU6O3ASOkFch/l85G+zcECZOyHZIGQwbnjkYk1Bg25ogb5zOHZiP60qpv
l9g+mZCmTvvcCYJZsPB7ToUSrwcFGzy/ss45KmxR8ExUInsB6DIwGNbPqDQYG84lmkZXePWZMtZH
tZCLPuQ0DW3UzaUmtW4UNS/Jk5+Ccqp0dZPcmeIoJYUiMKcLSA/Dt4EP4rv3FUBeLMcj//7aUx4X
RTRt8wSBb0u8A9i8zso6KbHHmLfEh0UvZ0wTWIY5WbhAWzh3Ea32G6JXmOtOUoVFXkgbfgIqnSQw
w6GmR4Uh80Fn6ifw82cDnMtqQq8URetRgTHZfZwD/KWcc5F/3mbtDeYfntySrSOUd3+XoTV2c2Ev
n3XzYTyCNBfSjwdG6bIw6dsR940q5xJzdZsi9Qmu0e/ubP7qIyn9A6Y56BpKtz5CzBoeM0Pzm3mZ
XwOKgnFiR8brIP8pcxxBfvmuBwIPgu1zLayopXmnyNNp0yHaWsyeSL71imrzgHTZzAoHmB2/OsOY
c08CfNSWdCcow33KUpj8A9Wan5nUv5eWsW+/8gyGS0CkuNlgFmmlGAnbjOmqnlrAaUZfAdTYHVOj
7iLu/m9xVaVfcW+14Ga+fePeLB+MYvfE0KH8m9dsBKB9fpxybHqVw0sTPDE9t55LuJRvzMWmgoYb
nohx4BbFcrTJwJGB6RKrx1ZDuk39g9aKB+gWf9JYnE2cmDFrd43ukuPJ2cadGLkctyU/ix7x4hns
TtD2M+OnLu7juqSj2sH1w5Up8ZW/CvVsj2T/C9u6VosXUyq2EMEXvyH0bTY1iorWsli2U9r43BMU
Odes4CMFl1K19f9S6mNi+BkbsiU3cKFe19OHpGgzwwi1E2Xslvfd9KbrBcmiMQg9ZQ+CGaftnhts
Dape/nJ6V2gugV7ouEhlv+gqgr3tzHY+mc/iDuQL6JFuWWRizp8y6ZchIrGGHavOaUMcE0I1Fgpc
RzvUYPT2xwdbI7vYdpxYzSwabZDptoAhvBA/ruaYHbgYJZG6ECoanO2EpEjnoRts8hzUFqEymAbT
rRk940lL/ZzeS1eSmUQiYJgDGqYd1dNhsHtOq4Z4JxNlm0VIkhH1029lVdpb81ONsKrXUgFs3PFu
5QgSjevP0KC7+RYyKOB1SZvuuDE/fS7e/1EAkmp4gcCNqApy3qGvumgulNZEh1Jt+zJcdzoOkQ76
fFhKpPerZkjeBmwc0kaw1O2He5shvGugVTs07WZfvvYk5eTRfA6USo9YDpNGXjJo/vk+Vw5OX0ez
cQIhpU1Q47fzroV1U58Ru7oaSUgyayK5RiZW0xl8ZGKFuZhqcofJHicnLGUQsfGtFJ5fP+7XSab9
u8RHYDD6XVhlMLv8BkOZby7FhHk/06tuvjFNB68r5+YZ2HSkDz2YXg0FJ89fMlm5glxw2FBsFoFa
ckh+bhXNvFQHm9UZXX8IidM29Dn4HKQ9RaaRxFhcoTotGf6em6/4KI6DSLBGvXwy5G9HvbhK2o4/
HU9vaQClxkke1EjOvR+0GfluWejrFceJ0BqL4aK7BwtpmNsBrKyTlRuj0MwPJ8qvWXjZel9eZTBO
wtVQeAT1IQeoxoOSZssDM0sSnAqrdLGzW/NCCwhAbUTPrDgiPWiNBR18wTXlO14LGlH+LYypiqz7
FpPA3l9bWNm1uCp1WVIsFUgZx+IFSRlaJI+SbSesHGHW6bDUg4QA2I5FlJostzd3pJMhiOQ4qQ+Q
nAsM8J5XYV3zKSjnP1tMI/hOLjWNDMFxAl2XkiP1fkKyF7YJnfEBRG0RsgNESgZmarP0MwgTgTDg
LM3tEucDN4bDWUtwVfg+JIxGL++kYrVIFqic284n4gsiGJuGOTPdT95QM6acoXyENs1ecTZA7BgZ
ZO/vPWPHNKF4nrGX0ERNOmkUZ1pPVRk4+zjcBHLiWGfXC1ZfWTt9N/cgQHJ3YBkYV+5DXT6jMBcf
El1CUdoWwI52M8Np0+NTiYwsf2/L7gd5bIZaN9m1DHZWFcTPmoRkTlgUHmu/LNyGHerCiK7Eg5UZ
t4WOiUPTiEmYNrWVaWa1lzAdPOC0aOcv6+dYegnVNeQ1eASRy6RknZeq68QM3wsjDqfiM/FsJpGG
RwU4hmQ9r3nWXS8aket6KaV/t40RStr8jWwUDpUblN/feZ6Vz8dyR0QQHjWLv4kfe4kw0ioWxB9d
6tx5+PIxFUi6iHKUjLFOJHfgVylPc/vGHZ8zz75H7H0JJgeWF/3xBUfwsyPkggggAx1xXC7DQf6K
wSYTL7eFNgDPrZ40fedfS5v0vR5+OyMjljByl3jgFCYH45GsFjtt85vwn+2zS8zlNy2HGhvLrXKc
/kVyJUPVkblh0bCUGXNxGa5wZNvOmPbHj5dZ6M9QvwvsLX5rthYl5A75vrffOVGxJ245AA65Ukjc
uUIdtqVolDTwEO40dKYPXClYogtlf2nweYyRJ4jn6pUmqMj9ZtAUNhR8QrOlM2daN2gqSgSdSXto
zQGKtYEhGdNpsPE3hmHXnod2/0VvZImy1RqZth/ayswdu8MdPoiH/fmfOvW27sugL8zbJFnnw7f8
vFv82SxOBKlzmpiFiLo38eEkVKBvCsIUEbLbB3sx7JoC743qIMNE6bD//Ft8klW2s9gHbeoSAI6+
mpHerRxUw+l5DzH1D+FkEIsuZp0E9iT1fRmvSLWqwxkVBQ4oj2mOvb25C4JSabS9ywk4FGHjP83D
99uegcfrJ73fiTm5Ns43uzNqbVEH35Xpfv9CagGnWdytD6ezoyC3V3wnDwwDifmWJbd6yCOlAnIj
8gPeCsDJS6ArlzlnbIiZwf4d6rTBWeEECUffEa6zsc17y3F/VrKYi2mZY5BxZnWUawVlmDqI6eEc
jzBqQKxv8RoDYsU/Qn3o7zp8j73al+WvoIpfvrv5YJfVGDzV9XloY9IgjdREEmw7o+/adO9/ibKR
kiHkVshtnwKTnm5lOuAW+drMJtD9A7MUe2lMVdYWKYuHv2YVLmyU6/nYL5bWZBkxz4arojjl5aE3
rpuoCNpVyN9Z189O+ETvkjrHVsT9dQyhJF8Jjx1RlNCdHHDdR3qynu+4ackZqISJOTvq6S7azW0i
Zx+7YS9QOBDTETe6yaWIOefDtHZuAbno7PSSXoZI4rem4YH54hGJehPf/JXeVOdF5h35lhmjNwR7
Bd1Sh01efAsXMYcplXyPUr/rBr/dTr5N3npY0RLfk5CmQz9K27x5yMTCFo0V4y1PzFgEcdy+dQbK
vVjTaSVHAhEu2ltDCeVCX/9mRgSS2vyGo5n9DcVamlELP0/pTELepH6Z/igGbte0LQcnFs18mZ3+
clhG5xx0HjZStlIn51k2w1KgY0Vae48I8KDSMEPwJpnEXmx5lzP/L9WmgznqBnXYDZt02++29AFM
hQN4GFPJcwALIKx/GJm15HHDnx8YHzn55Ld51G3zX9A1jai6RqEGLT9CO4eF7hhKhbCv9SoFLOLO
jJzNgnLVthzbevH9Ki8xS+ZUcWDs9LK1ttJVlPNumHUS2E1mhrcglBjMEcd37jqAck8n4YAd8a0I
aoYG/ruFBmQhHzSjDV0NgS77aKN+RqAh262Ay5D6to/6SMJ5EKPFo9sUDY58JHp5/y5vsPoTadmK
RiA+xe23uptnWV9T6NYgxUuqWPV0R4f6C5N9octuvlSTIJFG1KK4BRkcQsEhBYV//cH6iBFwdSfA
9PE7r6hA9ao9blcqMhtJebWfiRJhRs2wAaCw3h/6QonX1SWxET13u8bXWygYXl2eR3Uyj2wRqULq
6Aki1YGqowXoC2rHUbhU+yH25eSEWD6MP/rAfuMETmQfzpPswOQoHs+0tnKW+0cj8VFwdqR7YcGc
jX0X8PhDL0ewpKYxdNR9KJJ3iz5aAQjNQlR9ulkP3QZg14CIe/tCsCyhTaNkncc51QrX9R4r4ghG
4xW/ILWU5GKRl6NDrrfd1AXB4XIpKrRwEJzU1kVbbJ1hXfVSs+vRK6L1rgMA4K7hfvny/Kkn69HW
6n2OaEScLmXpuE8hEon8dRTY7kCREXSfcDXly8ql72aL4VObHdEmrlnoKwNuJ2yQfX9MLYbKaKsK
iXJ3cVg6hhqiOMldboQilN1LgWbEheqHHqMxjSF/0av8AaSMH+38Gy5XzDo/377/+R7pPNEuz1ry
o/J2HAQ3peYRfjOEms1aBwqQFDRNqSnCVbyD1HjpDtElYiG46WP4qP9dW7y2yO7hKechoTfrj3qG
09IecDm+GEW4eQ0qDfSdJaFlzhXmWi5KcF7dzgU0Bt6EsBl6gsBClL+v9b119e79CbGJFeeB8SUN
O3oD3dgXLixl/kXJjnbXK+clyHt+FsdilNs579Y5ueUv4qZ5wAtcz4Z6cnhSaFcBYF3lj1jTu2Sq
0nuHrO3OZRfXFhyaN2fojdFKTvB74U6Qqz/p0ooeDAm/zjJAFnpZzIwdU4bqAbfTQwJX9R/0XMqS
DAG5pysALN8Ub6g8dMhUQBljb5i2ppIQU4Ik+1COAtvA6Q0KC1jrNWfvvmiinxzdaPTpkEdIzHQP
PRpCLA9AF9/3SXPrbgsdplJCpDwl3QDjl4pfe7KDt5XPXhmPt9VWi0RHhdWpf0n/v6d23Ya9HiMV
WVykf75p1P3yyQ63tup2/87vPNoTuHtw+N6muyGi0VI5zqn2sJ65qcHhWiW96HzwG6Td5UOFBI3E
hXRJLUpUuftc1nDpc/jFIkIzMyILI96P90nq0O9GVyyxb6uM16HCOeWdGq2JK6tqCv7YMLlSS9YN
7oYTmh5sdPfPUQtzfe9QUBR5aJLjtZ/ciqE2u9R9Axwz76dtNjOFIv0MYpO8H7snJHX3NjirX/9S
YrrgT7ozOeVNo2UHRXKQHpBKf4Sv/dbai2Nqu1i3jgcT06ji0Rm3opZcU2G0T0RyiIbX/rrIUsko
uqpjN0Bua18GJInZgI4pPDsy8eWqXdaFZfKi4E9wSvLDy7pHsLe+vifRp+Z/lg3G03yFbx8Q3Eyq
z8StSxImiqw2oJG0jQoLrAX1ULZNrDv1m3h8pU7HCY+XM2e8GiFG+S6rSh8ZEn1/8H/33zkg4XFv
9yfkI2JxGu/wqnfCPg6KaiNunqSLNIg50b0lCdVjHk1ikVk0pCBVvTCQBWK6a8f3E/PswoY8xMjb
Jwy7fPbzXgrxRYD8FuOLX2+yxpBdu71u9QKZ1IZHZWd9YNQ1EH13TL0v4K+075EyGUI9hP4elfS/
0aeU5GjUYH7okLytFYDoetZhDU5FtsTKKJjEi2KB3VudNtKXaCdmYq5EW2pcmnJDiVZ9i0MO50Ve
Hz9SLbfaj1jnbM8dlOQ1KrfT7u+6Qn9bopyghfUgDQ9gMHpV9IEoj1X3p6Z5viB4RBeljOj4Hxts
wQPlCFUW/MSxf9mMD8CE9zgo17VNTANGZ5ndxYJgODU2H8+R55m2DDabrvhCOU1Lkds2d69DwWEY
eJ7G3n248l3HSqUFcoj6qYJN+JezHcL3AOf8xkRkxGmSlgyU0kOnlWvXKOigMK6c4tUc0jhgnQDE
sLfzz6zXUl28U34wxQpo+t8ylNSGo/OH4n1vXT4R7hRupbRgkc+GZcoVPakJzQG98cUjbwGTn3u7
GzcveiA/vtU1z34lDpuHCFcpGALFg6lB8YiGfb8RMJVDhPeMraZlIr7FJa7O3I16fsUKSwqXByIx
6IQMH6T+WP8R31o7HZqu/sBpJMJofippGqnjfG05K20BtUclGvUehhtB3bsgXN4D2airi7qmKoA1
+YfDMB4zcYMxZ2TjHYXV9//00J0kDXyjdGFvr0Fs1OWmPX9LLK/h8aMWMc1UyVsGA6RoitxbXoo/
XkBbAw94iG2LTfYjml+29A3xnz7EeN2KQ7+kVWutOB1/Yte4evepd2kaqhoqt5EEZunwnmlH5OMf
WbDA7BxBToOFPqyIFhKyEjaee/Ih5Y9iZhgYjpVUyHTlh5nYFQcjZcc5/Al9dPjaBma2zeom39Sq
CSQ5VIMld1cOMjvXBMOF7+XSzuD4tQgJLuDbhcldK1sFoSSqcV97/jQtG0nshgaJfMZgNfl1XyRw
dFyTxM82bxYYqVPfn8T/cRuAwklOz1CzRAxYr/XCwj/GLOy6oMEVpbv9Yf8VB9B1h4ok4M1GP9YU
mEP08UHk25hCm3FN6BoLZymsHZO31pzcsyqv2cNOd2j8zOUnSx2dZQXLioamNDRGrTFJ+HKo4IRX
aDFHTr5/iYx/Z8vf8BiEo/gnAIzIUOzLB3s5ScCTwuiPKKj94TiuxvGcO5oXRVhORdCuPC18gi4b
bESbLjL5zRNMg6TQ/b07BKuR8SeXwKnke7qKDd4wnKROTmokK1Vq6HML/b6SIftuD3QkioXnUjNa
Ge+KUDFUup8rqC5HFRaRpH7odt2TR+OrJBHUo6fmnYehSNWwtTb164eADHGWuFCyhjui+gtWIC+Q
z5h1Uc0bOh/YEHfJyYd9WE79aFg7pzeT6spROyBEWc8RvOYZrhJev9zJyWuQaVQE7ocb9CsgSNiS
OAe95BP1KP+XUluMoty/ufPsckRS3YT7LkW7NOxoLxNb/LcVtd4+6EOL5+cM04aRwu8hfy7rjPJY
DDiy++ZS7DLfCh5i/0xb6ZLdXs1IUxVyg+3YbJ7MPJ0V71iOzfVM9SUyB7AzE1qLIgOtlpKJg33V
1kTz5pSLZGTKtv7o2KQYBghoDvjTtNCQYlsuyGx5O76KU0RZa7GuhvfoIckxGcNfZ6eC2arebIKA
cqJkmRqlqwQ9hlpbSrT+boNT9TprrozU2J6TrEqXCXIw7E1upZKMs5OOP27kLBF+7ut+NRdbTvW/
KCu92dD8HZX56gCd7JBvKrDfC9Q0nk9AMu3zoxFL3AXRWhO+dyVzDJbqneYdxry8bnGFbw7K6Rim
ZXJjniJMYfeihFDsgnS4yZA+Ksc+hECFpNE4nq+5UD39bVeqP5UsOsPvOIUZ9HJCl8BDM0eQuzix
VZW3r6yoyC9D//41auRHoxDQIPVqSl/oJP1SDJEElRkJ65mXRicI8uJ42UMW7xZdifW2F+WQ+unV
nZEUWXVMMAcZczBeFlWGoZjMUNDkpFHat0zDguPlt0hhev+DzMQcGW+crkcq5B71BRiCNcLkg8z1
zg9b0qFCD07VsTfc/+zadEEKADQaPts6BppozxK0BZk3/vO5xDkw0b4fpJynxizROQVwbTKqDDp+
mkq5D4Tlew0ElBgCIitWYEQK9Dv2noSFOrgKrsjakRVIVayJx+1Le5vyBiOIwNjXADzj2V2DNplo
Ljq4SZTnXLkDNKOmJFweZGfhTBV7tJiSMqDYOSAE7SD9kclCI0GB9SgknuXeqY7mPgUhSHCLzePR
ZHt0j7RjbE8dJ38QV4FvBoY0blEoSsGhitACOk6V+BCoQ6vtVsrgH141JxDcl3zPXTy8m4f+gEBd
NVKMZ9m2jkLX8SCzLUhIs7msqxr4v+SWC8E0i3uv1GbX9ziHhfUhYxq/aNiJbpFnK6+88BMM1IrQ
mH7gfag7di7BR0Gsm1Fv8PrRPTN8AOQNAUqD6fKWoxWOh6uR99tjbVeZeozRzhMrx+OnAENvdeYq
td65gfrC8238hg0GKHtJpeQig3TZkjCQa91+reG08waC04PxzzZBr4x7B/dkfMSbld4RBcS8Kcc6
enadlEmR9z+0GDq2slGDQwKYBL7h0QCI/4juMRO9wu91eJgMBzK2Srp0Czn9UEi3TF0lsLL7zIYn
YMPcNn1hwZ/EkgzWXte8OLrQW+XGlX86qY0iJwrttuhn5eab+N6JvxsLjeUG+V52D9L+WY++6GqG
hdzIZnUt0Q8XCkvLQrJWQeMq5JFMD3eKLu46KydyVmc8FqmOy4znMyC2e361vjJ4/rfnleCo/59q
2RoXyxqls2jdBZkIg0i5SBhhr+0AWSTLrgAKvNYo6wU0NWz54z3o4U+zg6mcm/7jSS5VZZQ4bNHP
Fmw7aX3Fe6uA2BJbkMLdANx1RiQtdxWYBUYu0JqiB/KlmRYCS98bne8Jrrl/fgtzX71mqyfWw1eN
ze6PhHQo4m9eS82JLt98Xb6DNs4fmW5nZhkV67fFvSNx25/kf5L8jBk9e+JbAsSLSEtzwAGeQPYB
eR7IOC/EAKDudo9kl9iO+kamzZyqu37U4PNZ7O5fgJ3fFeu0gyvLAAFn6twp8yqHFGFdeP5ZvKOK
JZbiKSaqow5bDGMD/lUTmagOCBIKRRvig5pLEIzp6NED09vkRrMP9ka+BeqS0az59zmSocWZg0Jl
wGE6CKm+xIYkTdd7Fx4FdtbFrbBEWOZBtXZC8tqoQ+h3j9PCUr3RQNV3k3cF3dSAYHP6r3EUkOYg
PAK7nNC2QUE5HLIaDYfWGqVP5sA5KQEH0t+K8JnuXsKFpKZgw5EFboHj7dai/r9vZ2dl3Zr8lZq2
P8r4ZoB3Xrm178P+eySWBkfHaEzKD8P8Jtw78vFv1CrjIrrbMnxP6/SSNkBcJtoDGkBrTIRgjGJv
qpeyTdek2pqmd8jVd3tC5g+wc4+N2PN+xe3Ol2BdDdQMVlJ4diQbDYbvyEru31nqbX3DxFyVAh3m
QBqfAyY0HKfBLJ2RJy8vwKZfCvWLT3jeoPpVGKeYJfOe8rAXmyDyQre80rF9FFhzcbfLfwehmWsr
zUlexALqv0jtBeB8Nr1z/QHA40TLQvdpMqli9PUaWFUA1yF2CHMFZwVlZEGuhDVrgggb/pQWc0gu
+IzQX3dMzh5TSLNfCUTZtyYdxqkeNClmwQUshxH1CGCYDsYXRQIzs/Yxd8ABmphnfNMa0he82Qlr
GQX6syckzR6u/JXzw4Z7SSIWBt51Lqhx/xwMwzuqFdXA7rx64rAjNup9+MmEY0H9vdskx/0qkvvk
rmWqSS6Oz+l0wgZm+kNo22xxhf4jo+DJgL9ItaOVZSVGyIjhwSPBgJ63yZz5CnhjgnK5ZvgZBNmg
RCLpvCNBALkebuMlCvHBNo9OafXb9Hqf0PjRtnxs8CpKrk3zM7whhkP2cJtP+M/ASZpcEBqybmiz
DIQhOgaFAy9ocvz9BHIbHV78NYthDgwYo1M58C83hry8LZtPmoI9A+xahQo3tpvQGs+yazXF2aLG
wd8VzvSdPEqxEhLvGnTX14fJgtGwIgMK/iA0/XI3oL9AEGkm9OXpBt1btPMiFFVjVOXVl4nbdzrY
4M3hOrDE0s4csjR9FvdZEM5UB/ltILYbmWH2h7sgN+NBgIa8SXwakPHJ9+rZcldlkTryVyjU4di2
cNImYMzwvrAi3y3Wl0xJaPiZPusHjcX6njR15KTlSufg0beCpHaBwSGeeQF1cd7VuZ+P+Afrosp2
Lt8UAskD+gTnase6kK3ruknNYcCZZVPg2FOdsWJNrZhSCZqj1CFOy69GoihgtagJdRYmz0qxK1kY
k35t35Yd0fc9Y7K2JYy5Me6WUk6Pgl+Wz/Rb1ubuFtR7e+Y14nBMBHXwyldEPCsaKNvGydjqBaxI
LVbv7kmyWAKwFCEdP4gZ+c2a8S1LmAXraw1XlFdGRqFVYkXJBm6DWUl0Ah9A4/AzzBreqsSIPqCk
lTlPPFdD6hWBLInHKg/SzaGZE1j7YxzE9x5sxpkFdUp80i1V8R9KYBKB7KZOL94Q4rlK+NN1AayV
RDYDhByDUKFivPvpWEjP6vywiV7N2OmU0Pccvi2cwwN1y3LbKVhhq9kfLe9U5t8udBWWFMzbIIr0
j4c2+efnNtyRzqmsNct6XKTs6C7tk0SyTLK10nadx6UKPMscKHmmjzNwf/Qu/nQjNGMJSAjvK7uY
7NM7KG9U1+zV5D9NNf1Pw51m57NQm+Fjnk0p24FbHikR37e4F7JrisU/vJdx/e9+gk9rtd5/wEIH
ajjG01+hSAk/RO+rAdEUL14eSkgaNlBd9lmDharCTXWEbM+RsdgXcR/dnbFKKZk9tBkKlp/5EmPs
mkby4x8IYWt4Q2W0oqXrwaN5YKGgR3OcgE5fnujmWiBr96ESAoz6LOQ31JKlAI+dsoMxN2R9on0y
p/3npvnnj1W7Ns/ZI+0Z53FscvvI/ROw+U+WVrNWwIYqjEmSa8jw7W20R7YZTPqXm3c3iF0NCvSh
GI921MeKx8LwEx6JkkVj/GZr4exDWgNKXQbwOnH/ZSvO6spOSMYw8gN0NAwIBNTykHyoSz100iWj
byN7BP/xCtigXgg+HskO0KNmuWh0UgEZENg27yp53zJXAU9VJzX2w5bzuZGyzUtScmLQJnXlhqlp
2StpldKskXgr8BQo2J4OZwZxSXeHl3jK5rxxQkM2Lzpp41TxCFow/6hCyQomCGRwSfcicxUXru8D
247iwyei4T0jEmrTu57mrFwVVlB42NFYZmDGyeaEfgu09LdNlMBHUii8XUpIlVGH3IqigG7CScSN
+zwcSCARcgCa4QQFMVvwFcZhYGV44yXHT5nhFquEQyKKNGzAsGJxIRqW50JojAa39FZqltXR/8Ex
Q14xKfIgO5Fxvw60jS1PMCSXRSPlzjvz/nDvg7QPuK1w2PGOHMtUtweSNiX6N1/dc1g4cJCtN7U8
HlIyjSGoatgknwwiDhZLju5x8JOOABSsUB5DtgVMO3envUoNN3SAtgOHeMUHuvQc0cBR1l7VZKxR
1BIOj9c7DEtTjk8I5kmVenrnLWqG1qinX7FReMChIjMn48pkosfs2+MrJQYBt+fouiDDJG93GyI9
LvPvy9KzN0cb6rEOylPD6NmcQzFtp7ShVgjK1ZFljOnG3o6/D+GEGONOf01ONRIYLzdtWSzCfWI0
dsAwKWdReauujcmkolvzBtPN2J+8bu0r7vY70zsdGL2AcrN2l7FzWaunLGM/7qXPpofSIBxH4ITK
7Z3yegONsnNJZT+bETcvKbcG6/aAKBZ5z8te4uAPSlZSNfeVAxi2H6staMcogAmLXzD8D5cGCDba
QGBYimTl+AOOu7NIEzjO9fWcivvQVqDSa0CPfv/nyopJPpoZp4JkuC+N4nyKyINSrZyL2LJkNqt2
A1635MU6KyS6h1SXlr44kYQJfWgMDZDlGjcaf+YnncfR2Yis9Ebz/Yc8yQ/FDSiYW7fzrYqoYq7s
4omKon4sS893JguPtSsIxPeeJRgtTF/3ka8sJodY+yQ4PKBiuGIRfuNd4CUNdil72SAo7MXHf16k
WnGmYC/VRXqc7X9WdRTXEtPt+qOeuDOdWaQRop++eEyuqttP/GVY9MUXErdFsfll9rLiw4UADUHL
0eRslF1outRruczCUfCPjmWYrRCz8leoILGZ58am7dqONWOPh5+RBAxh2v/i9ALHVs92FdlxEQNS
4jdzSyUC630CNuucAxcSQr9srrSGJHFaibhjpnNGUnU2wwFh77PtyNGYQY+yJQq5qAqZsFvXFPeE
b4o1ZErkd902WQ7HTqn6qLxy8tToqNQTGfoYUpcQDVh/xXrbEEUkkeHM9Tq1pj8VbnOnxyXoEZUX
zc+YPjF1eYH/0fQbOv8MtBkdY4DVGi5dVcvujK9Jm2G9oHdWnbXEHPUDKqr5oqxb91NAvFu2wZEk
30fYW0FoVmLcrL+8fbeXwgt4quRQYQMtUMV12uMlT1PA0KiR1wLVQ84YH3t/ecCpyMPCTPszt8CR
A0LRTNIcC4AcGli/9VORlA0RvCIqZvFWT8Z5lGbIkAcpFbykuscesj9RwY1n+cj9hZkPUNlKGkm2
iatnF3+7Anl+hwUGQ/msPEAnAHbNPs0pqjis12rCmH5IlBs28rcARzQf8mIVLR3t18p5LEWVDsF2
NlAWvPBfg3O2aXAnH/BbuIOMQ2yn/Na2h2b+XmPzkU4NGYLLBLBziOeYmn7VHXyu+GRNEKN2Lk/H
znNr+plm3Q9WNvubJKjX9n6gKKbyJU1BuCUki/ha6Wk3b6Y+6JqTTIOvlSWdk9suwfJUglLxTNAH
i0GlkzqDanYv79yZ+pTlReSXbWcaA6ReeMM5aC59HFO7uSVG9YEIr+kIR5x3g9TnbSV2JaPCuhTl
nbfCeYTSgulil4rSiPGH+hC6M2ThifH3TDLiWQ9iHwLbbLPnj0D7e4JjoTTSrZAoJT6dUTI1UiNb
P9TTc6hw7lPuD3oinzq3OzQiTr97C66kdLMc6V8+5MOl1Z9CR0GkbBXaxO0j6FMr+owYVsc+lbAr
i6JAbsHx5K+6zQq0Ia5hpWO140lYyhS2kRfwHrFwkzGDIc6gDSuj4+3mkQH/ox8V8WDx05X2B8Nb
Ai9ublzRuMoom8TzWOwLUm98UnQY+Gz/7pnb2JNOq26WSyocpdUOo/6o43j5wlkW3LP0iJIoU5lF
p7XnG9GTf2hUGX2oXfX/N64mn5ERMbmqBXueFSeIsngDf3bDtYnvbb3hEypjz0qEvspXo/aWfsjw
KDPQG0yr8yuhNawGn1mkktNMAlc1IStbOVt9sCZZF3hEPp5N+xs3esj0GYkH/7YQDWRqyQOvGluZ
J2OC2YZajlmvx87LpF72m8IrYz04Mr4PjZ/3T0q9+0szQ7JVxN0AQDx3YNWXd87zkTjM7RtpNF9u
BxMSQVB1+ceEPn97ioONVzmwYp7ZpydoUeIEIM2p5wT/w1ZE9TJhby0wF1lHtZTHppmKQ80VJE2n
8REPMnSjD+aB0wb2WCIX0zf23jlf+krs3ldSE0eDrLpL9Jn3lEoj034yB4Ez37tDevJppcM0nKBM
WVsVL0WWj+esbWq7xPUpfgM1fpmPTqdxIICHZFnGVluldapNfhgzLnOKXIpnvSsxPi7eKjilvCnH
bDj5wx6DJZES1b+xAUNOohCgcc9oeiEMTgOFRPcThXr4HJIvl1vPzEZfIBPVN4/kO/5hi08ZI6W9
R/o3Cy/E5MFbu6MhrpfaH146X8WB/AD6wLjtgN3BFQ+sS76klslw+7fOccR1iOg0rrqpxj8Bilbv
mIxLnKN+8vJOAvkddIiCBRJh1kOrAhfnI8UimOjDD9XNBJtz+gtWHOnoYN41trqL9g/8uRG3RojB
QW4iyrS9VNlbhXHnjF/2lHifI1oUtCkVvLLbTG5qyrIK60/N6QsGT0IHYFMuv6mSzNfgykeQ5eaP
wfw6dXvS5YGi8iVkvoDveZRscKB5tS8kP+gLrNv2dNA+UaQjQbaTgNhMXixqgfyA6wZcsKcAnbhR
yjxxp8osqYqaXuD2WPATMJMF0AQnJ6UEw4tHQVKIVK1pctefW42mx1JOuNpYG36UF/aAMeejpEWg
Q1JdD8tS9HYMEI5VPfkWdtV/AYmrEZfNiDOmx3BZh8Vsi5UyyOM01ZenTLjHdKNezvHqbPK/aGlD
c/dcziH+GAFJjlapAdwwtL93Y5GL4sW1TZs+hC1hnWCyOj+d7QxYqcYwWOBGp/T0LpChnOBEMJUo
MWS3IH3HXlvb0qWiFzNHe0rcQ6Y8PQ3qLB34wttpbNB7o9R3T7EkMeSYxPGJD4MtKhsYvCmwscvw
VBjuDRvfuarlQJNMMkaG9tGaEg0p+Vi92mbyqF9AQfRao3p4oXdPdqDyMOz/V8lnFlwFnJAdiu47
z2TCzIafIJ7xkastkllakNehROO0NvGTEh7hxmqaAGRPp0y3lDmaG59ESDP2dr5xyJyW7be51M4a
Pz9VPha/DHJiIGqBeeDVPzViWU9tfp792QIv9gWToQgRg8fh1hnpObYYgrPhANgKEXuD68m7S7OH
SiUQQsNhbpJUUCLVOD1n2PjRQCf4lN5wCV60zMaupkKARcucTsq63brBt8WnH2JcF6+BZM2mpj7U
FYmq8Wmh2P3wVY5Kwy0m6nLghSb3dhvjbHh8z2jEngwCNWx9c+byxo6uc/dZ5TTChgLLDVuF4LD0
2k49Mh4rEFiVRFLprc22CU3w9HZ3x5R3rab9d9k4eSvHBnU9fL6eRWa5NhUgOoVb4J5wdkAXrI/w
MY/YlcQnjJ6pcYZYAOAlE93TrjL/HhHc8E32Z8SJ8ko3SRa0zMhijwjcKsTYsb0mC4W0SKT4Mwsy
FzMR4Ns4EL45QcjvmCaT2o63iPAZEQpf82bqHIPrzDbfbkO9sDL9Tfi/GGdICkcgZjbtb0gOjNVy
mHv5wo9kNzp7A4ZslMzELm2xgK1t6o8G4qgoV6X6Dwq0jxJwDvLmzKLqGqOrN2gmp3217wy1uwXk
n1WP62hYQbiuQiJC7w4cyZJvrXSR14wXp7dNQOFP4LvFkgLug5OoxqtjIDVTYtoNzD/hw/1AK4LV
CG2L6gFAeF2DIS25lsYKQ0zNH1lkkOKTTsFnTsSOqJMPQInSDvaF6wUG4dkG5HqyAyENUbmJYgIu
mPIzbKLpKbeMf6wSLO6p2i1faEbkq3gl0THGkkj+lLCoW8FeX13/Mw+L6o5zUFuH1x2nt64wOZbq
aUAaz+hLcjfonLmnCmOI6jfaS3h/4banRsr+yvdp6+oIHzKlxBXXQeH+UwdBuWS6S6bKmCZOSD2v
uQcOmE0Vom6C+B5jf0qogiSPqOXeKIJURVbH6Q72KVGt/5QnpR2BxBq9LiMT+ThMNujyUca+U41h
b1wRzMST9uXi/c3t0/7TEezkeG6oj5qMOy6UIDFfAek1oaiPsMw4Eg/LCeQNLIEJszTYfBkCgwOq
55r0XBZyFrERsNJSLdukUmo4iMa1ZhMANB5jYXzocba7zijmcGnHaQKPFQuuxrVEDexRfuG4FuFs
gnvyJ+/EWzhTN+bcyzMj3QR4gdrOu6B1m06OkqTesCDpNTzoeZ1Gb7khzDuYPmTCM8Wtg6DUUs1P
kDfUGUXtUAFwyHhIhtwZwOkeF5m+IyD8c/lOK+DXJx4/CIl/NpzOfWFTqPx1BoPC2756Ra2JHKTn
UdvABN8SPkbDaotvEEIZCvQaLZFsP/Q3+Y2fg5rtIcQ09gimOaoTMIH0tn7/ezeqNDAAlSW9HOkg
s/UbdPPf0NwO7sMfgn1cdO4wn6JTiD1myMOOD6B8RjQJtCeIqCAQ6UADh1DbX2agQjshJYzeyELw
5bVbWaMRn+x4J6ZdYMidv3ERCsmD5KW+WOkn0wtn3sd+p++EqV/37tVAeOAoQpo9IrP+lc3JLNiq
E5vidvIciodq0zGT3Hf6vy2oJrvRjGi2QRwSWQmGtL/KYKgZjF/geGTV0RTgXZpq0P42BqaxdY6B
D1CME7UsWbU3JY2K5H7o7wcHF4lGpIMuzOHhxCZYol61tDnWZOqPbNL3B5GH8auvVmsCHRavFyKB
d0DNCj4TEd68fzFdFGkCo41oG4bDvC7It2RxPOwq0G77C/hLkLT9o6lEY/enPzgiIpwb2GrW8FKo
5NjdaKlGQ/KPywZkdAB2cLbZRrDG32gX3PtS7Mbs1hXXM5/DG9IrTnz4I0oA5FDJXu6tMFCqmn0F
me/Hjdq2WAezJ9vmesqQ3lisVf89sPFpvOxVXKT+/8wwDfGrqxZQ0g3n1/vxdr7STFTXpxo50xZr
DUdr9JCDqiK7tpoMm03rJEER+jNsjehIRtEMuAhYHi+PA83cn3Z3JetZVgZetJZsAVwQdp79Ouyi
C5BICH4hPOAt2/NyK3p5+aqiy/LCbSrjzGaJICWE4RmYn3R8rGjxsfWb3H0MLNz8yIgwD0mTALML
jnmdot7yVnO92cQdsXR4KqIQ6tySdBt75RKxJaMhFuWc4J2znBwXUp1zdSYTuzKkwTXyLE9UsRe3
v+XvllYRZ/w8ivuvLdVeaJB7ZbKSm2XyRuHwah6SZMz3tnTXR5huFtsSyQ78pdjhIjN1R40kykS+
EobKJP+7zOf5c85lN9XqTe9Mopnk6VhuGqflhpkE6OlUlfG18p726Mh1+J7qGNFAGGpJMO+PGuAb
N9bTe4Z/BK000jSvqH+7Oir31rHIcPqvafC6B55xf2VMJfjeC/382LgfkERlBVQfzyvJE04JmU+E
b6/R1YsCuzq7HxpfyTSIGki79PQw3nSCZMqdXxq98QC2XnPkAW32PsLwOyLjgtsDnmnBl6kj3vkN
F1Qk6QzQ3BW5kuCJyQDJoT7QsYtZfDU68WiUVjZhY6uwzMUQiEGsDds8tpyWjWpt1HvwAieyQWfP
SY5RUvK2RsETqnmbn1l1J7bzdrw57vhjV+D0wpY7SePtfW2xlhmzexCu2OxVMDsZBaSgUUs5tcPz
S6twlmDoAstYoVg/JA1Yj9/88x+A2QURrF2A+/hlO+pP5T68EnJXBnr/6WFyplfPqr0MJZmjNA33
VURbDgd87VJ14qmq3b8SABoMp4WqCS5AisVPz9fhc9zrSSkX0K/yFV32WenlUjZdz612Qrep3xXI
ox69Y0E4+/GnczKwPUDxHSXXmG7wytLW2zwiECUlGjeaIsiXxN0rU2AR4/hhY2OEwtp7MIZqLSor
bk2b31WdoK31hctiUicj31Jvo0tvSHQDNP0PYtECHgi3Zxia+2/AroXqa3n/sd8rlHBWUMP2A/UR
ITY0KXRkwirwXD0TFNtb4OHj/hIxt0cZqrdgoQVlWKDcGpLtawTzLWNQO6ge+v8yzb8AMuqjrHd3
5HKoZHq4ulx5c9zF8nnZ/fUJsOyT29iAvV713JV0bzgRhFdt/BySXwNlK4tn6hD75WRf1WHaAoLS
lzKOqy+KdFqet1MLmU5k6orP3UAIce35XLOEJvbcPsy7Y2b9VcaDp9whzfR0GzYVF0pQwnh58/3o
xNdM/bE15HKIGrKx+JfqlhaPFyveNagBI6w5EaoqB2ev32RkfigPMf4uwRjDljzpAOkIRTs37LD6
5vTrtrryIeE52ryKH50ykbW6vxAQk/J2bysNL5RnTNOTcQj5fX5VVdYKbkLsfoAbvMgV3CqTta8P
RozvaiC7nBuU8k6eUNxMock4xLC53Gd/QOwUKOfgnanGp96XRqS9WxybPTGDMxi5rUM5vVUkPVXx
LJpy/+DinB8PzJn1yfxMGabuKYkrMQSxV/D79+fWL6lr3HaIDjNH91cY9F3jDd8NX79TfQITZxne
BAWqI2iko9OV8qPUZLAtafk8gOnfsgw3Hvn1K4yKoBwdWHPdVfATl7E62b6B5/WCWdpnnUO7JQKm
NTdv+HxUJynbPB7xHsr4PniLc3/L4tO4s2zza3/106vYMW3nBX/KOotMMn8YAjxpJi/HjC2cauNQ
1gs52nHprn1ESPM4Nxdbonj/0zilh+mveEn+5LHkW5/NXFOtZQ/MefHVsZQZqiv5eE/57elbyNX0
7dfsYMLlya4PeIkmreG8gsUAAQpLMml4GPpMe5k4lxtw3HwnJCFQFwketwdOn2Qt8qxNKBNFqGYH
lvlNm9GIrB82wATD7ETEAH/LWvIbGXzcpPLi44tv6KtQbqrPJ5uLgJ0/QmFAojRc+2Vgnfx3cFSz
ZZYh2F0EqFZ7aAcojMfHx3uGft7fmm4rS0gZYET5wxLaJDjU0HPN7d9LxhcuQ0QbuIusycfa3m2f
+kXwNzJsKfmpX/d30t0jVVChYLUA/G0fUanlJge+zStXfDD6Nvlb1M1JuT0M+AVRaEV9WZeTd2bt
h31AYE0BTTOXRzgTPszisTwZpVOkawl1yqCJbk3ULu4p2BuxvTUp1d9ecIgRjg69I5hIpNi2ZnXE
DPtR3dmKYSaRIXAKB8WPiL8Zy6mysevLmTEbC4NgAhvAfUQ0642jLJN/emX9NHGxOfeR1iQOiIyw
v3YLSttcT5jGbOBF6wS5lmCgdrq1xYbExgtzgdQmkR75d8pU+u2sfipO9ZFcUgYQKX6QYsuSd7lH
PmJ4cs0ZxQv50YO4KKP8toUX4BzXTP4dHulSF9vwE/cHFxz8JCPN8vlA+EIfb9DEakyrb/dsUWfM
9YS5kIf9egcG9DizkFN7UIDYRRPkJQXa2TqLfrv/fatmByJrvakCttI2w4JUiIwNpfedCcBqfUDO
R9hfc1uD3X8mit7xxMzuXeaugLP1TU2/uXKwhxj9ZKSI55REXqI4Odg9fPGP2FgKUmHBiltYLxly
PpQKrPnQHDy67g+8DY+NIe3poAiGrMKEAeokRBl6NHifq7ngIQKc8QrrCJJJ5dDojkxNLo4oigb3
y0cKmxxrCin6RHMiQkacdVKX1Y6GJuf5kyVHmc/JnVRyIQTvuY/PgVKmhAY0a6boxxWIVIjty4J7
Lqkt9nHsX08awK3Yl0kJoj+R76StYDX8pVHk0dAoJmMrTE3v0WT04ogdZl4gf+Q8h+LYZNEeosM+
ZuUqBU7VtHIK9sz01wwrqIX8ezKXIV4/B9kHZUdSyw98gsdAqrZSbHhPKvAgX2dv0+LQjsmHmBj5
Eiea0cGKOvWHVtj8mQUJ/Sl/VyKvQfti+tdciZ1+/erxoBgSFLNtifK3MgnyF9LSRfdcx4kbPO5U
YY8LEyWWl7NXbZt8WP+T7gSpb7MyWi4004vMzyUi+SO1qAo0qeX3iB3JNgoKDcXhnnX0WJHxJ5z/
RKGKk+d+dAUjxwnwIL2kgtlJKs9ahtmJ2nxNnA==
`protect end_protected
