`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
G3hzAzj5NNov/IqtEWWAiWy5t/AR0VyHo/S+kwttsfB/NeWMrzC5pDAkXF9y+L0rBw9ZGZJeFYuK
KHr9ijWKLQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EkHpQkj+0xYbYgviyS6qvQ11ynnP8f89hC03Q0P8bxG9Z8UmL6wSEmhhkiXEcQBYAm9ABOhQL84H
jcrtwgYIe8U+u6fRO3x891o6FDppMSPTIUpqqeTocqmLlkMY5PqPLz10Rt2SPUkomQqSr/zPqi41
A92omHGFt6CRIglOhq8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iFcSr+MbAwH6GuNjs43t8xiN8avus+PbYq2NTGV3c0az73gTYDbMYA2LslIDsJxfjY1mv4hWPFs9
wKiWXKINec5c33nnupXgtM46G+z/60q3e+pJdtcaQuIC4nmf0rNGH8XTgYWJOts8PBNctIF2+7aD
80+XUOanW0j1HTsnvX7OLny6vCGap3X//2+vuiqqz6e/85txUsMCwvBmk5nrEGzVMkiMqrgZkkTs
8SiFt+n6+kUoscZ1dvd/qvtXkKaV6uH6OCVIwft6vBhyzaN+8pereWQqRKhP5pdURrM+7DcOlZ9b
CZk425UByit880+vsKDGKmUnTOf3p/WVBixZ7w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EqrZFY0ET8oR5BGI/slbIqZhNqPRv38CJP2sdRPQimH91g/dLlVjlTwNhqSWDCbS5N+gLh0XTkV0
RJHP+iOkI5oLaHO+JQlgLxbRTLyLOjGoc1j0d7f153hSX60u1EyE7OjdL49s9RM2oI20kOdRcDpf
m+10tIKM9mc9WQi+IR1tmeiL/4wjNjPe3d/m7d+NwQbwNBHVN3sLu5W1vlkTG7sLzx5ViuLJbxVI
MWYCg7Wc/Xkz0xKeZqrqikgVPtpWI1nZ1FwMVno1MymDslSx0fz1C2vuGUGft2a/h4E6OlxzZM4k
s04LWw1OzynZv1VwrasFIw0fzJKaiO61wFhJeg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HB6C1SPVefsT3FY9Ld7wyB8wrp59Xn8Wc/bH+XRmUp4gXXLexz0PEANBQ9R/Ldc9+8oIpTq9lYGJ
4YWsa9yqYC8h5jVcTWdyKt9LrI+SUagzZ0tYyiU2DEF8DGwv/a9W5DsfNLlGSsPXsnwnHauM03m/
q3OBSzjejyYdqsTDn0VVIpL+H/68wxVoQmI4qGCMnMSJYBuU46S7rPHGT75rVa3r5K1Rp8ara3se
5vNxuHIvfHaTHjNaxMEYw0uemTY3oWlZw3vFrg0AXhidBmaDtvA1DVPHKnAbCViac2/lwjmGCifq
moOvRET0ZTrli0r8TV7p/g09pakmrsp8KaFOWA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nCMfbA+wjeeX94bo6oWED5ln6VMsCcyObdQpsgmbzjAmeqlzgXcYdbJx15tDcvpKqiGOtP8CnfC7
Ni8vPSAmF738Yh+H7bLmNMRznm+NgRo9H5GGwLG1NOJa8Qx05Q++hAEbX+gUecX9bxCWyG04PjKQ
BmkStJWonJCWeJ44mVs=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
foEhLl9iChedxElF7DMZQnoUwLLUNYma6V7gK29F+oa/MqpE1PExQ8tm1Gq4WKVpky6U7428IMIn
J0crMpOfUqOuMWdf/dZ6xmaRKidQU1OCbOkls69o/auMUkbqCeAWV00lU3SDaV3gZ/d7MMZSl97p
fTNohr5lhYIZRuZ4ocWwoL52I4ASrmvqxKNjSEab7lvQUyExO1PHkiF+0bRk5D3pzJ+JlOmGFm7f
Y0NDSha1p1XEFgpt6dg4q4tBov2ACpUTr2/JcNb71xAmXp9Z4clB0/mb4eDo5edc3x6ctsGd1oEb
gGBG4gn0qrnK3RHvptZh0mdCLCnYRGQymLFe6A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175312)
`protect data_block
A97UqZbRjQ7FTZIp4ewix7kcCkxm4PgDfCk3/wLmZZPhAUhcdZokRE4AX1yk5zGmFb5mb2knJwgP
lLwZrMyL25yW0VCxZ3qZ1IVEKKPRCsaBtcEl50+oO+kN5bsFwW9Y+W/3mAnHIpZePxlP+u2ix3xh
MoMT+bRsmuni659SzN3l1REsm7TksQdnQrsb3ov5+3CrzJkPXksmfe1IDyn0imiNab2X6iAy+z4p
gUX4EqdTKhAIe82phH0bJngKDUMOiNSxp8xjaq8d2SrDxoa6akPQyFcQX2Swlls2eUWgXGgJtflH
RESwJ2muxEb8Wa6yQIBCfmWIe2HkrWZDtvg/NU4iVXFJAxCJPN0Lk3SdaFdrDj1zXdM7kS2Z9n0W
3kXvA/VHj1ywLdDjmjrFpj2T41030DmjJopcSTqkoZcOzPTcFOMVrZZsbz3DCBS7QQ6WtuJ0WjB3
P5v4Eoja7QzbdxqqPx3Nh9aqNe0fVMbvIvdrNo0eby4vEhoiVdR+ShSMeCQSGJSS+tDHqfpoHtJt
2ZbVyMS1FXpWTtFLl5apvI8dpuB9kNCiK1g+J/BN6osEyxkymQHk5lTmwrvkyzqWXlgEit4Odmdx
i52X0gS4x3e72cKbqJr9GkETQr9+tczWYDcHMoq//dab8zVYP+1Po/ZQ06Wxd5dUbNUUT3PbjpvC
L4pDOJ1hvLIL3JVfTDYrBUxPAOyWZVnEvaECOKKuRLsuZ0c34lQlm8tGzfJTLwD0z0ZoU2eoOjOv
l992CnZLjuvwWKiO9cIMkQZREd6Mm80htYP+vRkJqwPCiVpTNwwXkWG0ipM9LuQMV8/dB+xPpkOf
F+O835X+h4nkUAjELnYTTIGERT7ukGzZ42LdLWUHsojIWA0zB0jnN2jYyEN9Sz15eZfc05/+EFPa
bwBbS3qTAi3Vj3YUQppuj0wmllAZMmF9So8AKy5B/Q+LpFKK8ijEAodB2MDcgcORCASvDia7+fsz
oSHvVdPlDv8rUAZwTUgfTRVaFUD0Xt3FJUjB1Pkx+VryinhFC8kIv8/ZUb9ZyyL9tnu+cFV8HTUD
KId8x3O/poJZpshzTwhdglUT8KRjhC9bKMcTxzRWMloJeHY8j84mLSkicgoYOIEckL6QsVxoCSk5
cyRWt66OtcJMG0H6+t+8ABKmo2CbjXsmByVmeMhMGB/wVikia4yIYT2L7gFRu5sg8ZZm2fpZlB7U
f6NFSQgOwTNlWnojJVNyBSt1uFgFd88ijbalJWlsCyBvrOBdtyhSeEpMGF3UPLC7nft9YmNYg3tx
Vq6n1SRc4BsmzZen0rNifSQTpAoWp5z72cyCWsh1uRopLn+paO+DwPjpZV2lljOkkckLCbMilf3R
4xbc3kePu9y0u+XpcOBncSmaldV9dTVx0rD3YM4QcRyHoIJ2OHLUq5HmBeylH24agK5C67VKw+Pz
tJBulKfnqEcmeDrngOTO1Op4moD8RUp19DP/RQZCnFccXWVjgubxrzI0Ijb2WX9VAOFjoNNar1IW
UBDUKpEOocEPogyDvi/SkxcauJv7vLjktit5ofG+l+G8iRHXLhyScB7jwgaR3zSweMHQB356b12e
NCA0ApM8isWZEqLPCSfDi15rkmNfHbwaUQWKn+GCR0lI5/D0u+VOjCXBOt2My3l1/1ofhcTGVp1C
JOl+IS8FhJSaBV3DB4FUg1ZCkXqRtj4KLjp1b1injPKmAJ54My+BnU8DJ3sfC9Ojn0nv0pVGVRgE
DyQ8ne+YFL/IrteJBMfVVHcuWZxbTIVue0v3EITAtIfHa1mwLhQ5WQ/WXt/rn7/ndTesJ/p236o7
kIEgT32tWfnYZlX7sLbBawcOKQWtdLhHtUvPah+G+ISNLAKmDGdLRqXCisrI0ofArh7fx9XAIbG2
+aZpnYYVDSZgiBZiHVHGfVzPRlw6FtIraDGOf26xBk3kL3g96oPE8MooKyQRRwXOII8HcXD0Ay6g
YroFoRV1VFO1wBBLZuqfgM0higDk4eUshbB7zBqH8pVwKr8/VNrvpFAZUFWw5kY+bQ/ASWx8gglt
xgasBW7rE+f12Bgk9ioxlzddexDtiUu0tPn9UFI9D3ayw2zgPacxrFP7K5DVi1SObDmJY4AEYtN8
vytDhOSDm+E5wlZe1gKS4J/nMddYSJRbvvuqsLs6l35rNe7zKBriwke6kFe29cWEh1QVsLjkIxJd
fJL7Qj8uEnXG+SEPKwyZ5PihM4FBH3TfBVMj8nLc1jUMduyMeO7/hMGhhh4RtLxD/w9Y2mIgatnd
x4HKOiGjqMkxr7MrCD9784kx9aC8GmdgcymWMmSlrNf8LUpkW2+YwgAe7nAjn/kNBuKp+p/R3uh2
VdtvxcRSBeYE8K08IqZirtWcUv9pY+l2+Qdf1/KzEN0bt9ZuaQ1m7g+8rdSAr3hO17w9x+e8Xq/3
2jVlHRDrcLFgo/CVeqnArqN87BQMUHTxOg841JOaKoRf07JcXJV3AchMTXiF8+Itlrts7yhviSoE
LT36Fd/wIXomj/okGvUTQwip/6Gxly701L3nVeiXEqxINKJAH2seDr8GVf0h75v0b9NR/DePX0Xw
iw96oj17TuxS9GHeyzRhQqyQCw1LuQjQUIL+CTS3dsLlWTHwHrbEot2DYaI3QbY9zclbC2TEfQ3G
D2Zw8S/FeyylgeKhZgl5e86N0je9eXIDVkhy8h4vLzgA4MMlU1QTCOdfi3CcM7AAy0cIiKI+W/m1
K/QWgEKH9cCTPkfZBzmlvjxX9b+Yuix4jahPJwLhUtYYGqi9EbRyQrL752l9FncYTTMgPJS1IUZ5
9hXJgYPAT022Ez+29+3BzGhELKgxTcIiolEn3RTJnb86MGe3O/m3IFKwyY5M2vjL6h8YRzGRq5wc
PtPqhLzMUbXwasZEUIwwxD3VSHfrDDQd2FrlVvjsJNwgCrbYna1Qv+V8vZomxGZjIgR1qSyAeF9L
qex54CBSlCphmFwzgnxtyICtwlBQuUJUxNyP9GpGYiAALdPtZhipRhV0Cb1FYGNCPXru01tOLwNh
PvRzEniT8d/nzJJp5P96V8wEmGWj3D/h/VtnbC9YNxbXwosXJzb8tl6cGs3HEXMVcSh4n5ZezSgG
4C94NlZStQ3IXLuH32f7rVJMw3RTPBNWc9ulPWWmLWzGqwm7lLksxfDKWW3rpwZzIGwC7jy5K1Tv
jpbFjFVtLCFd2vSHOlQb++3E2ITDqkqPFOnYxZXvrEus1WTxBHcstPKql7bVV2BfbsyPzKBo8Frg
5GW6G0ydprUyde+fjwjoMatP9UymgB1zdBklXpiEt/H/zRiRUEuQqYqfdAIDdQHH+euAeZD4TFeG
rn7n5tfuwoZJ+oPXETQj6Und98UeWm+OSlYCoL1HCdiEI2nK5oWtL6VNiQesKUMSl2yvxfRAtsgU
ns2e4bEqtkF8G2benlcNYNZ4SSt241NxyYZ0D5q/AW67A8jG/Ryn7C7pkQnsIdCja9hKq6EEZFDj
u9jr1bB6RCw+7krtaMom7LjXYJGG7R6b6qRPwwi3Is4HMDw+FxHhqQeMTvaJm9ebLwUbf9mPYCFP
aZIb7JOzIxfhLPUR6/kLGpWsUrh62tM05TpQ9/VtkQCAW8drdmACji+/+PVwgWUt4YBukPtkFvWh
lfne+rSv6pAUziOyPDFR+h+WDQOs8wRPldWLNwPbWrp+U1+hpscZ1elhT0UOcpy3pThtjf0aPinK
hdc4q9Dvw8U8Su/dx0WK+sZx57W2lEEWvBDkP4c1U9ZCzXHBF5FW4r0JyY5BgwUXw3RyR7oHBzQi
7kZit2r+yTeBjvsKFxDcIUm1dLc4gMo86d1NKkWWERblVOzZAqHQRXZh0byrsPjSdD7uOHmqnOBW
2ho7zEN+1rjh7FZx/oWjuqTlBJhveI55S+X1KQCxqq+6wS/c5AvU3UnKCLvkSiVapJP+SccLbSjC
W2PmuPjyQ8dVW23t9TNnF46REHtqLjIHRiIqZ4D7vf7rL43qsP+TGQi7VRc5vOJ11ZSeWL/9Tl0f
ObCRdw6jpN2kSwlN1saGgcmIvcMGasgt556ttWs0L4zMMcyjppTCGmkFZvJGMRmB17sXOi3FSrn1
dmQvveVueE9Bw3YSGAWNFbkNpuZWiW3Ahi0hVFjXUOfmwgjbGN365hKPT98Ai4RBdUxa8e4lVxPB
RcJn1yjZ1PL0UTGbqahUZai/u4LAYWmRXm5gq2UtrSl1VMoyQIjzDjdJbU5ymbCQSAWEpjorMRQP
DYaPE0/w8h9GQ82ib+++BjYDnKxp0aARUkkvpg3O8TaAfdwbdfAo3LiqeVYJmR0GVKDQUUvto9TZ
yZ+eAOG85b9f7ZYOCvBvqkO6/2lkEMEjIe9b9r66WVwgZBGKI8VY5dvZ2n2neuz7bLhzr6J9+/WR
8DpQ1Aox8AQv/faBRtGY7rubxh5eYkGIuFiBba6VBmjMF3rQ0lQIfuJof/UOJSrxklhJT0nKHGzL
VhrKrfvD7eavyFQfEXgHU/dODSdqRmH9FIhXr85w2GSMlWD55PIYe0F0+ixc40Hn8gmGcRk73/zJ
//+f4H3h8L5I9KFCGWav3bplmafZL5eE+VAtqxHnr7+IJ9ZaZmffQtyVha0El/leIdx+HFZ4oWYE
bhOi0aU87yKu9UeWtuKZQ7c7nZIfb/hQm3xafVNH4bWb1YkqpACROy/7FCGY4NwVhDV2WHWNdON9
5mI9vLNbDy14RH149bOxfve0ryOQ37gwRIrajv5cO169a5ka3IdU5i0iFtqgkLnwXMkuKfvGRXJK
Fb3m1bbsuWNZjogrCI93CIvtff8WYrhTtRBtNP9GcENrT7SYJMoUy63IgXtUQyTKhhQuKqrjNMeT
RV3evUVJlFDav4zJJUfnSEoRKFMAcl7yM7wy0c7A9sPQJeGQcvlvyEU8UDQx4GmxLBkVlSXDYcYQ
0shK0ytE0vz67IO71WNlfwkd+wQaA1JSrZCVCRHg9Xrdq8uUAJHjbJGpfELlg025+yV53V18o21j
aGfXRzBxHEUeUNJ5qTMgYOsaAb8qz7Ttwy+y5hDMbUcAlPcEfVH7NwNXiT1q9+z17gOT5XN/bKsV
8aN5jETESv2f2hylrK1hjfdo/e/7k8emCGdI4W8dwEgRMzt4D6uFcSJtl62ylZMLR6lNUUFEyRbY
gySKGnhLt1Ccy6R1KV+5D6qfcIlVBd8Ep3RSha8xxid2x4R/c47ZsZ6qYzD3m9cg3Zcmm2mfR9kH
VnzqsSp/ZvHYDtOynuQiawbuNi0QmTxb7XWJPxuaCrueskqD5ya5Az+W9a8yhSWNrvtxHMkuGjOX
u27Z0RUnOZdMt/FEzn3JGAhbqbJXzEmstd9r7Auv4yXZ7bDkSVfd+rjbnWwlVzbt4xzBzFGgWNX4
d84tVHw75AcFrHv1eBzioR9Difb5/oR9C7c0q0IG6fLyyPSdnZukLfiFCMjgqVhEUL1T6PkilKYE
G89oyWMyBqw3T28snOEyu1MyduZfDXopDoU8y2Ogp6sIvmRPZvcJTp3LlpYfzX1gOGmusnkSy7W7
aeK+TD0b0a01TbSRXIfV+2K/MK2MJeokwRLG9s7tt1/tIseFNfoMcEUgd4MyW9OV7cCCGaORlJ32
VfrvT6SdqKHKSph7JEy2jf7BPiO8OrARtDnXnRM0AcEoU6qj37oR1PcgNVy1m0WYpNMNShg4MaP6
LcZ6ECprxMQEnDKv81fvZqvq1EMrS9do6qNezCgpCqDL//HW/Njf1T+RFIXlko2z4C80sOxlZ2sK
DZoC7YlMXB+22pWFMBwA6sIM1zX1RjbokH7kOkF7Yco+5ioG3eKGHpZ35ByOEJS3yXsO8NAPZQ42
OrwTZFIvDCcot5KboWSH6vISFGjP/lClCXU+sjefOnZaKTU1nYyMlYna7wfiNnaF2DwzWTF8BfuB
WxBP88vF0zD6NzASoP5vWaEobOiVJfiIayG8Jy6jXLzgcBawiJCMjQFberfJvva8i5i7uT5NC8j+
9ANocsXt0HrSXi9b5fJ5a3Vwcsl7by9d9Nv8JVowQcQC+vy9CIdPWqAGiRBG1OALAsfFkxOWCRUD
wTpC90fl+MG/acQZmfIOrMd0OoGGXDgaEpgBRr7vGAIplaccxI8tgkfOrBHRDVhAeC+Kjpm5+hss
1xSLxpFhyRXYcw+N82z8pHNFOO2aKMWCwQIXg4f50gxi/Ttv757I3VyePgyNVFxcjy01OcC3ylm+
/RJWtMkYZzCyT8DtECLo7RXypZAwdDpzHm1hDtVBqCBKgLWcQ5YtH9+C2YA6iueFHu+kQ28vea/u
NVcCplgAG86Hz6XvuRgKp9JUafV2nyUGeCCIsF7vttxYkfW5gX8BAE5OHXrju+PpoYoKHS9XDrvN
TAFs4YnZUpSY5y9GQyqAkDhfdmt9+Qc0Ht5xiXn5GYPnkkvHlOPoQCXiqfprNRzvanQTOPT8OCxv
GSIIGvgNCg7aTEZwtnOTnwfmOc97hUHqyRDYxk/P5fgBPFi0djgIoAa/4SUnW+CRumQvBYxzu53Z
JEdOttzssSTxrkOB2t2nFCCXR6q7ydyhIYPq7YpT1ZaOrhnoGlcMbUXMgMFzd4QSZ7PyksjxJevj
0uW1K3l8e+nFyJ4jOu9YVMknSBFAxmBHPS/4AjZAhFFyKhjNh6hCSIpvEDCtMtT56pmMPWykoGrI
r1Y/XT7TkGRLObyTCi5+Bj4lCaHckz8qh8KmfZ44huxgAH3gqkDkoQtPbFWqCroi276jcJauie43
h+Qdi8UplZ16UcbAEigyFnwoyeDfB7TZzjk8LAHvm12w7R5bsqhQqNXTqVJ2NwhsszZ86F577+6N
PV24vBpPtdpbla/cp5U5IwT41AHQ8MApS9MGha+Ya5X5Lb2VhwnVNKgyfKbsitpkQfc2pQLLMtyp
tIEs+AQEtzwEzp1Ax/53QmPDtFkzmaEodTByOMQah24Yc84SGPfkocFMCj9gOq3qOyoob0NMy9Gl
qwcZOxbVzoAoTrK/KJKpH807xNAIbfj00IwjZVYytQgwDul1unZN0MoKbhjBIXT6gMr9XUXm0T5Z
cdbY01gRPj19eLfXZQ+4jgO5OF3u4OV5XUxdF/6J/3AaxfQPtiQ4VdbHtScNQyRwCyjnEARHFLOa
uJC/Q6PrKIh8wmST6pcVadEpnFLiFv4o11wCkNtD/1G1lOgTFPTExiGK5aUpBusU/ilNXTuShKJR
gLEZPfWD0aF/GObLPqGGp92E7c+dMUySSdYgjyQegjv5CHrTVB2KPR3JT8Sb+GQKRLKkQZhvm+Yc
uKYYqn2E8e6yxgRlbQw4Bfae0T/DT3d1WrpRg6J8wfCUEU7lr8QFUicrxGiz/T226Xay8Lw56T95
2cgqWJsOS0w2r4Pfo2t0bG4xJZXQ6EAHju7dLF1trLAaFuwxqena0wNI0VX+pspT+DDg5dJyjC6b
14cIU19w9fOv54InVJ7VZUOjYQ0I7vbb2jY+t85sI08PYuLotQsmlnkAHXHMwQUMfEZvHvPDANem
tCl9dT0hO//oQIm5NJRVFAAN3WMEepi9I4eGDlqneD1Rv0jvczg+T+QAwIlL0xvInS6pNbVg4NSK
JmKAwv7kQt6Nmdaq08/fIdLiZMIqP7zgldokaJHkDMfr2mSDN3cJJO9U+LuYIexQcqPpcvVWug7O
P0c/QXgAf39R4H5Oyvq0mcsIC2uC9LOYH711E2f8zoHl2i7NWITnJuJ/VpwX+q8Be8Sob6iKMFnY
R/XdL6Fg4iFJJMxiE9LogPh1Yl5cMIg55cRafXVIz63tYGY2x4W3zQr7v7N4X089Ku0+xuo9+J0E
qY06HIez5BCN4+FMzeEpLFnrgOI5xWrqQipMHoVGcDLemiz9j6LH3nO6aa/elfiM7/Zhh/p0Q0pq
1sMRj5iN72qoSDMizjodmVX28b9b3VS4YAedVEfHfFFBiP9P1Jze7baSCW4YLJAV+X9OVxEnlwTw
qPWvHFxYimhYyTR2s2QEvpXDZFfwn8VH4saQ3vwCah9o07hULSDOC3DwSEk0n3veAAGKYnfHiKr+
2J17QG4kF+lT4IYj6KvS1SOCamdq7rqcO1jW/fLKgjEp2dKB8NJkmrlKTSWtIFC6hbZ7euv2v2i7
c4/lEGJ3t8QS95ITnOnjo0oAy7tYxHbGx0KDetzAtZS+Ipi2z4u+AZnvrqz/+TKQ02rswJWfP1Jb
UsRIAXmuqp1m4vLGurwWWeQmIxSxUvG8gUHwBPH5O/0MNNX94B+Tkm2yBCjcCRdlzd+r1d2//1Hu
emf8MigUYH/hZ5VAS4gt3wWR2oMo63iAcZJWL7k4e9UdevrqxJgClFHMsg+o62lFqenI//yCNEIn
hBF2+4ZA/Q3NYaajO/wz+2LUWv12/B2NmN/pb0lZbMmo5eQS13kynbSmtTJn5mfgVCcF9pdRiw8/
NyfuXZ/NCaEeNB3yE3CrVbxJHTUS71XmPJPfaeuumcBMe9F6q3RLL5Orn2kJJOggX5RBlECdEUFG
MZ4rtxP0K62CNFa02gbX//dTHyqBn/sJsqdAXd0BXaxFeK0d1uQM3GSmBQy0xwlbGh5HvMKL0YC+
9iNsp0Yn6Ko0UGRKgf71dfY8MmG0dEK8jtAqveV8DzFBmyCPJorAonGqS7egyCp115JpvjA324QL
FisN13iKUwV5C5Qf1I+wc16jUgVd9EG6H1HpukL+hkEkC/64Rf+d4dypkzYgl09mJYYWEdaVxsKY
vO3ZWBfMz0p2MTI/Biyc+MwykSGlMaOMkC8IIaQpDXlfpl++hlFJuuYMLrvs/DgLSzRbVXCFQcxj
d5Zl7Pu1/7qdcZ+m9Z2GitP6IPyYlPWT9HqdvGtHyfmJ+K9lFLk1SG+VrMM0S591QP39D7kVW0tV
VbFp4vYWtii34YMF/qL6NxbDX4yFb5x5ggpdR5IdkJ8eEYp7j7TRPuo6zMvdRYBG6ro3VJS2iZQK
LqUIEQoDU8I6btkGtgjmd95lKglG4r9jLOZ00kDl9JmrmggeCXmYWrLSAb6pKvCh56k4rU5OPnM0
SiZkENPUnORav1jFjLxhYMCGTjAjTMriMAmd5sqlfmdDQazehCg8s5NYl4JFk3ztEFhfXYRnXzzZ
15AL1RwzGwucObAWr7YbRXxCgXENamuzNSuMt3jGeRkasPJF5xpbBLhu0UkPhvqR83PvQq4Olu+L
EYogyqWncSrZvfXNp8YvwYqhJ2OAX6l/E6hChKNBXMFi4y6keztGaYa9wjpBqUM1bVl02Z5FDMBl
bCDj++rlhLE/I//aTsxwi11rQdjoxC+Hzyl3RgekebmkXcbjg6iINAsyGqtFcU9u+jnQZgbP3Jvt
m8rozxXEWBs/Ctv2EpAHCcLV5XXrAYW/YZUSLrEkZ+llfzPo0Zpalk97ARrnsnbvEofHAVI57pUI
iKwFtDo8cYpTFDpG4R8xm23L2nshXAornENzPITAq15RCFY1Ua2fgutay8pq6+EYgvPdfZE93zgU
BbSAXPqqjaBXFhb37OBH+5D1o4DF+rLUYFgrAaOEEevUuy7y0NOk3yateDGXussiW0TPwLIvXZcK
ir7L/CxqemWYiJ3ywRoyDTRS6GqvAjHocj3c4ko4dyEQoRWlD/OgWOyfXM/+c3QyP6JKJ0UGnJQT
Jp1PUpZPT76F2kc8wHoPuCfRzsQGJndU2uSnoj8+TuUHZlTUqzMDe2tgcoqrmJ+C6c1Dd9rnAUc4
IIFTKAUyy/vjD7ZSydO/ZaLMyeSY2bEC4D5IBjEkvcpSd5N5c+ka0d4JEaiPiBRBWjHAKMap9Dn2
hm5Tik24x/ebXux/y+WJQjeoMqHtjAb9mynJYXfBrtbUL5WIXaRaBupypUXM2/QX7n2YHoeTI+ym
ZLzgKe84l1Kx/G/1qqoRMlxlixyK/a7YN/02PgBP4ccClWSj3W0qbPi5ZEbFET2bS0M0t7WaCfnu
8R0j69GsrscHl0LrE+Ao2NanutPrMLHxml+NV5ebdKx0+2bPDTmrl8PvAJrtyzhVgzufUfgQ9WJL
wi11KnuiOElIe1ia+Vdq+WFUOqjzJMKN+PtikKiRm/BJVEPdbmCA1gXZ1qHJsKOg/KahXN+hapx6
S6720WSxrGxKyS9BUu6fa81Y49rCj0wH0Tge1j8MrNInb90uv3Y2BHyWAgwxMAembrdvKrxX/6/6
4Nux4x6OdK5ja/87JoS8+yVHF8bXCJPhPfjSnYlB7RFjfEx72MkxYfhflu6yURExsUnJJkum7IZm
bTU4WXdv0BdGuE+ocokYcX/WtPrHXaos1KlAOVOYYd8c+ztcG/ZXlNJJ7VO/SpxieXvrdtLEwuYm
6suf7IMav2HDiINCKkmUNHnUVeN6xqQ1CKqDXp6UMecVKDXLiFtW12meuY9OZt1kZ1vaarmKACQ6
VNnEz4FzElKuvuEtuDWifaRze1vvQFDSKhUK/eH1yuWvEOJWqOghq2qkFV8A9TLu/j11I+Rp3iQZ
++y21GZ+qZSbC9cYlqX+pRqhWQr93MLBiI0LBMLSOFEgPaFQYWR5xggi4aqWmB40KJeQ8ccYR28K
9E9rlYdM1ghxBCD7DMvFKiCVBBCAU+LySKWNwiE/8Tb+gIcGchmqz9u11T8XPzQo/X1cnw7QF48K
QP25FgFaGvdim5R7Qkdz4hlpOMVryyoAe1V9k+x1YCzKmQ/KUEhKuSNnncZ+7x0rI1t9MTCUE0S3
XfGW4EcsTASAf3kTPER1ilgjivlOVdsaSdHMtKs/UI7oVFKmzXx4TH54tHmMr3FYUOUd7mC7aF1X
OeOmub5VpI39pdXUYTa/CS9MaQqICCFVH/zdSPBJQzhKL3+AJ4s5QbZj8EcjKw4Q9vFDyMxleqFs
iy1rP7EgWJJPtMolmBKbjP4PIn20CdBY1aiy9lkIUB6Us1TkPJLYAc5oSiwGA3kXCHP/GUlgaJax
97Sw7jqfjHPQCBhkqqlCm25VfSUhEd/LVtlK6UAglsFWuIFyUj08fkD7RO1MMJARenvo4DN20XYQ
e+J7Uh9n75YT+vSqybytWIlfvptjEn9c+UrA4XZ+IcL+9m3ox1YKzydSnp45LMfn/NlWaZU8BeUN
Xz+n9nULbeXKhcBSPspbSwPqqBGIYhgSKSy4uTxa7ElmC/1pyq4cVe2uG9FJzpTXIdJ4TTRquiga
7QWgRMVdaB6OTOTENneR2pz2pTlSgjFZPgisl7gZlLiB5VbPJ+iyR8GD6nfHjkZaNd+jNTpydWGz
x0AkGJrHh/m9E6n2ZhhdHQ8uynSwY0Oub1sWr5K6NNY11OpRAY96rd91dskb2Mo7zlKCyy+QTIyO
eLxMPaprcBmhRy2zg4g9WleGR8EygspP2PnW7DRiO50JYrZNxXiN+6NCi35FerLILQGwZz/1DfB2
E3Hm7sma18GWVNB8iOS09+ZQ+vpC6+U7TtFg8mPmOoQI6gjRExLiX7+vtRKTgD6Vi/qfSj9jMNoJ
QDQHT9ugv6hlNbVc02vWbt1W8z/eZ3CcEkf61GPQCdGZQj1ZFg1wIqADy34ASi8/ygoHkeC8KCd2
raXNkhDkaxnBCxeWj0OVto5SpcXf+fehuiwOuACXQ/oCkimo418T7i17O2n4osbHZzh9pgWg6oir
4q69c4DzKGJ1Xba7695lyMNkv00v20LWpZvZjRwa1q3U393FflmkwCgqaePqxoAofzZxNqOO4vhz
lyQmK+Kfn/r+R2MeZKVahWMRTVcxkwoEg+/dRnL4R1OWymuq0eAfPpUcwGaSQ2rj+mTjus1lsh8T
qYnUnGDUz4qt2LNuhA/Oy0UmBTcPl0mZF7K0ejkIgcA/vcotM9vHAZV9QkmbJiY/rzzqHgA6ujqX
0q4VPCwL3wvP3u7fZMXXvv4O841Dwy4rMHsJdWtqtfMxEI7vIWJAEAPdZsxSN5iKxtGhuht4gyLD
6habJQEE0qb3U3ZgawzX0h2oWnPQeR6JkSo8YpvIr2juTJYvK+gfhzLrpCFdbl8bdGeVO1vlvZdm
QXScCgDpCLYwHrypWqUSKzthTAWFLyXbExtfugac2vdsocX1vtGKZVVi7xUazsTE062wvmhcVOG7
bmrLEMxySe1smJ9mgpPTYsx72EYaMSYf+6U57vuWqpsPu73NSU6n1IyYpaW0aNLopj+VXxNSnTUP
RqrIQ7450nzDele9n7ZlSnYau3NwMEH+7PTxOpmf5SGsiHSdb+t/WxOGubucIb+K6vwTbOSo1uj0
PtICdMoScfa/WkJdXjP8DWXoDN4VZrJZD3c3+e7BU2Hv8OOzzgg2WT4PgxGemVomBO3H/1HVDyKL
8ZMpIDODHW0H8Wbk5o9T4bn0oCu2IrlBnccnIhDf+oxnoQT5FchysDerKw2vuNw5xUpyT+Uf7cjh
CfI37Qz+4WmXbDF+2YTuvdyNtK/ln7xNZZ0n2L7GyO5pJi8EPyE/6kroMvLNnqFM/qxbhoPjRtiV
DyBU6yAiU2JqODPJEpqHCkGQYoLFl4RzWZ69fHf99sGZavPR3X9RCIPgq2MG4dEXfWjmozq3Di5B
FdeojYNuFmc7lKyFtoWfL/xQDNSpGpd5skRpwBRo9iozbJSSK2LQJp9wvMuCBs7oa9uco9KUWBIs
iCb3e07swLough7HtaOmOKFjVomvs1vACLFvKvamSsWOiunKgw/oSSX1Vv7fL/V9gaLqZoraG0sK
YFwBqKp8l+KFYjatgn+162DHmapaFw29HDaNya//r/831wtgE/DTyUsJ5WjxXl2ZEhMCiqAg5Tt4
I7pRhSxxhojKIsD2P+wZcmIlSggQjEg38t58xmyOpFUHUqrgROeZTXQS77OpOAHikquh/GM1o91O
8jpgiUc7BNh9bnS0IlC2yloMRaFQytA/lQhJgOn1f9A74FA18sMdswqOucoOL1Yo8NskuF3NycUi
+6aqjsVKe6uXJCErm6KizDsJplN7XpnSI7eYg7t5BQTwc5u/Dyb/Km1eAXngfmWVhik/cZH0FmEb
4iQYc8bcjTc/SERdnbMtmUDGxlMenozfBnyo1Jrh8LULtjBHhjTqn21XhgwpyMBse+MLglvgDCYK
Br2w54HhZ+ce7rxpWNZz5/Y9x5Pvzh17JP+vZeUJ+gbAr1GNIXGRRrzWd2muzXVZq8671mVZN6Q4
QqcWueydEPtbMKu8yttHBnEgNt3j34fpr6S40ZBhE1NQMmo7nYXPPqVoOHDPFvQpI1s1P0gG1gYJ
gAbNO9ea0i+GrUoYBKbtbFkpIx+RTc/w1qzwemTw2lGTk7ZLk5IxLFbtksHFqXqIzdGwX+9nNX+P
D/1RuCmb+itQhlHYi/50xNrPAFDoWgXK0BZRHb2np+M7B40rHpB4VgvszhFSjdGkfJrQFbfY6jZc
VI+5Au+MYqQrNs/YqVtGdrI8i3x1CYRP7aeKJupq3y7WoR7Kg8h5TD6MTv5Pr/QxTj6X8a6hMo7E
VyBYghaOHJowY87xxq2taDPCob0V4Sx3rNdsmDYoxv1BAcooEUhmFhtiHnSmxYD9vYzIEaX9HQc0
MJc0ALRZPreTPmbDB+snROdkwEeBOY/Ov5nPjT1AkeGEBbval3/tL8YK7S4RI+99glimzr27P3gI
vMjVJQt7pxLrHKzeqvvRkpaYnyzotJJ9RNigT4bx8kPH38iZGDkyQUD+5wtdDv77j8E80akUQQ/t
V4p7LnxLcYkPw2WM62/heGzDPwvZy4Yoy8/9VVlc32z/Ev9TX083k87Ti8/1PBFVVbppvtE3ITKg
kNzptNswF99DICHO+CDmhuLUpCXXE4+SjZ07L/0AYTyGAYQ+a9JvklIZWHcAxKkjl8ewh3XNr/Q6
IdfWcBK+ONa8aHYrW+y9uqpvbyjQJgRUKEPf5rzWxMXSgdjifaqYliaWH45KA3JY5iZNspndaUeI
m2HYFi8yK2TTFIwKreDDi28SvgGLXP7eCVPMJjzO42wSWCS4vqqZGFlf7oo5R7IfWhWs0PLsrujF
wXm1jk+75LUi2oVFnerlnVelPxotGJlRRcESl/Y+20JvQb2EZhNP6wOuGVlSIwzL1021tBLfITJj
G9UX+lcuRwKYg7YRSAhTK53723nhYx/aaeJedAuAz6EYclGUlmLKSKaynau71wQS2mWAauJdmpG7
TkEv8ZM7aS5w1uKWDVQw0TqkJRyPE50ZeNwQwU29pfRPb59KZbdh2E9o8x9sdIcpHShPQ2Ql8a8k
SGdWyTUN0eOWQy1oHewC+8qDE1oiKHEC41rTFG7nUuKS+OTWmY77qFsGkieeQJvE8T05GuafV8dX
9g5uf6AaRmCHBchepEdrEFuBUyLuOKjjUY0m1O9lk/nlxWurVb/P6wsN+Rh1k3gpX0/ExrmgGO8X
s57cIXllRFDIJX/wiexEI7V4NESM1eFXaJjlJLwmRHD5Qfhxzqz2vZ+wfdGEOnQ2wAYM5elSoPsO
5Aas/KJ73n6Ny9Dy28yWU+BYkbPGoyRUO3DUd/AohxCYkzMTC4zQ/438j35BYfOx7WqOk61PPNYp
LKXgiPh++hpuVFfeewE4ftB5W7ljZQnkG57qM8YHJFYNetjUwjcuWskVQXI6oJ5zLAv5BZm9g74V
kI3Km7p/AfM3NDhpPuHJ9SGVxTa5PCLOKRZWCAqwAGy7ECselQA1von3MIYvleoVcQEZ+DYYHF9V
rbX3beUglwC7POz8acoRKTq2SsvNmdLFo0JysJLtsy3gxKDOyNs+Y+BS/e5dqchSPpK6vMwRYFOJ
aamF6iNsz+OMFMRUQIkGJ9lZw51sQtY59iQ9yyxRf8Qm5r83KeS99JmRLE0dVQAndyBCCu01qvkw
wVliDe9c/51dxMPJmrsZN9bWGdxsLPQXilAYJF28Qigq7551x//p0h7TnSJW6WJpiSvWT+ko2HOG
AsL8fb2MNphaGjA6iRaomuXuO9KBycLfU/Q4RO0nf5qXAep+7W76XqV067WLlxYiqT2qaQuCSVx+
CG/CRYVw1WfHb3KAyknj59dnklj1xaxsAuAhb10MJvB+Vlhn0rRSrPsAl1bRuVs83A6pjI5JVHvY
AWeDWPIGyWREG2muOQsGuV5jGhp95hQlJrKdJ2e4Ym66re0QafZTw4DgnXkXeQVmoZDUZiRa0fLS
cywNZ4BUfKTicnyrSe7JJ0/5JvGBHfYg//ADgpA7mTabVri5AZh14WqaCc1XXEmKh+JwNafxYzLl
YhFrLh7eg9+YtfuVN+mJXmUVx1JfRE58+2tfDxfWz6mtGFrQGSS/LWbBWvcZELJYudv4T9JcXL6J
/90RyiKMTZRNIWpYxJSM49nF6S9zUOlCV6yMC86qUm+KrlUAsT2jxmi4jCAADotRTidzIH7lSHVs
CRSlQ69a/aB2Mcl33bnr8RIruY+z7EAWCO20ZiExw67cqLf+Uw1iB0uuR0A2rpHvY6w+X0ODxVFJ
Ojcos71jc0T+lDCICFwNks2TqESO6cmA5GatZAikWtyp2OFTmVEEubgMMbBtGHxq7TjMF/g6/Ydl
nJo27ShtREdkKPftEHhnYSJcN9czUJ07weIU4s45MVZ3uZ3241eOACsl0Dw5sLjSHUGqN/vD0dmj
JxyF320r22sY2lX3YFu8u3sty3qejBoAhjNch/Kofplr5KkFrSGJGbWeDq0afCRFpNDi0gCbiM9n
MZvpRW9qYOpKX+zYUQYixjDt1kRnJnNTZ2+Opn4v7sqfzNB0H1NuFnJHIh3DL++v0aLt8DqQxxfF
esYYiI993kMcuOpADnpb0k9ZezFk90wr3lCJXU2ktO9kRvez+JdpHwqeJcOwjgjKGn9uN0aTYjxD
83VkgFiPavGap+/1dORPhLWt2pSsqaMTOZtgNV1IHJU+FUsyNxaOiQN8faXLUXJVdctceKG8eKjX
2bx0RV6WC22tZSVO4WSuZ8iTgjhbhCbMByf2dswNsNcTmiFMM5wHAfnklJEo8/WwPJomy08h2XVl
iB11hqcLSZGPxhjtlokWhqOPJ+fKVccsnAwnzyogcMPoAcICHyI0jPbeOyileonPcHB8rrS8dfyn
wdpmd6KjrbCNA7Z4281GYM8YTnR9zSUcFm/TAoNJa5bnaBDk29JA/9YuIwORsjYqw10uJgunnPwQ
511kjrPNCaswJ3asfxHmama6gCBJturVo7CUIN9qyl/MicjllatI0/8F7x+BokX6NpvSP4Q+pYVY
i2iMcbaXlR8/v8qlXrqWBJ8LQu6Q399zuurdoa112BjwKptZLfJulasIfV13cqZXJNHlwUuOjAq3
CyczhXK1ejzQs8b4S7MJ4LiFWmWRRI+UFjrOvzuSGLQN/q60z8FHa1VgbwnmR6geIsFxExLgFC17
3MX1UG4Hr7DoncJPCkM2orupsrL07iYKUAvhhlIt5IcIm8mlv36F+P+CDkoKaKGYymNTzQLIT/AM
PaM4opy6bJ475/sXmEN5oz7UgRXug6ZQxqT9+p4uUq9vewc/GDm4hL6ATg0pa1/7R7vGXZWDDVA3
uo866zlpThrecPpGkm+8qkp+fo9n+rCL+TmK1f6SpupQ7G3yosIsf9JojQ7hXlKXIVRXwe/JIGQ7
DA804511PkSaEhoRJoCKpOTTRYf9Jko0H68DVCE7wjUajwaejIsM4ErHK08cwr31PNKZE7PXkHb4
p4+nsjpEh6ODtyJDqilBAwP5jiwFDyB8Elkuc6f/CzqhlV/+PeVcpmGBf+PbdGriAUpzsnoXO18m
79egTwg8UmEvb1Bd9lUCO3OeJxqz1IS46GCQ2T6ichFp9jwwshxNNlVQeb72lPIa9hv7mUVryv4v
GBiDoiS2HDWFfPHPAMp3rhDkwNY6+HvUSBNxgDQDkcRtPiDGUr8H7pxVSaTaiqgx3gvPRyLJ8Rw/
9HZakYTZ6Up/lH/jsv+or3y6FmezOVlP1YNd3QXcrmO7ryR4gzuKQ6A6OF1wt+jwb8uC8Hwxttth
b9oHhMNuKDcESbN7ylk6d+K2D8QCO83fc6NqiCy/e2vgBLiR4EEAH87JBvVCUdYRmmSJNSSo4juC
/FTrPvXs24E3k2P5qgUP+QDCr6NRJDQDrfyWQfMnAhjoUD4OBpiomMmcZeOje9qJwc7h71cYF86O
THNsqp9aAO/zPpnc7OptHeJ0rrf3zAxhbhkESvnKQRInOVlXBZJcB/OsUW80OJ8RvA4VnMobAJmB
Hue2/I0ZNKGTwuWUk6jrahxU59u7xKcNmbQQ0w8x4cyBf3OhVqrJEhx7DG1lpy7ntrrlXbR+iTys
GXg6fZO9jlicz11LsMJHc+VZ7OsudS9hxpHkkp55ykAqz1PsCrVfWr+ZZX8hsVXFth+Bue0can5w
vZPKs+ejIhFh/6KUdk61NRs26PuEBH23ffWR3ejpVmFp9g5yZDWQ2+fgcqAR6nCapMGtelWa3OdH
uYYKDy40oDh213J90NtTd6dq4oVP77P6vnRMVqM8esgJEDex5bQB66cA+/gjpDHJ+EhhSeRIGpaV
ncQ0MkeovCFtDTfqvNfIw/f64xAgkx/1lZ9HgJVz7qHcssE+hoG2xUqN3VUArzQ/OOlpcf/6H0sF
wCEjUfZpRGdFQIit38PrEr8+e8xymJb2VBttL4xuh8QNTL/G1JgY3Zguft3HTMn8dZKxRbyHM6Sz
JcJcmdte5101sJFfPek/CAaZ765uCTIk+/HFvlZAY4dojm3C5ygnaDFb4vrYDVQtBgrQPZlpQOxf
FGkB1yjXfoRAjqKyD0IF7BnghdrRC9onTZSTmA1DQa0v+Z6hRFYkBUZRTwgID6riYh6e1h66Mt5D
P9arLqKl6peQ5Z81YLk6Li3wDj7aV+IWS0mMXnea1K1AYv8S+6wWM5P8sk62UaTKnJaQTxrBLEMe
Qyo1tv+xu8q5PUN00zGgAuHYnCWp8YDGqL0MrVhu2Ynf9gRO5v4z/jb12Y72/xa3v/AjS8JfXFnm
o3v4OfOc1XJ2+a5YEhWRz8X1tVCDrMzf7BMZ5U5CDiFpr6okB3T+uBv4lVHNbecEgO7cbYCu/2mZ
W11H3iVnN9DHVfQRh9tsMQT+C5OHJecM5wZvodJszdruR2Ojeop704sv4TzARPDJvsJFDvtSTsfU
pizPgzZs/g9yH8AzB2PAHlYo8mipEtPHhkV+5LBFf6N4zIFCTWT3fVozu85Yg6SzfhCJ/gLwWR5N
jymBqYi3LeW1UJ9d+kr1Y39WpW9/0cgkseWc2NKMtaZ6H6v2KbpM5els5IRBkk1J7Bz832buBKMI
RpPKGBXV9BI7sLx1S7Y4I/ceiwBmRuFW5NCler/4p7kq6dkpZlP4gnbJrHL46h1z5+sdpX9gwO68
ZWB5/sN5WwmWZlJ74UQoWeuLMLphJVp5TREQjoc3dkpRJn/lVsRjFWrcJFOD9CSKdxk+iVeywD17
2Kxk8+7vy3G7W0xMlqUnDHfAM27c2C5F0AVoqMk3CT9PjtZkDwPEo6efxXPIItEbrvd7+2Y7MQMj
wZoKAGQFokBrlCai/wdqSwC5N+8CF/1jNZgR3kwXauGC6bKls/TztlVF/Qqhk5/eKU9i4ZlUr0B5
tNZmzbaVkYJpaduR5L4kgkHLjTKs/6eHb9uCE90C660VaR0K8kUEOA2uEWDvkYKu8xEdgiRBESba
c0hM006owPcZlbgekJx1eqhzE2JZAXXxlt4SaWpOq12hhgQVHfxWlPacMMAk90Nbri8ylUnHs7Lm
DcOZLWF5J45aiw21YJeScPSZsMdZ8qxa8eFcMKguKNR5m8NOhSCk3FuuWuhKOyDjtyqazF/TH3uU
HB8ZL0gOXQklHTEXmAjIhdZUdamRy43ZfSclXIZM/4ZwGx89tH3ATh1n4vBK22R9tF9tqh90K3Kc
2VjOG5lqchXjqeVd8k6LpLmklda1qO7YgImzI1W+pBl9Ai+NXNoz8INSe+lHT9hOlOVxLkLUETrr
/PHmuJ5nnn7GX3AmuiL61uCbaVkXGQYI/RxFk11DTu84NE1A35HcL7SzWHquDWlO9diXgLFJyBH3
vP+qrMCk/9lbgYXo/Bu3A/G/lLr1O6lGIfRELOAYl2BD87qvrNUceTPu3pxNqyeGlK54ux0gKDsu
M7vn4rmjkkwI5hwL1gUOwlKdKSQZSo5UV1d/56/o347ed1pHYvtX6YW/LGdYKA2GXspAAcmpB8UG
KCOBRX753jGXfiXEftYvXuIYr36mA6NhEtOV9pa4sVgQ5FWIjzDQ7LayrUB7dFO96Ax1taB1EGeA
DCxmKKznW52ghIbe3fbogc5peP+deFT/6h15Q5fB7RQM8n8l7bm26ZqXETGi35fqOWF+0CDNY3AK
i2WknwwgI6HY9bnEZKRVYrSifpBrIznDhXulCQaJpL+h+Vo1wMF+AN3mM2iaedL7r4UzMNXd9sar
zlWhaV5A6a/kVLaI4V1pfZfZYXCg8C8m3Lqd4RuOGS8X8STDLB2sPkq0Rcn98aDp0BDpaPrxLMU0
fseRUizu9XnTt4V37gW6HA/BKYd1qEOqq8h6dn7uIySfgPy8B8hxhzYxYg1YY6z2xRsoOz06BGdF
Z2mSp7MAunzeKp+Ewc3PFLT197l8WtRFkNpDdgHCrgFntCQoQHZ3S8DdVo3Ppz3732NyqTl5jWkn
GX1TPY+aG7PLqVqZ6bMN1oIOGs8iWaPEFHnhTnZehIxJy51MzgSu2HGuiA+zBlxEl7OTIS+p2LT5
Lri9c58kYKHEMJaU04XaMtnmsDw6bO/uERH/Bmryf6lfh7BNzuFPElRelVwQHxsi6IlDxPk4NiEm
mOuVlAWwIA/81qyrUh6tryYRqYvYVgJycE4boOHOJ0ZiEYE0HJZnvSYOWPnsK+lhDjWVfLsq666s
XkDB+GwdmfgcmZF6/AgF6/+1qlxCrtED+/l17s/2ooUxmKnFnc2Brl+gRgbOY3zMeC50yRjeA4Zr
d/aZU1zOaVkysBEce0/XnRF3MROuGv4ALmqb/HGkHcJTYg9AMrCYhS92B5zrGKwCuzls7GRtIkIv
LlmbyviDNTpbs00SzQchVNH5lcih+rYZ//9pEdsmOWb0pRncxmjgYHP/VddZ3a26qA6EMqOQvRlA
AQVuRXRlPCi0D6qKyPkSOktTKlqY18F716q3eRiFkA7rRK7qcNHes/J8pbpgFq+DhCj+A9BSQf+a
rS3q5rbVcowmfQLgW0ZwCS2wTSm14FSx4dFqcTjwRZEc/LLV87FCTC5rT4FCs0buI0vTw9YLL2bs
/0OWUY2ucmt7mINNj7T1OY+osVe5ChgKTdJz6K4vQUdf039SJaIXTBd05jOgMOeI0gDqrY+Zc1lX
nO1PgN5x2k96SFGA7bRznbqlRmg34FWYbS5ZUmj43hVawCVxtiVgSI49+k6wp5qbGuZPH4yaLPiq
hKshKBLKBKRmYqEgbkXLxa5TJ3BeLsP3B/1z6lbHqyoEXen0TqWE22h1ETxXdzMgco0BrNawvHwM
28fTDj74RsiQ48ZaEM4CdTxBI1mf+eqOBkIDFx2iq29Tl5Z7zV04lm8c4OCMiIFC/vT2Dx+T+9Cv
GCE456PNrj9R7OFbsimbAyP/rZL+zu+PmSKnlNFFs4Wz8SZ3KzbHXTVBvCfYBt5Saks9ibtb+3U6
v08N7bS6mwaWe6wzHagFrnFNoYZl2z4rZcRwE+m69p2OYxiJVcTPooSr6RNKqGcLc4vXU9gtPE+i
i1DFgzqGIJlPoC8Bxag4i1fSp6XeKbarxs6ZmjFoDyQXtoyhfmJo0HnJRm6xKfFPtIL31DmVFKXZ
HE4eCn51aJKH7YVRhM8KWizZWw1a4y3oQgw/+J2d92/wG+MY0A/OL2oC0zTnGjxe9VcUnD/0O26h
yNAGxlprPO+sHlMO/E6+MgsZR2EXBP6XONV7PdnM6mnunNIMiNGwF0o65mvVwwsOR2HE+uJgSbWx
4xuoSfU/9IBD61nuuAExUCfhFG5pH2lRCEz86a8EJtLCIH3DyByJbUqPQhjR8uYuZq65Mo1IpwVD
gZYxHWP3VWk7EaU37KAeh3NNBtWND9d98c7fD81riQvJUWm8vqkl/5fVAKFY7OLQHGSzGTmGu9x+
4tIR4eNdnZLmLYi92WSbXsEgvz9hoEjtiwlXr0W8UWFtM8Yo81AQef3Yy5J/kVLib2nmaKAtt7zM
Z7lPpO4i2eKYB1E57VVuOFmHNDVEDvciHgeFQYUiK/i6pIq7mAK3kFDVKzuvUJzyCkeUzK/GHxGO
Ycg/9AAog3PWBWieEtkefgZ+xN7ydGhS3qVyMEOno+lo7YInxSzNa1T8yV5C8cMyObYCovzKdbey
dKLd83341vKjSRWmN+CdyaKaMK+JnblYzQk36IaCXnuYGfmHPNoRs9fkQowo4kZtcw4PaONxek7p
OzDcOM3/rmUMWlfx9FMf74po2xmtE5q9XqpAfafHWyO3s+nrulrkNipieg1Cr5f3K7cQMPw0yOBd
4NDD3w/V3G6wJbIbKbX+06/Tjo9l2QDAQ7o7nyJL0u/53+dDH2We3sFMybg/OxBLgpQzLmiVh3PZ
81h3oQcG1XzU17gA/TisqhiPWeQCJE0utAa4B3ztBlMxmi4dFm0uyc4pQ6esC07YdlJb/u0GVmMs
deSZAa6jYW8bzmBLOmizCSCtqw427rrihbrIn9X+p/BBKQNlG5kyIwRLESMWsJifnOxOqfwjdsfl
R/lptzgJDiW3TKtqTMFwagsrngNvm4+dnPtxkHSqaphhIvz3lLzeAVLfNZ/QFBEyvUrRKJUO+wg7
Qz7GHazOlocTEHEga0CIeyR1+ZI6J0XaPtUWYfbOiSdkfUruXqzthN/GEKrUZPEA28VL6s0/zR3e
fRYQmbZA3GFHxIRL7GDvIMOlmnhGcNRci4lTZTO0ZxtA4F78U9MK5X5Wlr5rFIAbg37U672zjlL5
KJzvP+SZtxDRLcQhBDOM7eZ9zM6IaDlAqLI+gwxUOZYxdgEnFC/9cRO85p92si85Tlyt1n0J64+3
h4sWBi4+Ue61x27TgIDiEYx1Q/vULeo1lk3D8reYQFn+iLAtW31fg9HG/Tpr7p8XVZK1b8D877ZA
qWrXQxq3+sOqDbYZ5FuEhbdvlOrXjYXcCseIlK8T3AQ005TKxBp3EVuxGwnOqDYqX5E/nJ95MNT0
tbF7H6JsNA5I/TfwpybQcnNzf+LYiOmo1Hur0I+1GnUEwAqf7leN2B3C5R1eVhMDSjGK2ka8Oktw
hRIhffvi0S2dkcvVBtxQF9ZGnsXOlr6sRENiPu9V4NCBt7J4ZSQPDnInMO5RQAE+lGDISbX2x8+D
JrCfhqm9yIZD/JSKIpt6gHa7wfKamwMta1biirFgmGKIalzF575fiHRQ0ZcbbhP6z5ky0vTlgIDZ
gwpwbd4Zesmek7irPDogd+SuI0DKgzcRU/euVWumi21ibTo17IEDvTKYqKM54BI0cfbXlLlgE6rJ
hCI9wMU/sFYmk1VES17nMPLlIQUe9s+D+WCXUpe/fSAwTD8ZqTZk3AacdCghYw967ALxJ1Bv+o6r
TFSYkhzcb2bhJEwWH3MwAEuW3r1laUgFg23UGQ8OQwO6bZdawX8fD1I+U7QoVPByMQi9HunD8EXq
XNBFbJnCcSbnQy6T4QRrmpuDU0JYTTRsnJGq3QRJn6/Mnl3LrqkRwhyBrYg131zndp9DTJBEUF1z
cRr18OxQ4aCquDjUq830fOHes95GN7rK40xIEVfusp2ae1nwmArEDmO4eHLGPxBVgnSQtoB88Kh5
ejM0kox/wbzKalNPLqhuKyEMEyHDJXczgPOVl+jNS+GPNG4tPYod8E4BuVGOdscI7X+f/R34nxQn
FJVymviH5EOwgNRoK7tywk0w180EzOf56aZbJnpWzVwESUyCsGE1CmEpd4hbu/pMFQmkwnGieVK/
HFp18qHuqmNZ3Br691b+IQwP2B902zbEw6o5swu+V+mxCwPOb9dgHDs5gdW6ABdg4hvsL060lP+R
ffjy7hyBMUhlGxWccQwxw19X+G8/AmH+4Fzoa8KPgCH4Nq4yepNRGu2w3PicbP+p21pGa1jiyx9C
KuCmNWKWy5ObyOYtK5KnWAgO1vQZqtfFHm+A9k39q22jyxTq7qlS42N3yEOMgtpb8kMb2XDRhnAk
9ATu8i1qbG1er2NMq0JgrkZuXSM+eXWSeC3PHza4vKaTeUruvmqybUmciNkptGK/+FV18rni/oep
MRZaeYS2PY9Mn57YQQRFq36/13Sj8K7cq3ZiDM+kBYGvTRxRYYPjaBy2hHsaIZdcpnnyQTGvKU9h
cXgVkEcMBsWOh2AIa/rT5vmguVKWSwIYkfBV1VqieKTUKHDswr4BA0pf/3bMR5CetzLZTX77NPi1
GbKcKp32FHXy4R3K9AGDQrjv3UFHal025wi5liiTkLY97IwLKDQv8IJS3Mikm91e7bSMRwsFMfU2
XQctwNujElcRX1h3grNsS7XJuHs59knyiYwEeE14FrLTdqwSaRAesqiYYxjqkbhQDJOnBQGMDwxP
TZYcW1jDOvb+WQUCmnVxPb4rGOkFJDhoHAVCLMFIw+72/0VrEt88XbYmzAL3ef8uUMBWPVwbXlC4
GgWuhJy9PXIHNkDXAe01S2OTPs5QlBJ7HOOK30OT/f84oYjR52sgEbAdHsWCP219FFrAjl1B+Gme
r8No9/b9rTzGa4kYoCOl/OtwjGywxSi83cl3wcheQggq35DPQPAu3LaGTXu/L9sSceOJclgnwBea
s/6tHc8ctcAHKEsjIRwOMIiWGsCkAzTm4fJ9SiwknmcU2fpp9+uuUIXwVvcYPrJveWjqf+aPEOKM
v7fLlShgyU5xNxu9O0grmF8lQO3AQieCqBo99ZWM/NskSGvywaCVjhT+ztIVfAOIeQTQhHs3spty
erTDYQ4bCKu7+6jM2U6gQz9B+H4g+acR0GbN/tiDXvO5SP2WIMl+mSjvun7d7LinuMLNf0zuV5UV
yVvZtw1QTPl629L6Uq76P4LUZQppa+YhZ8cWZ0X/60Jzh0BuKTZpXPQ628QNaIg3VQODQHqgSiIa
1p7HBFRwzI9HK2WUWtacpJEcfE+9U7zqI45Elbwl0tl3PQvkgNWcBQg+UNqDxEsg+K05gNSKJRHj
8aNO0bfbdMgDZjcOBsBcLR+i5z0sSa2ycrFqZJVFPsbDKWG5NKeLvSBrUNtWSQyLEiBa/uQSMEx7
hyEsaq2fwkJciOhRS8wmprJpQgQkMiUJWq/cspD+NE10XaL7gzzVL3e5SDM1OGSgFk+l0vZUlO4R
cMy/kp/uqOGs7zFeLGmVuWLUOxsQnTLg1vVT0QeZYUg5m3kWPf4yRFWViQHHzEhBK/c8nDeOKHvC
us3r0CEdu2i+tdeqxxhAUv6TKfup0DAJ4sUJfNfntm9Xfm4gXdUeERF8KLtkobxrwJmD+h+8pvJc
YCy+dBJz2+1MCbq6qY3WLATkCAb+zrwaFCk1oOcqfALBbO5a6yqMKWcqcFIAiCL30fH1hdZjRgL5
P07PYFT8t6jt3XQbeyOFgdiyWiMhVv8t01nTTmHUej7SXqy/QJ/OfguPbyCOzn4kt5hf5XAjJ0z/
3JsSqqtFhYgNP+yHMfip/iuaMzh16h9VyxU+2toi34unssBj99R45NN2l71O7rEvy+5mHVm3Oo23
WJWhKcCYbGUxFszM9F7T46T3YC9oOEf6zVh7iaDEeHlh4X9AAoq3RtxB+nUlmzfCBeIsMBb3i/lD
VhCm6IcPH0M457+wT8aIFkNbwa65Usu88Sw/de+aiUoQzeuMVxNyNCD2SHM2t+Nf1x3QmT8XRh1H
G3SLw3vHwEIMwz/j9UJTmdJtPvmQ21FxpiDpM702wu/NHZLWHQAa5/8mI3uH34vjUAb4cjVZRW/6
SmKHqwyjJRDIP7nORZF4gbcR2Bb9MkUXFhLHzsK8PWYIsy3splm7Mbq+vVNpwvj+snFFLGzRMiyZ
0JGswDrcCJHvDSfM+mGi48M0DPt/IUnhHpsTAZVWLsjpuQJB/FA1oGlVQZkbxSfCOS3J1RfP5C8b
E2RXSqbDydRPbxxV9A/hbWMSUvt2kYhE/qnELHb2Bi/yp2KTcnq97+UqXLBFqq5+zgt2Hpb+Yvs1
OOXYHSMcVoeNvzKNPjDQ9EiysqUoPAbD7FfuxCS4oQm2O9RNypAgd6KMUIyhhkUFgmQxaS+gbIpd
aNXNHfNGOT1Z+KtnUt/4ct845F7FeTg3J1euBo/pLRNq0aqN523WMWjJFzCk6mpDkKy/QJcNbfvQ
vY5e3Af0IXxnfzJIf7f1+nOgVZHVY5QGy6MXBIw4gAQvzVz3wUXHiT8u+T+L0L1nC5R5qZdomi/H
cDjvjxBVw5NZ/AGIOWvBOPdEDiXUjaS0QCZUTs64uOYinBMkhSt8Eu91Qd8MhkMYW2TcGjAwShlL
MSITQj3lrKsCfzxh4r1Hu/Yq9in0HLI6iVEUF/F/uLhZjPOE0BrY/SiWhSQBi9qUsY2Dc2JnTuUN
SUAbP0BxViUj3HZY4HUwi0m/tphMHPTbKrw6ZMAYnwfYAPIB8dghZ5FuvGL8PZDDJlXWmtR5hLYQ
GuGK8cV/9P7qhg1utBlFk3tq3SEqmU0wWIiDrFHurE0zYeCpwm7oMBd5FKpgfdz33YRdi3YqqnCQ
yRnCGj/9FqUFVOJk6t4WOldRBpwVP7EA5P+xep4VbxQHAbtviPjhvewSnFiwCMwVrCFNBfU2iIMb
Hx3ArIMghylGUZNam3xM5ESyXEUerQn5LntuCMiHalDqZ1AYNuyftRRuTxQ/tTatv9x6t07v29HH
rz2BAgZJJvEFIPQ0BeBxoc4iMYpV3BFi9xmLL+jNUmzrlG+jneFHeCHPGGQ4+XJOM+yw8a4X9S+o
DqKbLS9XoyYvlXOxC2UTfOcWlDg0dsunbvGaVxAeUyRJxp8xIikgmHeRzq3m6eqkvnL/Oq215heD
nDa84yyWqKN2eQSUD34TFpzodr5LLMQqO0kXf5bYsUEX/xBvuNYcIVqGf+K0RgHqXy4azxRuSLv2
1H6mGpawJQM60I5I0o3QETdosau8vFHpNj0grJRYjAXBoULGz3QFHPjwJHRJQ88FbDNUegEUIlxw
ya14wsv8ilU+WuI+g1Az94Ap9O5BQfCIRaD1nYlYTODEkxv2e3XuxPoNK1Sy9CLykU2rIdCH/zBI
baCMAHEYb6l6NSCMYFd1rXabehTCWNPxWM044CHNFGlf9mw47rr2R/+8/xEKApprUaNxISwZN9wm
qyyO7MCEV5Wn/vSrqN+15S7nVWz1DmHYHayOsc9YSP6ijyGDFQEyH/AO5QX7YzZ5lLOvvg6gEygV
rQa12/7oyqCDw0Ok9MtN2A16kAp5qq/PY4VMwSJef5SwuU4ztXGar9S0EVaMFM/ViV2+5vjAOcc0
5FmQWFECkJZ/TZNVSd5jA6LUVad89F8SaiF7QOHogx5apCrXCM9scnR2rBXRzbzbA4jJjmeXStsJ
9u9kpG8hJvwnFArCN/iTcWrEFwwU6dT4aL9mE1KszTdeSPydkeQEdIZ09pv7XUd0u/QhV5EsFMBz
gxo4uVBBd+x3116aawSzsUCX97dEYSO3bSJbZ10Xdc8QpWs39vKszo14bGizkSrof7AQweejmVvX
mUHxUsRUhdh1yEIlTANepWOUyJtmNWpWohQD1IwgBjw/oB8FXCAo/JWpWB4N4FIMfJGTNb/aAEcQ
ovoL3xsEwFIweuo2466y5m8najjXGyixwhE5/58WRhjoxbbJ4UhhS69Alq1lmANOyY3xoDe6cR6y
JiWH7zwDHdul7TU27S8rkWkd8Pac8x06Y/YpQzaylzvTxQmq022RIltt4At8C+bPIJP7r+SIXHN7
Nwby3wuid5oSrDsjJ2H/3LJABgA5g0cAfyVtU1WSiJa80fTlFSjcF8VCsdlKIaXQQ6fuZIfuRA3Z
8u2ZBLJRvZF0uw5sDBNcZYJ5bADKmDk6r6fbp/wvhbD77v6gYg1PeYDlqt9/B1mueWUU/hcuqAiO
eiegmnhLyzYdiqhnBqeP/d8kY/JSUhYUfqfawA+uX9WqFyPIWqNa+89RZhARHD7NAmlXDnnN00OU
tx8UD4Cri5ZeK7Rc8uKJhZ6NNCGWCN+yLVM7PLvkt0QgRQ/u1Lf5CnfiPD/8S7FXlzvOPS4AFMeb
701VC/yHpy1igz8UOzwRS4nCrCgjk0277GvxLgzpsflsnADEB7Mwk5ulCEj1+slJFnUbaH6Fbz23
Bf2BYywoKQKzuVjNOjMYczc5PfSLBK1mefugpX94+umu2wr+EvzqSMyGOPqQWXLswQVTETS/sTey
9Ju4bFm8esbA6LloyC184EocgBP/fOTRm0vH2aIvjwtwtUxKzaZoJHH5u0baFiIujyThtL1wp4QU
MxfTnHNkjfZexEhVBibRqFmYHF9emMY0D3/aCTG7B9Ihpfrl1roS7XO9dM+m2DUBsiAQ+7CopeUD
9pNyjAeTExU8X0oSELuu7+eP7SzmfNa5utr03EtTXfrThEEMtPRZYrzoZhYbdC5pxx03dkOukMNx
ApEhh/B7/Tbg0SeARu7oFsnaRAQy89NcSlnFs3RDqJhYofCfVFbhbNlJTX5bn2KBZqY0E9bENsZK
Yr6vD2T+rez2ShXh8ebn6EwxKolbP8REE17MjlBgoCkQXn+hhpjgaUjRjoft4wb2ZAqi6BdBopD3
oF9OtqAWrRtcvoBZLtFvOu1K5jKwBLKxb4W1u/tCuShp7jmYTQLo95N7FFPqe+G8h31gv8aHsJV3
b+ckFtdj+K1vzIQRQxsOlltj3sfqwmgLDR7fHn0STr8DHMpafRNJ1LbfUvnndf38rmKMzUgTyaIv
/cToDvqBcBV/a34X6/0MRvUibVZGQJtXmpNQ01jYFQ19LEIrmmcy8sR9V30PstfhoLObeh1ZZZuf
mlP5qrvSD8aehQqCk65p3s1lEfHYZWD5W1uDygQRFk9F118PMeb4OuEAeO7TLbayrcqsQa1kpO6t
Oq44ms+82Qyzm1iT+mt5EaKZ7mIbAv68xsJggW94jLXTzIYg9dZ1N6x3l/hq9VihYQMMjpzF1NGx
V5lFCg9ZrP3tRG93WnSA0iOMfMkWHNszq5lnwpGDYe9l5BkqrmiXs8zs0bSFahGG1O2Dy4qXvx0k
owZlqXc7JTnBmf9eetLi1iqLxdxW7nS8a86zYLhmYNpaqNV/zVtp92LqiOu1dhPiE7WoiN7JDT69
MUW2e/jNcfG0KIaohkbU1HCEDqDHry9pota/CWaGrofN/YFJFBq/TD//Bl4Rq7iPtjvBf3n4gw6s
j+g0sUiM7GcZBlCjpp9Ote03wDpZ2QbbQl8qaPFsULlVlrbLLcQrnEGlvTw5p11mp8YTfpFh4txn
zAPoWdVkgLu05m/gF0JikCh4ofoPZwGdp32mhFeS5JtbEO2DaldPUBXVi0/DvX2v8ozq9LHi0pc8
fw2peykJRB7yhWDNRbDf/dS+GtTl5nKkWoEC+PkYN6jQcPhCNOj9paRY9cWnByq2EEP879ie/zJK
JXEmvJDxjKvkQHbQQGnHLdb5lIsqUGXtIZPunUQ9nqQIQpX64/SqR1n9J9af+7r5ciDTatWPGxD/
JXM9n8eqJm53VAteNJ91VMDm9N2CH5HXwxwDTWW/FogDnWRHQi3FoSSWguHHpHbjU/7U8qDr1iHz
3hKo2+cDvC2jHP2GIKa6ab0o9pUlwkJN/lIxQ0e/4pe86m8+ISdZotieLVlFP2ZhpznYTqbrhxqu
JFnYO5YkUuzXPTF4XHStFi2cXTJ6pCpg6+jy7pThZaQyZCne2C2xjLdDI6euXPR8OZuI7f2zSATX
B7PE6sC3U/zetvMuf30lUMrRSk9je5FyhhH6oaBfQC/Qex+JhDQoDf1UcE+DTCirX/xPAZYXIhPg
Hxb1kW/42i8KkLZVN2h7wzq01eMaxjlvO/7/o6Ew7XnWDbxWjkABn10Af+vOU1mCpT3371I1VFeN
nYVyXRPF+NP8Iks4LgmmDd0nUMwKZNl3Df6oKqkxJFkwRCwNOR7aCIN1FGXagyNLxwOnnMUtbNMR
GkUOahzOHSffckCFk67ksuNRCzIfdXPwnSMuqOFddqDyq1eE+fSlQMOMyHWg/bIF7Kc1Rk6MBQqv
DLkeLYpOndeFQy+q0gyibv7CHaJJO2vkHKJ1MQHskbSBT0bk6AX2JgbT9E6kyibcSIOrAR/n0Cpg
jarxrklU5ubCGhlNjv7Y693bTMpoxqM8g2CrfsDv29ZUhTMVQiCc/8iWcKNa56k+rTl76mK+eGuY
mLzB3LJ31hTFCqe6XsfctxcqWtO3ySIxcmm0SgpcD89C5ZeNXPtenAwRA0L/bgH3QOdMdoO9anBd
LH7yViSItas61setR0wlUFWw2Slol7Y7I0aFjW5iUnl/jR1OJdac7vOqj+Ly2roZ+4VwuDDaKsoo
nYzi5NAZX/JpVrs0YZnhnIvwjzfPpzi0P78NjR0b6WhBGfAoGUtQ9vKVINUxJkh7cqRsBJglxBoe
zuUtEbG3zmwOYEIUB5wBelPejmBN4FlJJMZcCnqmL/42lESoE3gFvdyFj1INqEYU5hdhnEmYh+Fq
xdVnVIBF9fVIquL3LeEy+n8eu7vBEXIqQ041rUmdrxtudG+QGUqAyEQikuMlU9seTT0ny9tcdvwD
/zy+G6oqWZo6gNebN0ysMyDtJTiNlVEu92xtM526jyfYNP/UAurcQu2EsP83u4w/HTLwc3xYR6fb
pIlhwt1PH+PEtXImvQl0bZayH9cDTJ6xRGEr+Gb4DWT7eRuSZ/2Mf4c4Md7jXkfVjrfri6TByGpC
YuxRfTsDKkVP8E7Bn3WQxjbUp7jvHjELaQ2bVgcn+24rKM5beHy9CivFBILWbeTpTkSc3pE8/aRt
VsD8WQkUwv2tIFklSISaIveokQ0EX6eQSEGUUK8/qg0z7GJPUMZacsVmtPehHtqK9dt57pXKo+E+
qHvPMzlnC7dGSALpy+wFAn9mxRDAFr69hh6amjWXoeUurCszZYdULgsY0vfSV9bR/aExPqWfIb4c
2wxWoCS4YveHxwNpot7uaWplaao3XDdK0d7vFfzUnFwjqK2zz5rr1FkBoRvd5T7i/zCE1/MtEJr6
bnav8MHF+zflth+gQjl4n/UTWS6sqUQR5vUzSX4EO64BmYTi24hgAcHxnTcaIRVASrxTlTr7FcFl
Q7R7z7Kek0LeDd/42Kj1lAMsRaww4QyhlP+567gIqdGj/jXgcC48Evi20CYu+re6TQ0I8/xeXWSm
CmEKc34gRmoL8OQc8gs99lXnWDDBs91g+xUDsLDAeLN0GaSoEofuPafRJyuUvV0qNAE41SQ+ANS1
xyVHjKmkabm0RNy2rwzvEGQAoOyjbPJ1hQeIsIazA4NjxkSqDbh4Yw8HmfrovoLRoL/4OLGSF+4j
2d1vbOUImMfUOhBqF7vbKEfAv6UglSIOVSCqgS8HAQXikwy8E/OMCObIlTob6b7vML9xB6pK0yds
orm+XYDeTkUjUXvbbYl2WwsreFOKuNRpnplIm5OKcvq/79gXhS3ND/s6IdAFIwbS5J37yda0bsUn
Y6AZWpSpDoJPrSNA8vmebFhQOWXrCh/kHT+CAYcPS24/Xei559O/6kGYhCvVllk7NMoNfXWeVcrM
grQpKL4iABonNr9l9boK0M5EsGolKhZKWwSS+odUiZ3gpMbKnwBW3QoHjn5XLvIx+muyow5Zmx6k
SVfQRxl2Efrr2JEWw5A4lg/rrKWVnoj/ub7zoRSL79IkCwkLUj3UR6NriNFGwBAT7JXgpiSBaHYk
nQ8rcFAKeKoPvt3FSbYkHEsTpUjLUrUUSTSajf/r7DeDiu6Y+V5oRbAQs4kL0hryMm/JwFc9nVHQ
4SYMAjDYhdzsaPXSn7Pp5Q4nQ1Jr9N5EPBDu7nU+8Sz8xQwajx3w6YG/JUVj+32AQJWB2pnfn1Oq
nkJYRGGRZg+PAXoyoYNbcddmLMunYDRlSY5EQJyIG3RydZXAN0GU1GZ8DfnrNAbuOPuhY5r0H6Gp
FkugE3gROxVhIm7kgkagXBCDUO50WiP/LnsLVDp1ZIkuw4g+tEfZTfbiNBf2QLB7nUuVJiRWGWLY
VSusD6NAeTE47V7BoU8y5QooXaRNKAGLbrRJoPccl0ufZCXdYlqSLGSeTza3kLzC2G8EXo/SzRCJ
UbWYHUdHrQ4Q0/xDuVPFRKvKLjIWPgtd0prpsA64UC4psTkNoViMQcyzo337gf0fc4oJDLVxWjZk
S67XMJFfi0LnK7uogRCc+PyH8hWvocUtI6WyAL6/IS8xnNnS017bGQ5zLEVPBT0UvU159Q9aK3H1
2mGK06AiabIEIidcl+TRRo8e0/Juo+GLdFZaYO+VwDYw+1o5qrEyq05Ie1g723fbIdzCTTZFEwbB
4J53YDwAZ88SCAuY2mBxHJyendkhv04DAA4LDwfZXm+ym1FtBvYeb2olwo6taikt7ZKo56KUzpUA
HBt/bwPo22RCyHsNREIKxymZdnaz8R1pOgk6asirYjmXnvguBVYfYecNFTrnIrSV7ogCdQUIteqp
C70H+nyrUAXF+G32n3GbJo9iQb6KQ6nY3RVb0qGhoB6O1MSaxgk9+L+L4Zxec0wjhypZGhH6Befw
8ruXIJ5wbLIQooaqR39M/1fjyqaUF7zE0h0TdnGCE+MPSj1jySf8PJoBP4dYGwRT/LXVHRAmZqP7
+NCTt8V2KrkP7+FBXHTTYd67AMgJS+gBnsHDW/VsYBg3LSO2BLitFi27Fx8hvgNTgxqc29xwtae2
+B/4S1WS4WXI7Zp4RxELyZ6ywPGjey4uGnCYTyYkkouAMIvuU3pUuBCNL5jk9UTr9D+9pEQu8LgL
dd7u4Xg/zOZD/h/suzwhfzAU5s16gRbHq8elMejKWx1tEeItFBzHumHm4VnULb54N8k6RFmwF3op
FRN0UG+WZeEy8EKtFbThe/3abEM6LGhEiEldF20KipAMrPGNcnwHqPcL0VhPpu4BHMw3lrWS4vWm
vIo+6rBAwn8DM2/+55jxetELhLZlg0uNOpRcG28N4yNrSwLGGeR2bNiulq2irPi1i+fNCA+p73NK
Vz9r35tvERTgkh0BxtA1pQXn++vHZW32XfqEcL4moVoGxm77xlzWWZI4YPzA03pKPvxyAZ0GASSo
AnngjLmfiwnGAQsvrluo/UajewpOMCvJkCVj6iNPRRUwnKmLiIn5AsYGc5HGpKyfi21LsFgDy6G/
LzEvt8mg/W8KMz5pDQCqBEinauuMTZwp7zFT6rnUbakrfa2oYFU42SHvMNZZWxRIqKt8VF4VbQVW
oQ0AL5PmyTCqwbUZ/q79dXJLpQBtOGLD6x36xA4M/wETfehdm5rPnemutQrN3XrPDsdU5igTNgMt
DGI5tsKsBV5vDUS1HMpY2SJIPpHGDdemhillqw1RUrHUKsZchpZ6oazC6V+3L0Q1Hex3z9VKhmII
i2VZFh3157+xcjr7PzEP0KxZR565UT5OFDcxLU7zF1m7nHiUTF3H5vo7+xmblNNYVlUR6TP+531b
wmTxAlctb5XA7pNYvUFHiFp4+OmBR9pPQ3VNK39ioPki1UL5hw81XNwoRX16Xt2FuR5TIrAwR7pF
G2orrn790oystiBeoIZTdgp6vNnJoPUwINZZyVKj3ocuUx3yqPvZtCdktIFQlUKygl04paAKc6o+
5Sp8cnEA1HwUIdVkZpi+ZOTwNOWJHy2kWyyv7auOWyPqzOqTAtyaD63lcF11zN2ZxV0XYa2TGNoN
ts8mi+Bb5HglbteGM/74NlkGLysqaEyTXAiPz5FlwV5ZeyUYAH/u6/7JQtDiwRs3ldI+vkJd2Ilz
AE5+NZxcU9EZRu1L9XJPMzxxWlEAV1AvY8BnNEpF+B3NjIpmYPTEUE+LhYQQThLOPmjc2YWFHV3B
YaAgV7LwqhRMMOQhaH1lFDLCFA0cvXFlgYxFkiw/tlHr5s9Ut/VvoXzslcq+E8HNDG1qJOHQiEnl
sgic5GFFtCzkxHNY5XoMgJ+HP4uAlWEK7WeopiOBJFx4ox+KW8j+Q4D2KqH9ouiPrZu011XxQjPt
YA2G3jgwF6X3JeVuIe4bTjOceQwq2O6BuQaiKc725r26NIppuzPkin3cJmrxaTcDvhDJJSEA8Odn
JdSNlcoU5/HCskXktnKEnrAjQaKWaUNvYq5Oq9KViaIBxNWfQbhzW8ECDkmAw+qnrWo+Z/RS9F/J
cT2gHaJtU2cl/jPp1g7v5LnMTEaUbEgiiyfm+bxAG4cr6SQ4NQDm5kTgoBnvjgLeRslrLIAeX5UO
ig0wa6twlWdfzu/zW7PaMmfCr3637MJaJkZVUOjz2U68QNYiDsQ+Eu/DGAIZi2/Sh0ZOv3JAz6Xi
8BqYtunul7XOELfXPxRorfxrK69bPO39LVGg5nsO5NXmpuK2Gru9iX4ptJmg8uxEB1n/diLoUjYK
RSWSKRtqdvKR7cJrMO4UikfnJP4Fu4huyherC7azHQ8gIpXU/yP6UDbs9feZmW1s4nsP0fMxUzoS
7o7D/kBA1oUAPd6FgmJvLK1tras4MBWcOooUfXgvU2b8Zu3QE8kvTv3u02eZDnT/rtL2Mu8zdCsx
dJW1RHo1MTUQy9hZot6q2Fug1m4e5Z2VqbQBc0Lr4BE7T2bf+QDgBrHs2NcOJ040WUJFmP53vC9r
R6xJNyvOWmWqBLWk1uERPATMB6Gw5kQkyGQvHXub5CHBY2AkhTEWaJe6WqmWFFEQNiY2J+C+iW0w
CDn5DeDVMouImHw9upcgRxUCM5YgIFbv+L0SJ85n0/RXsdAW0XCn4FxepRuge/E6lUEpcHtUGGBU
ztvHarBbnozGDbQSjQno2qnBecXEKL4u/SzZDu36+zQwLqHHMwxgb8owE0jNxRSBGq4y4OxNaGbq
TtPnNfY+vcRXuWP5re1uQHmJ0R8WO2bnN4yi9O8UB+WdQBvT7OnqA+jLFbSe2Jd9CU8CLOcztpRU
unbB86VRzeuCN9V5soJlRSWmEAkTSkyjxcFyZRyBfSXEeDHPwNRDbx+NmeZPlGFTVFDrY6BHQQhv
u6o36iRgjG9s227CUNnBZHRfUSl0edy20HklELlU5n62ft+IRioETPrRKPJ6s1Zzt3QElz/JVjOo
Nm6MjF1RARi1jVgV1zcKTexve/z2oxoaoYCHELNNgZljhVtHEsUCxe5+c0AjoHXlY/QpBDgP7ZWB
kdVOu0wu82RjLwOnbeKCW0lQnkxMZiItasuhl8kM4Opa8+Otc5QzpVzwYq3lsDWnWGQDM+x6je/6
o+PauuQKOizxuNScp/GnfQnAX2Pe0EkOWImMIebUWNYZuLTKwF9wRQdl2Ad8cImEXK1sUfkW70UF
Ln0XM4JoqHlTjZ2WIZqreCpARgVgTFci8LU6GweXMDRrlW6/79uDJEm88inwV0J0d4+b1C3ygmIL
VPe+06nYU1IuyKfdWlINaVgkPqTdGv76muTBPYTrAGl7HN3cUzWuLelXaq2CP31mY5qvgc+zNgFM
BKzd7Wo8JH0wrbttbv/8442lDT7oI8VdkZ95aTje8qCLngaL4Mpg/O+ExeznfwPkjsXUOMMb5hDi
7VvMnmX74csaRUZ2CvIZXm6mgaBNdEpGkwFOaEduYPFZbwkzMz3ad3cHzNR5CKzK4gdcnmmVPWKc
q2aSbWizl58ArKEBuLuISUPhh8Yhw/DUdfo/KVpfKywlxSP0wo3nQ7fzpMD3/qj8G268imBd4e9e
GCm10P0IzVpnA/xXqjgsDWFjppgZKwGLNhlRoppHHixBMweMdRfUV9fEzIYahaSyTWcFZoQvpMPo
C8AGTJtbew6T3eWdm4Zn8PHYMXesFC0LEeFGX1u4MPQH6fio2XyEO5ASpxhJC0U2wDRX2dYSwSle
xRZP2u6x+pWYNh6TO+UbSr0sc8qrhZRFp4vKrpahiyNO3+/YN7cKJlH5yyKpNPGZvyEe42f6N6lK
uuQfMW4DVAph5CichuIXX6TvaZiL81jrY5JCqpifgBYnAGgsJP4c6KanXCS2kFExLAarFNKCnJHi
d0htAHMufI0qZAlcQUplF9bktTtScAJX6O2xjKDSiFIibLrelzAj5HPWfYUt+5379gMD+rDeZseV
ZfYfs/UTRDS84STuJ4g0xypu2qrj/g7PzEmvtAAe1VlppXgFxglIcjPZIYy+R6lP2xt8Jh60wN7i
xtvmdMef9wmsYtQ6eSbrzJu72weQC8or4Lh0r69iKoXkPedBNWg3cA9amUs/keOs518GyvCiPJca
qWfs8bZ340iTL/Hha92jjpkSqP0s4YNMHXWQwEEr0cQQxLMBltxsNmowYuDblxCPWZKQ5r/iBX1N
AzAuzPXKGjZ/bw1rYb0ywsNnyckcgbe498KHb1gNDvIjqklNbpdvDg+ZEn3IpmE+wh/rXHo0/keZ
ihhn1tWz0FcW8OkkNkDMEF8oO1kQqSsxEwhzoULiPdteHXqkuyIFoNm+jrccHreT8Iq90S9PS57Q
bwCrvzfPq9zGt93s9J7PoUQkJf0mtJ0k6T+ZuItR2qpXIuCzihnjxkJWVj24l8C7vV/kHWbqp6Dt
gHL1Eu+DVzvwi63wLJUZb3a6m1f1GEVf0DQV3uFJ9fltmm2v+s3+fVIRBltrU9EJ/G2UlwXxTngS
p7JyblnTMop0nHL+edBpGYmZ97UdW7O96+AESZTjZgfqokD+s7mhp26boeiKqUDXaM6wxywCAmz6
tfUPB+f/ATCcByFumAMpiVT5Kt6HbRlJ6M2tTUu4LTjT+orf5gOyJh3iqf6ipqTcUDrG8TQzwC5G
tUtzNC5zSkBE8aLYrmY6oiCQz4QfdmIooyMe1c5Wm4ha05w9FiP7VEpAAUWc1W3TlEuPT0GP4gMq
U14JNONzhPvxhi+dFj4KMcHRPIUtCuSLzlrihRITyXk55OCnU81r0dGC29hjhotjr9e2DvBPE6Jy
T45ClirYfptSVOABBOgs0n5QJOhZDdGZFjZLn4VxeUeBnCrug4XjysXlFk9brLmudI6VWDHm4lxP
4NX0GaVf3yadbq0MY2GOpXk9SArpH2VpfIV+XTn/zOniJr+woNviiSSsMb8GerC7sVdMSCkQIlIj
jIY7rni90hjA86Qat6k+VDMyPNwyCEdVkPwFTXzYZQVB2+cWzpd1S/v6o6G/BoVZLEdkobq+3bkc
c0cmZOOLMg/kognohO+Ye/Ivp33NvFmZWQXKcpzwFAnzcpkyNpaRSZrGZgMpBJY00Vvnx243fJuI
WynTQ3tvDs4xgO5tAtZYtyPrCJReuFU9QhOp8TgsBeousodVgqgNCm5Ssl8lOqo4WgUEAO5NQT5r
jP54afEwfgz/VV4DNVClnKFy++eLYApWvGDPPCfZ2ODE0rf1YQUTQtvWxRfrViGmL1ZcPFAXiS7V
baOMcKAk34Al+1zxzOKYRNUUacKdLj33njzihGSwa5BJkmLNQ5gwk4caqBx7ZicJNpdpdRfF58Qk
g+qn8Tsdm1s1Qp17F3TdNLjfjL2mnxT7f0LX9FmA5eVZAoTMa1PYopepqJ55BnOL8F1mBJHABEPH
AkWI62raO16AU8Tv5CB7RKM3lYYyyMF3Kam25DgbNYPXDiU/IXnVECpm7L2YwOq9NtxL8Kblnuyt
8PEMCIW0AQvS1kfZCeMOJtss/VzsztFKP1utGu9fUbcl1liDns4Z2SCwLukeVk28tOeC0HCiclY5
I8PUzV1nfj9b6MdyegH9L6RbOMK2OC6gxAAqgUhSpPvfCkGdRCHufcMQ+ykWqJaMB5BkDI6WR2r0
geteozIepk1Nr+sJnS9oDbPwKM1DFnaXCZF+jNB3q/94/tg2250UrQDuqtJCLjCsDz+CE44ChdUM
Y+s0tEqheDa6Q8LclDH4+zZBO7UK/DeIW97WiRt5SDfE6mzAxnREL5XZYnG+1IUxIUjvaQExzlOG
0hmJ18pPvDhUM8poNXmvlkeEw7apTw8UQJxvqcj92AJ1VhaLkTFHcwromuGD3RkbjIjGrAn2fZrx
T7KfdK/ZRoOiaRXvGNJZHpageLj3M4gteKqCJ+uDYi8LelCpwJXTyBS87Yc0NIPYsQSitlaGo8aF
8RKVDTRnCEn59uGr5gGzRjBMjNXiprxbPtd03MD87eCrRXJ6SbEQVLq+b0liMcNzx/KoCsWNg53t
dPciUQ2tprMw/O/03Xa54mYKNbdGfvRRTF4oe6up5ozNeYoIDTF7QEol+B7VyqhFtVXn1GO5sWQK
0skFDLFlya8Yg8RgPDTF9gYuZOuDnDQi1V+4r2xaHbTYP9Fvf5syuyTwgWu74KxZRHBg4+/IT2ZU
SS11DpCog0HGNtuhAweDpX/bN558ozODmHnh7Gr9A3KECI41jYQIHYHN8h/I2oysw78sPP6OIJg9
UmHgk2pgYN/tmFR9uiWIpO+LP05MyRYZS284/pAT/FUX1PPDcpv4VDDlqwtGt4jG5I77sfh5zWu3
YiPYlIMYmVGsirjVW+/qTXA4wILZ3lsY9NEDaGlAwqKacNmaDHfic6v3/mVJ+RWalrm31oQFDDTB
C7jpxXgryBqgJDF6oIniuYubMJAoeIThLD6XB6qF7cyzTthhO8xf84fYaSaeIlA6/AyUS9qqaf/U
hMsSBBWMuSZZeumu8iAGXLzWoRn0QDE7zdAJ1HEg+LwXi9wU1JuE6auHnMPHUtsdbea9hdEfF5IC
gfmnnIjIKhu+eCnfeeR59o/CLPXGrEGASLL2vWgQWySHKXeXn3IPoOV2zNXOimIOIdi4areOCdRw
GxRKRSAz3w2peUgXUf61M7taoo8meAaK65kpPRMdJXSwfE3wPF848bR8FJxXMrrzI/y0HoMPYejd
/3QKIjp/Aj1X6o+tumke4ybGSKotQ6u/qexp+Q06viOAiTRCSAGM3s8HYPH2UnN9QYhbD8qsU+Lr
xtMGvwp/DUkCvn7cdWeQ1W5D4zztzjP1/tlYNLIY6OfgKybGPgOYeSI1wDuiCSA4MEvPqCfnCicz
uNsCTRQGc1P1N1fUiyLf7MLz7pHwYRHCUodiH/FUHMEijT1BOiAktZccdN6HdlhyZEQ6tMc3kJsZ
ihyppDdbRzxMuIG7foBKAYcpV6Uf0a/vCnoXa+po2/t2cmghfFGoMNOrq0uNW1vC527L9m4u7Lc6
x0iOoJiKyXIhgLcw1VMJTSFJ5bne138ULcBPwoH1Iis1WAfqT/a9AhRTOuXXRNXVdWsHfjfvhBBM
t7AWFFiaHn12QDtaH4uXAl+3TrADBWLxMJ4VMbjnT5wpyaOi2dPcBZjJ19mUCY/8p7KW85IrnzGt
GP+nvFHAdrUpsvWC2P9IvxIcmaZPb6p1po8zsHSVyH3o2/PUQKm5MsybU32xZmtQWV4s1OgKtrod
daN2LCT2SyjG6HuiI6yaX4zRGL+rUQq7RCrLUS/65dJuQmeNQ8HDMTGnl3or61zyUBcIDJR1d7JK
+Can23wPUUY93xsXkDiAeuR27KgCfFq/w4SEf9DtKJbCST10zYgi2c4/ru3MGMxj2B1XTauDrjRS
EjBVlyBIPMyy2s/U5Uc+YSZQRGKjlM+A9LrJwOahnp20uEvCDpRoUI77oRx43TOLQzmj6ACu0gX9
V2Xu9/LXS4kkFcPBtzN/5Z8rUm0jWRc0EIxMBy4tiQP/8GsH2axWz3BIgTC6E+zFvCe4b6E39Aae
rIHEewBkGQKXq1MpNibBu4inJybZKy2wE6lhxL9jjlLrLoUqgdUtY4uyTBP5i2EiWzywpbsGlOn8
GUwBLz1Sam92GQ5l3WegCIAPlaMf65lhcHh5ekRS2vee3YrHl3r/2oaXst3nDeBcCNru9g5rEOah
yiL2wTO9h3Z8Rsf37V/l1YjajBX1H639uIhAdQ02C5NJPY9+3y58IXim60URTVxjuURkzg9/JP/+
2DaO8iKDAnhxRxpnoauIWh+GiDG6rRqXYNMisI6dNFSZ/zlZMVsOjeJfgNRuF6HLE+L2d6jXXCpu
bHp+a/ruo1rwlD8Et7J1mL0QUOAkH8DWBUzhuF9uT9HLOWu+SYRm89AjpHgZcvtro6rdJq/imybg
UK/iAWvOzxuYaHoSz7kX7o8y1ltwvsKdyTwfccNli4qc70EBpus4NXpzYbi4RnMAWBazfxwnmLnm
iFUeOD/Wh3VcbJtCSrRdxAQR6lDLyFDpnj0Dw1i7K2pUUbERvK95xtJqo2aqabsXoY1ubVUchK/k
3CCy9y+6jYOWPzDlMqW232NUsfVuXWBzu2+dsrE2A9XZSdGRn/7/RYY+l43O7g0SbdtqcEahsZGT
MuPOZyKRtg56f2/w6g9R2odamc19AnYb54O483q3seKRNY0dwL8K4qgfxnvB2s9qOcqeB2TdJv/m
pJdfeiueMjNW9TYwx7G2h0wJrT4IWnuTzJHI4pI5sjUsL4zM17NKCoN3bSl3KF0kkwiKGPeBBsBv
wxN+zF2JaxzyKA4dldjOdMtMLYatWVSy1a6ZqoOiH0AsYIZKJjd9n9TKtIRgZ6sdtR1loQsgRjs/
pcrbNKKm2y5EL+akEmGbXWFoMHzms7iMyjAdDYnAND791gBFupXLr0+K171dWqGqzJGXpeZ3ppWP
rJAjlgCH5Bxl2euaBAA1U6CQgHFhg9qYCEEsUEzYKHcbWZi9/hoPQHDBkWJWykKhexI6MjEMNJEr
Y6gifeS0+LX7Dcm38/Lroxn++JKM+IENaA0NLUmedQ6uFjFGd2I3HtquhsSQxUOq0gKAqS2b9BSP
vct4IGD+CzHHbC+2Sb12LLhmiwQr4zOefiOpB7FW90fjH4JZCguqhtlzI/JZ0Uze5yO/xGGV6Tqd
MtJEqMt0YdXMz5D3OyUzy+rDyh72TrthDxKXABibldg8eowynr18L99Ykr6cJBVMLScBeeu3udPh
rLGNcElcCHC32jLB44icqh98OxwN2WTuiSsiKsRSPdFU4MC2IRphqTFcG2cU48Im0eLq760g1zf+
UAbZLQuckLrlt0hDVstEMMAbetFcypSUD+chz65iw7HIqXo7OgWH4TiEEFRDuCpw14RPQ77PLdBI
hSPlqxC3W7pJTjkeyusyCWMoVDxB2YZro15LZ3I75GBXumCMJwBMNG2SFq8MW4Q4paIGAQF1kcOk
3l5Y/22Syd4fZxCCTd1bRMisoQTrnPIxwgv4V3cqShvd1V2WYdRNeyYY9B/3f9/YygkSL9nWF8r1
C4WHtSmal510TQASsCYOdnrURFlvVVviI1HhgyDhxsoVIyKC+QWnGh7lT/bnNbhyZ728PTlSOBdG
GBh8vzk7S5Ny3x7sjDm3JcQsuZeDZZXw1P+ppM195mtHLIJg5CsCwTTEP96vxgE9jUIg+O91y+mL
PCkVGhvvFwQ89C55a7BAgQ4sF6iMtK3t/GAJJLT4c9HlvEdG4ifE+d9PBVKYZOsIdObYc+Dkt3C1
oHN52itzF4pTF/FvM2NoFgEfGFVBHPLOZ4nlOeYjCG0grpsza+eV2VU1RS3DUUWaFicYcbB4n2AF
RwVTOrc47njoKvbE2SF0crC507GZoAseQ8+b//DLNCq4PwyO0O57wSEA9LoDm5kFEmIMELxBvSUB
9EGxpRh2Imq1xZuBWdM3pMbv9brDpvv0rzbjIULpG2GH+29xG3DRUnJ5vFsyvt/fCI+EpJDl2Uhr
2Up+bvRp+s+EfUh4ZgUlq++OrSC+C2Ck8XygTq6R3PWg6t/vCi5Krg4IqX36SyY5YfXSBsZMgeXe
Li7l4lsYR7rvn7SmQKlc/uASDosrfaWpwmbJwY+8tOfb/JBLE2Gly9zs36VF7cBdaGIMbw1E41J7
vRY7bqYyvcSx76sgxmj2ltmUizpJuz4YpSsEgsv1QI8daK1y6D+0Hlswd4Si45RXHdmMHrWEnLqe
Yn8kt0GphoZ4nK4xHgZu5g6+MRmIBLqeW8m1m/dhG1c143cv6WlZMhQubaundCX3+1HJNvkOY2ff
gxlpmKiqaOIXripnxWMY/jfJeXFXcDQaAf8Qv7mSGQPLDeVup+NF7JaLoOd7GkGz8YMV6t+auw6E
vMfrrKGU6NRkVYlPsSgQ74BtJVxdWKR7cWZRAzim3ee/Zpyjlg7G6b1PqMtQri8ukLj3t7Hn56Nb
3MAQqZV0Mr5KPvdvGmhKaFp6igF4rlU7adCV/U7RYuyYuH5t/KtIy9WU4eYVRy9jF3XK+CnrVCbf
Mn2mEsNY5KLAnEdTy7sL9EYwycOrKINDYlFWZnSJqJzENCml9PW3644UL4ujITV9Sn9cQ5TsJPh4
E4FJcmU+xdu+0gdp8RctfD2DK1tJpF5yG0OnbpdBdvJnBEHrcOUaE8Ry0Kr6jgIonfmv/+PMRuNL
atlzUgAn1srYUoW/vijgFxOTS3X7To42Wynr1K+h74q70oMneEmtqa8ifvQmi63WOQyT6ipEghYd
ddANm2WbeqYkz13IWU1h9VDn99KFOQX6cvk1wd7nh1MGUfzyD5KkM5KWqUOLVHoar48G9SmWic2X
IpUU4tmliw3v1Q/7iYQWI3R5AAFLsqZVuRnhdHmXBlXAcYpT7K3YA9n3YB7mTpDCz4q8URpFMiyD
9Tjq0GvgbTpoQFhgyHeioaoRW+dPs2r1HX6pyTWq4WRUN70NVEVZ++SKMY0MscraTnmnfmFme2Sv
hK5OW7JBJKaglfjR63djK1fVDQwP0DmztD+IilxpEiZCpgwScuciyGYQ3xTzEucN0EGCKM5r3Spj
7eJBuMdKdURJfCPw+6wwFyOwAxH4mBZ2I0Av/0txVn4NnVVkR0mepVE7/xfSU8zdy0snn0iN2dI0
dATz5VZYyzkbhbHnvI/EeAqb3VYuh3fBRuWXGKMjQ+0GNtbsYRodHl28ShYSgmrHkbid/pvHQEiK
PBmARGsqxoNRC4CO28EhPdXPbNqwchJdzVanpHBp3p59WkILcdSX5ZcHJvWrVp6dIViaY5dNTWTm
IHbcuWke5FN+z2ijPpvcZHX/sWsTZyzsQtTk1LYI+q3wBNYDlAaDLHDukQi/eR1BS9V0WQpDqt+1
4Bg2/AmlFrNafeYnmSMl/8tz7/NlZZxCkzAOJ3rt4i2SVB42qA/1l5oR9UDfhU0HDcbMusvVhQH0
LE/6BvZLjAiGvx2eo5EWQL65yH5TGHOQk2ouY15svft6Ri0vM8FQQ4wCZGr09PuND4JaqZGlxKZP
bkzmabY6oo4SWTojguVZ9OSPHCTtnJ116gQIGYmBUgxVD6GmVMIcVelJQFYtq1IYfPE7zjaqrvl6
9DgEOB57Q8X3A4FzoLGR6PiTnXt83ZprP7hmvbRPGS8/C9537edZZXZI/AoE8P7kEUpfywtQd8Av
KFBpO8qFt/POgadWIJwXs4VcHvzgJG2cusOGVgZ3Cb4hJTURKoAaZUUpd5sa8cmd1luwQPqx9dsr
NGxc4FfZogv7uNqcdEdk6zK2Z1HCTJRBwnBXlggKsmHqKrlnTp1DoiKiwzAIRPeAT4pk/7G/mDx9
eB0iMEJKmXV/Vq2pS0YgY8bIWnGadUUnQhK+pO95o6QyjBC3SxH3SL9ZTxFovxj/LuE5YFVDHuRL
6Fo1UumYXNv67NWidVbbs9acbTnYP6lMHBWwBHybnMB2A+zj/RBU05X3YQfkY1N3ZAZu3uwBg6Rm
3gv9LsiblyKNPBS4tkZ1QVzkNqhvjAz0fuyNVzhq25YbLrrznc/95fy4iv7gXdzdMr756IisFV/e
1x5DSHWnvOEUPtGHaDBqNww7xtclXI5qsNsLceqNcmPiTzw1C/yItzSdQVLR3oZadHiWBaJ9VRHy
DXm1iOXLnrOZUh9b4IVIRvbAFRvRnsd/BgT886jugzP/VAbQAqP6zmMt1fC0OFd6OK/LwNPcmyms
rqAPUVWxVE9aG+pylkW/4nFA8d07fQ92/WpqkA8UynW1ZxNRh3dJ23fMi1DcLJltomhjWYHinSLx
m162Q1gMj+oygoM1iI7AKseIE+IsJ8Aq9zV2rDrjL2fKoX3hobddSrg/9uHqDNQ2s+RydywZvmxg
fm9cWvWKLkCuCA5K1GP3PuVcfwwbsXrmKbuRGmpqRB1g224R+/1UfFqgyEkeUEIjFrag5Fm/gZDz
CHCLY687AcHpRBYPoXEB0ylYQHnyjM50mp8PeX0D8qgAmpWOO+YWoNpHlY5xwf+a2vPA3DSmA2dg
F0lxtLa9ixpLx3fDuLZ6GZzJDpu57gpYbeRD9//xWxmFfcAix1DtV4veNSVVH5KEIpqLZ0sB5CCl
6ZeSbYhssOcNiQ9IwoLYVrsOWTFU0c2w62CF1K4w7CbP9/gxHFslrS6usbxPLlZonFFLQNqEzQmo
i0oW0Qv65aGhxscH2uC/rywwgC0Pn5mOA3fQQmLm7HYT/oHc1XJx+5nmShbjeD32eVzXx7ykzcbA
uwU5AQtj4PeYiKKHPH9NeY0nS/g8yhu0sL78RBvX7zcV8Ur3zLEEBciXvSD+xw9TNKJSLB0t8YEb
nKaFU02A/696Gc4SKdaKaqUKi+qN7LG2lDzQz8mV2+j/ho31dc4ls2hqgcO7vtoeVC3dpc70ltsm
5M8vvriSD6+2ST8MLCr0rpOn+RJTT1YHXvxKSaS/ckN+fLBq7dbWok356Jn6XcQd5o3PjpJlo8+6
GOgHMo8E4MTh4TfZhNxgOAb9V3IPoQr9bzwopmF1pjIX4NtCy8lAARAL4gU6c22NgzBWLes4BVZW
nss2YOolMk/i2bOvoiSrlxN8zKnpfj7W+aHJRyC2QJC8SPE7NOFZG3nF8t2/yNhCSKgSzsQBU6XZ
0cdwc0yYCZ6LgESo/DdFZ5yqSxAijeGZTqTcoXTtHb34VXjLWO7BkyKZv3EeiBkLMecMDiSiUTKI
Xm5g1Eb3F2mJEV0qxJ6RJXsC35AYol5Q9IChl4Bbui9/DDpK3lH6vhmb0aOirS7cwL72U5dEHUev
ip6g7uUp/fLaqB/O/BJLg+zu+hYpEeosVd16I34kkLe/qZBO1DudZVfyy9F5R3OSEFCjkAERi/aI
nn7Fr8QdET9LG2jijhL5vHJCcbZwxGFC9Gos2zQCuRdioxZdkDvQrgAaslrVGdtDJgoNs7yHPF/X
qIu3E7YXDM3lo8fuRgEQbJbkLq9VseT7U/F51uxqEgUJTfTNlMNAS68wdFzzREKRbIAMdSRYpfAt
dGi3I7hDLbWYxgzM7OrYrtFJS2xs42jyDUSq4WtdVwjbdpmPPhn4RegmnuikRIZFNyqAqp2Z7Ocy
Q0azWqwQjF4Fq8s7upgt4Q4T+XtqUsWdvqJJSTuPh3TFaF06oH6v99vgjW8g8eu6EfWJsSS6BNrP
u/wHm1bXaJYc5gCtg81JxBjnrT6u3lBMTreITJuyMDJAyU0huwiboHJljP9H4/ShCSOLftov9cu3
aM7EtiQdzq/zt5i7xgHO8bX+FS8GyZdviR190Jp/xepVDLCrmCwW7HTlYMwX8gtr1zb/xp45uk7i
9wn6kBUSu+sV3weTwoLAR/GMCCJAUse4ZfxWchgwsrkdEkEhOodbYI6uWMXpSZpUdnD7ssd3ds3Q
Qe7HyMSHd70ZFdb09KyLzWllzcuYURYe0nWt4AfysGJc2F2EMv9xxZWw7IGxC+xTqKzP8Eg9bOuA
FsM/XAMkDH4SCPLJJdJHh0caAcHN6Z0qpP3WJvxMBoxgRGRAFtDnJJ5FUqNrOwC4dlRkct+5mxOk
J0k+sBfPxpssG7z5760Szz9ywqlEkVLaTtIhGuXGM3ug3Gqgi46pJl+7+moR3RQIDKazBlGjdjKb
t6MB5l8FWAe0ObQiJdwB+jttJqLIAGds5HA4BL/FENHg9czyKfiH0n6WPWdSFZT8805NmnaRQoSY
99SdTugKG6w7XLqAp9EnYtglRi14bIj3ms2J/m68lGU0P14UBnqoVH7+fEtFgSZuDEgCunrtFQwJ
NmNzyIYRLp4BgWOCyHl6hq7FKDnVM1ZdM7xBa1XYWJUifLIa5uhXBkyC6XasWkn44X7/cwgELgXX
iJEEiJ5wPhhnE1PRVfHjeJrqXI6YCWi7Bt52f5068q/QxrHuGEP7xowvNikzHw1q5pYZOIEGRiwR
gLDTM4uLv6U42EW7/1CU/8Ab8BOgjcj3Y4RedX2SrsFoN87m1xCP3YRttkc8RP+lTpP+EjsfoPht
uZYoiYWtYPHoI70bJ0pYdEtKWH93oIN9/dadQCj4/1YFY5GC7F7ZqGJLRnE9MzFSejTFW5b2UsUx
oRebCF+dsllWw/YnCWA+nuXUkcr0XErWlKO0joGq7TgPNrKJi2fStETlxI/j7M/re5dwDls2Wwpv
EDK4Z6x/pCbyyBr0oOCJOMkiU8vkMyKav476C5cAYExipJ+bHOdT1+OcEZTmEzXSVLb23WQUmmLd
+3NrAHBUhgBLUGyUc01hDIKdsyLaJsZMmICkn6qVdL97NI02yP9cDeZmaccCTHzsMOSPgLCwsXsQ
AKzrtdaUZ2YHiAT9DIi/cUurzT0oAAVXn/Ur3cs4UdPMMeP3i6O7X3Xen93x0fMhEjDryilDI3wH
jBzRZFZot6rr4SoTVB6UoHQ68csFeN5XkLnWO8FJB1IQglBKFdQW5o2gz1c0PMP4S8yiERFQm1mq
RAVhgfp+Rd3vWb2nKR21bi0GPZWNHG2WjAPvpTzIFjSc/0ctscIXoRhYifHvX+lUPQm26m1F5Vxw
30NzWGPTEJ27fvyACLJwrvPM1ZEoyTJMIrAcULca+GJ5Lv58sd08JvBz7AHANRzV/tHl9+w9k7Ea
xItnN0v4YtP720v0sMUixpC/AT1w1ruFz4EJnRGvqFOwAzOIy4PH2DmWb81X475sr7sHxa9LkZ3g
HRDHWSxAq3zZ1kR3vvgjbf34v88yNofEfpGlQZPsIiYAszJLGNL83Lu+uqnLVaAZyM49tHsP+kSI
XWteXyrTD3/hzzRBy5fQOlOpeuSHrShYB8Xw8FsZKeusl0N4LdVMEeLfw0j3pF83a4TmFe17kk0+
IhCjrMqPBcAGJJEbt0hF5Wz39vMwAsn5FW2qJ22XjnW6c1jaVlNudytXDCHK6TfrrmIRBGZ9TWhf
z8LUDzZWWgwZ85F5Z2FfpNKpkq4ly0a1rSEcd6aGqZppPG72fnHGkfZn35qQmjLGhevmy0t6uuuJ
haNW4y3DasTd+CSauS43EM9ZhM3/KctHAxpzSaeP/+cZmA75NJgVePElzOhNlOMztc/G8Vgim7sa
UXRB5/ozlF4u8aEZA2y5BRtt4Qk1VxWpnQJ5u6n+pfVDBBOHHQqW6fMlpN13ZS6HXMkhmpUY1g0j
7WDhheCju2/cOjslF67zTlhXw3/012RV2AXpMVtbEI2K17HRpaQcC6/Um3fnWApOOaAXW8BoOqng
z21Mr8Evs5oRw2RXEpdvnKAEIJxjG5C9FwpGlOs0UgOIX75pmLXSC3l2zn5DufvSZbYTM9nJbVk5
/SM5jidrgpg720Ooa9iX/U/LQsRMAPV3IsXq9Ze9IUiF6rJF0nCdRCuRuCp44Wwtyt6QNpYuJzU2
yONaUBaegFZd9wz3imXJYKVhG+8XhbCZmC3rWVSD/db7Z97mCgF2vsH5FgCTZscvGw67yzX14ZoI
n+jGbtGONV+vOIOfF7Zqe3WfMK1ZeZVUIEKZrS1a6QC6lzBTn7wgYujQC42aEAZ9YsTgz3KuVssv
+IV6nFTSqPTXtDNJpB13fNHLKSr9R2YyGvQR8n05MtMDWFTunKkInqXzOZBC/AaYPth9wYNKvp1O
0GAzOeVCSbIw4lChmQZNOfVW7CUA9f4+g35N0ltXZ+I4YD7vPd7SLTvUhr62aIccNAqTkQmNrtwJ
o113bAK9MiSjfPUIg7HaN7tAiZhq9QBrzOdep7VcxiC44QQUF+IIaHsxuvRJjtOlbFxXsZ24uI8K
a+/MFa/zCcgOEjX8iVPOmsyJK/8QIrEAwGDWddYgGwGlA9hflwAi2js6soN8bJSQv94UKh63oEBj
qBLhh4G6W9jAYpGN5l+NQB4ZLm9tXJVOrSKRm+r5ho4ZAWVvzU6/2MJ8VLWTrilTBo+Nlzbs4Fmj
aDDnrqmpiXT5S5vI+OCD7SauvFMlPhurMi0mFR2LODegZQHTCxcSuI64NgaQVL91fHrQvhGgbve8
t5kLPWNdufhFcgWYv2JjQEdyYqxOXP+4N3CAvA2VWh58supgVDVN87W/Or2N4W0lTIUqw4GMcNkg
I5ZFQNgGzLPZ49x83oTeVy6OIV663bJLdJFubok6IIBbqCZwTGaoVr9s5Sm985Cat/jTSt7teS1J
BefCBOZTvjIFqxn801kT121v4BLQrHYZdPpLAkZao7JzSTS4bEQ+oOjLlIOX6iIehSsCzUaBw7VL
2LuXMrzSscVp+xKU/Tw5AEl7tIjVIRClURFo6QBC+kxmkGKjEWOYjF6WRVNwS3M4bocxB5RHYd/h
l95la7htf9mUB15uT5OfReJU5juE4B1tEiVVRubCThxecGm4hBW20KkJiQX0OX2F5Kq6zdhTxYiC
Vx3RonhN3c+WkQhet5MZMNiZa6F9uRK1IeFqy6D0Ju4IpJyoH+sUCeT7N516o5JLpiEbKKbiexAo
1JOGwPGFa5+W4KOyISUzAbGuqY96CKCP1YCs43GOScBDqbjPqZcdFJ0mzqGzz7suY7XEjhj+YFs9
uin6xCYuS3wBu9QQuGXEcrF/KJNTsETZDQyZPbLSSujSb0EYvUeypAkHrsM1lzSB4UDXHd2XZpt6
9r4abrei/Nv1AkWErxrZifRDoeAw71qLJGZlPCfIebtfkJRPTZFIyX12IPMh8E54Zeg4/U3SxBPY
fX+/YukKoJJH/2d3o8sNN4Q7Wo3Ik18G+KQGQPjXug0am8YFF5jgUWycryRaKa4k6vkOZF7i5jO6
y1VEvbKntg7aYaKf95o/MXTL1lHTXAaIp1PlIT1jhrEooMFvt1ST4DFNgnuk7F1Z3ma6rF7TzpAw
zhBAyTWMi9DryMMHi477HGSsfTubjz4Q0r08+MbC94OjMei8sl01rebhrLLAPwILWqJz7wU7S+hi
5D6rFGVKQTPC5TQDTUcpJru+RVAS3DbzsqAyf1I/gZBw3DBRukcAgW0tF+AS9m2h+tz/+CRhBNwX
z1wXuDuS3REr9aGYpspmVcpX1NajJnJAts3UpGRiMY/oq70xJFEK3X5yJFpuylux3XobJK9dW7Ca
Em9lmLgXHZbqEUhuDwkQUEgWB/iPYrogCYcNFLfJ76YjeLY5Y4VYxnvUERbj7uC6LJ1lw0YVwRnT
x4yWhSf/CYjMgfcFeASPVNJNaiVkXugGCj9TotFLJ1zfVhaA5Ne5bEcfYnBfOb6cxvdvs8qSZYSF
Aap2L3vrebvdZSUKFypHp8vRqsQt6FEZQK8qi32ow92w3pJIDcHAn22PkMOjSELlP+tJ5M7Bzg0i
OsDaNXRehBEqRS1bbbMUdNAFsDLg4afg0EaN9qejjfeXmimoCPeFW30Vk9p05t1UOG0o183ofOvo
INR6HiA2OmA6Z5GhXf0rS1I3Wa0Vn3W/ynCfdZYeHdBW6tZ265T4zNtL2WEcgn9wAxYIoS4vHBMy
Btk6S/a6s3mA/NfoTM3RFIJ4WYcfWf/cjNIiaAU0HNl2Mo/Xoq/Kd05AurZTYBsqsHEEm+hqo29V
NrawSLypodikBruoFhaswQZSMqNjO19JnyB7nkRc5rgco8HDM13ZEKt1F3q2TLp5lynw9c8vCTUd
hUb2SyLab7d1W0ERMGr+rXUftKyBq5Lpm5+R7FspNWI63Nxf341VdJkfZboA5v2V0MlDCfGFlpMH
IfIbir0BA5FakCek28ntsjzzdIphx9i6yZBYEIuTLv1owhgMDiz93jtRrQO7Z9SULm2C26zIQt1l
sYklQXhCc0hxrT4RRexghyBsmifwqD79hw/vkqkfeItKPKCJL1P0LoR7DuMEKM3z9MD2WMpySMrz
8QESrItqQRm4FX+Vp4YbseZPjeO9CfnbTewozy/+23IRhu6u4aVZo1ajEREkB0d6hZWuxbiJx8YE
IBKBhGw1MXnl5y9Q1FoKgpsvwQFGb0gyBbD80vRcgCtAiXFqO6xewQV6pY6+dhveebZOZigCNt7o
Si6nSqD0oPmaHtbFoh+ED2z3MLpocsB2hTpE/gO25fzZiiIButllkS51kNeuCVfaIjuA7/tudzjN
LJ9DLYztw2qMwz0FXCaAQLr0aMPjJCaBsP9GXidgSS6K9I2BzrHC1YPKVYeOiwqvfPy0dN8rz9Gz
NwrSLnizvq0D2Wg5UYbRT/7djNt8zzP+C2dCQaq8CUTSq+7FxrAwu3zRdEyIh4g3aJfK6DjwdZH3
+YxN0cFbBVqz/CskZCf6q73bWSif4kBmV1RtFYzQsFikWQHlXIVF5JyoXslSsyrYSFcIAKc0oBOa
ZXJY0dNn+uyf0Y9SHAqzCu/o6EWKN4Iwt1BO1rJmWOBgg60dKV1Ci7L+DkJQJ+IvmeVYGneUOl+7
4VjMsuOLHU5GdgPfpGHUw2xNn0b1MG+oj7k9//8k5OtuQ5O40FFTRXKSDBNer6R4sRSiNCoeuhgi
s35VVGIxT9Zqp4UAlfaPtHRzVHL9D9ESte4r6XwxpnAZbpmbe45luk0A0fb3QdRG22ZAQYPi9RbX
EjhrIKTM2lOykrbvIgpiBKz0o9SNdF4XyQnpdQWEF4tYSQoWer8Sidlan7840zCqqSfBz60TsZfQ
1gFQpU/pLLMjr5ocb++86H7ioUzdRfQCi98afctZwvDbsIp1CZuZEsT8AqiJGtErHDdpepyfpPMB
lJXvBWfEoBVIM5PrUHXcsAawGk1qlHkG9BB5CHz+rJQ0JkaEupuGJfAOSmUKcffDg6sszv4AMbEv
lXuKfAwhbqykcz8fw0ocILCAS0pgZnjCUthTC4HiAxkyQYeiS2wRQUU38hEtakdWxNWFG6FETQhe
9nIoLg8R7ROZCj3XQSZRIa+kyZ1WLu+zhP99C+5zyNQAgjSusUsZYtdzq0ABVIlO/242CQSHG1TP
76sTZaibXN07NjIrTL0aq8uwD3xHUIE0x76SCEWhuQT3YKquc8io3pFBUuXD1pJdAD8J9Euucnh1
aMzy2CK8UTYYq3fu449C5vWF82CR+w3rZM0l30PgIAZXizx6RAmptjGLvXDP9P7D7Gp8rTKMDnhh
8hQhb8qxNa28bVT/h1mSNRM3j5ceksfASiXzHxoGjyTPuR2p4lia6uW4mDnAGLSBz76GBSLlgcJh
rhUUHk3YyiDI3W7PoUhXKPkb0nDvmhuGy4kwW2ccoQjisv7xpc0ximnV+UolVM489yy7OB5cCeKQ
21Of4jGg9ftHAL5ERoOc/InGe4aHd/heFdnIZH/s6Xv+7jCAG96g3mxCwcu8UtxZHQUitytE8fxp
1Bpq4w6QJV2YE50kiPp2f1f4J7z5v++N03slVRj/U9zP7Ctw0C3FHIY7OSaYLJnPX/QV/l8iydna
RbobkUDhwI4/9wEeQbhrGkZNAJAN5RK2dRguZhu+XOgaq/zWGnsBsPl0RJJD8JcLdlZIn4QL3Mkg
O5k7dfmJ6aS7xKDrBL7NN6Swg7x1kLaWITZdsZEorJ2jmiIhxX4/XI9R0mrMSVTHJc++aWvxX8xH
f8ps3CI/DbnK/I1WWx9pnF2Gs4esQRlnbJE4i5+6FwfU5DDoklFcAkdUD2YtJs2VH4jfH754MKPu
k9dV0a74Z5FV4T3djABhy147MihgB4xzbWMCNhtI8QCw9zQQk3aD4+LCcSRKhAbvKdrWSWHqPW9V
tkRBVQgckl26UX1k19e5XS7taTzzWXp2hjtus/kWbLX8qZVFVYOGKjxNQtUYtozc972g1FQhhNdA
xchpXgEC2ycYKPOQH95fhThvEvAU+YI6e6Q+XzISbc3Y71V4Om2yOtUshEod6v6PwTpfrjJ7FnXn
0JeFB1J0csi2yNX1cu3eAlWcWBJ6VVQGiWrCm57GF+GGbFm7igJBSDiRS8alPIK/NHKK3nuJXhTc
hmXYN6sy5Q8xmJhhXawIe5n6XtOVFQIOhM9FfSuXwmZXY1uRrlVbfZyKugri6BCABBlrY37f288C
qvjs75xejUdpDy7B9fpq7mtIhGUIIIv7xLwQ/6JGVC7sKAP5ZzNmkJ7DioIEC3Y/UyAvpFygeyGR
Dqb2mGhDrGyZRzAAItE5XgzX7v6KPkKuL203ZT7hwVnDSGcUNmc0vN2ASD0/RThE93uoDkqUMJAI
As1S5OxHplq3uKlpuK2NiFa4CkiVN6KNRpJCanYGuRktjmJpqURzp0ZBiPZ5N8Fz/fSZAYgURr0y
Fe10bsF08lAZcAJxILJiLvzRha1BTwVcGBHN5pip8IEic9/zWJlaywXwTNcu6uAzEFh3gwQ5aLg4
ApZshyzCFbT+bftVRc513E/Q0hTqEML9rRQDbV8OEpCY0leLha9WmRRIudfH/i8e+jPO7UsN6DSo
WxyVJYlUDBQTeNebaglFYWtuSR8f8DgEjHfeLKgQHeVMEjuwGCMKiSuvgFpc4yMeJAjbkowbGjRX
eV0YJHfMpfPNzj05W2GEud1ZOrh+nttHUrE0Xi/GOgyCN8AyxquDN2SRxgPdN5bnu3lql7XLROW6
Ve9MNNC93zATSBdfHcM6jzPjsf64rphAL8HKM3xRkJShqYUNnhba6gvKItsdRkexKKUGJ3mzMGc4
sTs6hvc+tn54IXi0FFqjxSc2eZqzSFBNXCfu8W9f9P+ZrGzl4V7x5P8r/qkI3iEsKWHAIufrpF6A
LecTJVeo+QM2sZIeDrhDPtm08JCnd/ZMca5gsgJwD/oO3cIBBQea9VPyKCML66OrvW265vLbgWZO
nUba1pOdyjqE6eC2yXUh6ZZ2So1k0Pn6ngldKByhLWiKvvBCUbX2VnwvlE2bMMJdyXzsIX9D0zyn
fxmilk3Jh3DQyLPJGYfwUb9/fxYLacDoEbb3asFPm+mgacpJkLJNi2t6WftkHNl7Q2k7oqCU0INu
UfFY+kTNA0lrJv1NLOt61nji2mUkhxdiXdh011U5hkfsHVbY/NWeANLkh5uECVN1xteGU2NgBvQG
3ZLNUqhIL87+2bCrbqXioa+PB9qEx5WZ1dvGfH56zy3E8q2FU11uE8S/JUYbGAV/UdzXVXcdeHO+
AnHamBHRe9XZTBO/CxqU8qkViR9rozu45v0nYZNDGr9w47x2BZsr6Qaf25ItWKPMjSYxSwS7JrGG
HNU2OoZiP4aK3tawkjlA7g2/zMlNiSuqhG20pR5PqfRwsk01NtxP02urZ6wLSL4635dp1xsTEUNQ
NI9o217FjClFdylW+jUxVttntnQQ3inxhF/kXg5PTFf5Q03rQsTpkGN6UNU/4q8i4slh7xnO/JDi
10TjJyeLzdubDC5CoLgghMjH8kXwdTvApukvt6S70Q/qqnm7stguhPWwRJjk8VnXTvxESeSZK4Qp
s8czr0P1XGGc62i3N8sDf+8CVG7TneIQ1SAa+osqLEyCJhrW0nLEzDP237jkfKI+2b6ByROXSPp3
C6TcUmyqR/ncc8VsSK+d3M+rXLddnGxh66DHfy+PXHw1K2sF/POjrlYXpdAMfsh3mELm5qeLchZ4
mayUgAgOud6CV55qV0nS2QozVGWbo8t7Z2qVoY50FCIu98En1ftxeAah+bvO/TiuzteFmiLVGsKe
LnJGlldNMqWfllGIIvlt0KiP5r4fQJRKYTNF0yJ5k04BuU16sMAkFWDO1k5gUtAdUlUUB1tI6fq1
o7CwBU1d0KlVwBCnToPHvZh6w/FOw4K2G/IuWSxMTXlp+MLKyxprHm2pXbQipjytPqTmysorZFmR
KDTESIMjHV9KQhYB78yG4n7O8hAPjsLqlMb4AXc9N7sPJvl+hbleQdmxJHQVeuRtr/jtwLw8kGeW
9Vw/iJvMPnhfxA7WvxtCe7Tz7Key5YxkaH6NqFr1xfBstemffG44/S57khNdKM1byi2i1YV+Mh6i
aARXl2ZQKZ8yunllHl+RN1A/32TB42Z1SUwBppEIjWLSRrs/SdZotp9Hv1rzVW+ea5X2iX4mwNFw
EFif4/4x6D0nvZukFZhPxubwt6Gtmt/j3rbdMsvrzrroXaAc2jr84naX2ufWkMqWO1q7yFrGVmA4
v9ajIc1i78L/1bICudu7+ejR1vbzUEW5VhPoKbxhwr2Fxd1q73whStjLMP2BrUToqIjiIq5WbnPQ
enT4etf98XC8Ij+EtJylaFz48Aeh0PialG/ZKxxCb+psQCoOTSZPPO8Y87PYv8vmtD8s/zp7ND+m
6H/uExTcanE7AF9QW7iOBpeQ5IE8rIWwKoqK0l49KGees65k5oe7yCDDZWD5WX3PNJZimQdA0s5m
0BrSQke18e1UKfnJ62UilYV0lfpo8xNBYiUNz11JFf1zNK03gzKvI0NWWyh9goswyCBZlsVO32kE
eNxJnMQ3SYMRvv8UgdK4fFHZNbVWlUDc1RbNmBoLCMg81JxrUffePuyLd/Ws61mWDK/L0zCTm8zx
n0n0OLHENnxgfl1nv/INpcg4OKoMY4vJ4k/C1qLwRXCUoW35qVMaaiyPdIWGgBJjqgeHd8O/W+Q+
Ed84PIP+ACbCmwalPzYeGrpEBIi9ydvpDTO5gtWpUp6U9xgZYUKFfTKkjlKtcDgeKmuLkeH0YzP9
xebV6Ldh6f1q2sKrKEe8ulL7QVFYbOjcQSFukEjkqlGNNtU1XYb5ns4sN7YR/xXMa/RupXK1KlPI
ugO7AJCll2Cpnq2+BiAPZeRiMcFs5pfBFKhGW+wkWD9izpnE0sfcoD+Zoa879Dg/yoM8c9jYgEbR
qX47fKnhun6wk42BQkX/Kwzj37t557QZayTKpf8KX0ZDfSzmYfb8j0JO453G/eTSsDwZjM7ZHX9y
nVLQpScR7sk2JQfm5UmfsvgXNZhUCy869PseVUjfSPyNQUy/aDKnQUGpJ+3tgS1RVeZoUYEIOQ2j
TJgzw4sTDpiMUfoNSnCiXAiqlA7BlppUlrCQh+B5rH0XcXu96dgULNE5Rysn9GS7/n5X1erp7wV7
zRT5cpi0ZKhLjkijQMSaLGl4HwTAQ1LoBQuFktfRRi9yvsKa/hhpyhg2hjnCOBgiekhibv2xYQAK
LUGwRvWNRZ/uQ2F81MowzZzCXz9msCKHrnHZtB+etba2XZew6t5tTtAlvtdz1vgoUvDAYbK/O83I
x3XHw93Y/+H3cDGjCtnWvYbKWWzWM/iTegUDF2zOfkVFPTvqUZ1vfns+JMCe8zQLMKBqH43pYNhW
0ZGVUFiKQVccIMnaRQrtwnKWBkZl0QexPgRs5d4PrnDJ/meNvoRsM/FY6A84t/Q/dId8vpYVd0j+
YZblwaDT16OfjqtcrL/V6pEeUSn0JyLSrig5Eazy/EdroGy3ruCgRsJSgpgVOGbOgMr2dac2WgQH
kl3OvH6XQPIJ+IJzwfg3vLWFTOhJ2NxvqcnsUgy4KTAEGU9OJl+LgVmNSigxtZ8ud0vswriACcn5
sLm1xG5QWikW81yM+ONURdWHU9YFzJzcWGCcHczXl1a8xEKakkmwZVjYLDKtKInOkXR5bZsaZDNq
Ien0kPCLq/G4ok9frHtv6Ipne6baAMOoUjrsA/7pFI2hygdn0nA1/bIIjN/evVIR8D/oMT6MxmWC
TFnEjPUo6oNsGpfL74zBjGhIsSG3PU2GT3YETjXEw2rPVcUiaXm9NArM1MS2fhVScgK0k3pksX2V
WUGZAbzax+qORm/nDI1p5FvsAy22scpkYvKLi20B8kTYuL9R5cY3Gw2AW93Cvd0XGjIwGbHUC8Qc
w6NJ4l1FJclikUsXvAHyIDKGO6akLi+Py+d+7H7lj1Ul9rw1gjyRRaJQUfvY37hRCDO0NOgntwrS
SDKh8jJi/+USm7dZgXQQsbsSX9Zt/EeAaNtVAyfgwO1Zc6z6Lo4j7ge3vlFhikhGMHUccMR1Z09R
QUUMYH+zgfVnNL2nN6CjgouY6SCyngVShEzyiXRSX6RzS+dzxG6NJyYKwRKjK7VBW9Flidwq43hV
KcxWpgrcnaQcTIHYcGKR4GD76YkRVNMPz3LwjvwpO7TzBY/aRQa3iqHSV+dJP3sDTDQo+ykffaVM
ARCrcsOBOU2w57Bs2jbbxRozt19R17WHIHyz8REtbBcQYjNIKRxfWiJNgLqK0UkDL7SqqFHrBiqf
6ILlmKQqmpIRGHM+QrjNEEX9Y6214y+P2QqB2NI2KStJbbFHKaFVnVi35Vo12IH2FCtso2wIL6rU
Ieh5wRhQtRvPnNtqHHYxypPagAZehBBzfxqcwlDzEgyeFeVh1aV1OmuQUg3rtIK/t1lvfBAcfTOb
MgqbHqrs9kg8IKRKvP/Y+vRRc5V6+bkOHydqMqmCw7iOJXkbUgOmMHiVBm5663RULfr1KyW9X9aW
Zj5nNjNGW+aIR90+xKvFQR61opjL1Mfj49aPcRkqCWkaFIUcb18hx3oOdOXehQDjxczkuQVJMzqK
0IrwtvHn9qwGslk47nHmaohzZ/+SqZBGqIfYq/rN9TvZo1qLRIOlhEjlg2wazIXonOzDAkrEOeUp
CpZqLxsmG2PgSrhQD4+CZsAogs8cu1g2edynnk+JpF+QMnyQHNiEQs/iD9IAQXG6s0rjmgZ5SKRS
Z4Ul5HrA1qhikHymbpolfizHUJokGXBk2vcej+7Dbp554zLEn9pGoSUmAT3DtLiXDuBjSwtAAJ02
uhX0JJOuC2650l0Zd+vZKvl19hUON23PJljRrBG9Vq65SuBQe/zmsW9QQAhxML0dW55lPerc3oAP
9tLjU3SmXq1ImpSBYWMEaCdwfuKtK962ko3QN1dS3HHTblF87ySIAbQcytzgVurE28A37+AIOUuP
P0sNVTPebPtJ2pLZPcl82VAuRY+kOIXp/9ttSB7TiiGDdykIA/zYnwSA89MyaWeb3q9hBBcSBJ9N
rcwgfQi3b98i1psJhoKyRZb6doEVtIiEUGi8u6Cb6Z/TewQr1I2hqOtZEmeNTSo9evStQk/N0LxQ
msytXYH22ltLXy+GfQQ5JJtJc2Gtdg+SbItUfBgxKufORbX309rdJcqR3UMofs2Pf2j7EYylWgsK
ynOLiKSefkgeUzVECSg1443JgOGPWkYhM+QrYRxUJP40PHeejAfEXQM7tvsbw8zKmNc6m6VVL9X/
6ds675S4b2vEB9xJMHTNzKSIQjL5C7JUH4n88Y8cWEXdOAL8wSLIO6yQXqm5iGZ4432b3rsspOF6
fCmMtaU78V6HgGriaSRm4+EID1WBR+VpI8rQyJs4NoNswxgd3lphrZo8JzO0ks1u7zzvv6jaib1x
uH+32fY1+wZGnQE8vRPyAIWTQ+UllMX4ViJ0vnSc4keTQVGp360g8OwuWPtLxxwjvxUjPr2SwUMG
lLydb//KOjTEL7XpqMDJiLz/E+QL+cJAIhk2fCOpBzNwviH5oakfCkoe+mccA9Bf9MaScOfj/QZ6
RkHm1oud5UJqEcWTQD970VWW+0DaxxFfghXNKehQvViMChcHsfUliKjgEt4YSwKs1yf3WDXTqdcr
37Vigw4YJkl2h/YGIKNcqiR1KA3K+f9M0rgqq+uFO84rrObGSQoZfns8DeVm7obNO0MUT+wuZBSN
lhnPyDhztlyoNrHl3JPyYv/2wXpVyI9L2oI5WjcQA+Um4EvOVXAw6DyinhlMJlkeXvoZiG/UH4II
FfFHzNHGzn6/9ZA6w9SXpCorvSX0WcGFDDguhPUjgt8AXZH/vMsR6qsHV9GAuSueSgxZlN9EA1lP
cPcDjutFEf7Kr7ccCpuxGOVU2ktFdd0ab1eidGb5Lrywon7Y4oPT8xNfHuJ7PBN4mQq2+DtlIbcY
dYI8fTXB/1HQvRY3qg9paMEc25FWss+nVCwITa0jkCmbYg3AVK6B0/PQvRCgq52HOAu0hceBIf22
H3H3LpwUmF59j1JXcm43QOYB1y/2HEGrARx/hQPloqILkLr9N9MTqYqeOSA2qLbvbT1mNXlMud8n
VeMmUm1l/XFw8gPYofhNZGgCz+JLewvc/RFOrJDt0R6lR4QNS/kUgMiQEeVMrk20FxzgSrH+cv9f
o+vSUEGDlc6hYiGTCF4AEjsyNcuO0p5tvmcIbepO2JTWkcaah5QCUzbWMjYxoBQHjV/PfqTldAdx
nISIrVc93zSwfJfkmHnbuiCFmHV3r60Wc9h+SqZ5fmQibQUFHu2IRlKs/BtI93bn6+/6RdzFZHEN
7e7L0RzaNV4MP9kYQaWITFPoiS+nPFMyU+RqhMQ/kXDKXfwJCg7Ydtw3LoNAJjag+mGePQPnEa42
xQeIALYxbs3Hmq0lqwUkxE8bIt8mh9Ffdc+HkgzgkvPdGjAYRpmiFVsatww/LcbI9oriSo6hiE2V
ubMZAdaGW9D1lirLL2eO4h13LZNXimPVPAfoPtjKeuAbHJbz+zHZIItSh37uPjQnEjrw5kXV5RQi
El7WCyy4O1a7tvKMOiDUu8K9YNYGSeY5R5u9Mzar+5gJ4OZwQkRWL9liPPF2QmMHVfGIyoB0vYfP
kW6v0Onjo7hevAe1ikYi50eEFgugVt1mHTZ6UQittM5i9/zGvh9QNE5+MHMgwx5WdHvWxDpZxduH
/c28qYlHjb8wCFNaBN3yms8RaxCQZ1Q6DYFZunpCAa0r8kdV0Bvdhvx5P8ALi+jLD0ZNALLSJOjj
Cj1oo//D13W51k3JuLlZWdxSqep6/lB5qXpFluZgBTLau4g6+UQzsMKe4WGQoC3ATAZFuD1/6isJ
Mn4Lp646S4cOHveX0qw+nSUShO8Euymd122eJiqro7B9wr4XQk5nLRT8DTqWivbx+WuoUsxDv8wO
b2jiAhpBHG69uFWMzMq7CVTYjB25cO/2PJse9hELQahe7fGzFOYaS2rbaacJTBM7X44pizdozNro
+PiuFcpB0i205yALafJLkTzh/cwtB32qVPKCSD17xHoF71dawQKYXUJ4sKFQJ8JQbAiN/ygme9oi
tJjMhAv4bvYyASlk9F3ccqsUAyL9fSjoCT2ynSjL3YFiXsoc8dHtnhIh6/4EZnaueprTe81Z+5pI
dHOK7I81eIWL/Yxn81J7gwFuRxzyrLQthAbiF92MRkITyTDL+yRmgVn/IrA95EmWvnt2m/bOV+H7
eh/Yvb+dSaioOmECbfKs0JPoCwbL0r2m7FDyeC+QZoeAeS7saVuHedBKQsM3Ka5EWXHMQ164WhKg
iua01x1D89WYrtnoOSQR2xMAzO3SaEuzk0SK9NlfiKqWJRk4F9FkNEaqEYiPdIBoZ2DE4Sfg4RSF
kdHIAPmIexhWM9Vzqi9lxMfvxsj02SOGAdFB2IJTi5c765KGkApeS4N0y0DK+h8wWzr6DY45yUun
pYIqn0fazNBxXEWjAibmwnlKD98hSraLBzmSPRxbR66VDNsySbMkDIlgZApQGurDsASUGHGG+Ml5
04WjTSKYBNn9MTjPiayrZ/A8e09DQLEx7RyYgwt6FtHt/iFLkcU1Agd05I7GDFqp5ZE+S7vwvpmL
/7DjxfeHzuR+2k6kNeJYrV1WgsD0waO01RBOvScwHXJlwkCcEKs5NqmP/jkfzGq+njyw8in+AyLg
G5BH3d1Yq6yg0dVAvYtOMJw5mVtkZ2CJmoepgiXPRJG1Yde+q9IUukvDiw8p/pWKsmPcHVhQj9Lb
YvVhK0OUNDgXRcOJe60n+J8NuU6unQD3YHoqHywyPftfPuGLJOQe17nz1lf9sESzpPX1N8Oo9Hr0
HrWD1LAHPny7/rK7jYEGOfGEEhF16Amipq0W+tNZRRcYgU6KibLaEJAPPM91+Jap/Ou+FtHNLk1L
NbCTd2kiLLCetUlssszJWPNABQYm6FCInAgj0tm6cN/FrNk4isQdiwYN+g5SdabsBiBnZ5SZDhLA
n6zCxVmB1EhTv2RmcEKJH2dHEscmc0I4llWKRyfkrPlCfvP3her+YERWBLAdUUdr8DjzEbrIsSsc
iGZga2az2YLmUXmeS+SFdrWQ6g37QZ/PhqcxN7Q0egmR1hadSiZdGSnBBWAv2ZX4yF74EjPEUfA8
11NzKkCJtDOTJBmnqz7vEmAVXoQph6Tv82q63aeTD7G04CgCu95CFIpRu7+njaH/8pj0V+3nUaEX
17W5wlQsnEbuGUwBxUmIjmp6gajZeMoYdgv8EiWy/v9IAWF2MXSkeCbyNp4ZlbINrzd5qbLMcK/2
WC2WCZYw1L8HZFGJrLBOvVu9iswgIRZ526zV8Mi7dIsF0SlvepQ0GYhvrdMcDgWUAHfD28SXAj0R
RZNDz2gHy+ao7hjYYch+ACP31fz07XvnOeR8V/wa3utOx3mRiJLwi+wLIjrvsVKjAetTjdCq0zeM
rP1rZyamVnIXJnCE0aY6+684RQ2Pz/iA9mT20KrGEwsTDjOzX3+2lGu6yqHz22ojw1ismtKIHX+R
yStioRp2TC9zlYlKJucThzhsAy2EgkVDg69gzkP/pyNRYms/ZVuYmKcJg03UuMdEPyeA5DIk392f
WJtDcmTSq2kWfpnbng4wR5bpnDyXnH1LI9oggURawwoVscmySzN50HhX+d5vCfA6Ibswi+pO2ZaS
nARFY0ff7hgqEsdQOUS6U8sMWeQdzVOIynP8755v0rBYSjM2dC3E8GTpZp8Zlz8aWt6iMRKz7nMG
qv/XL6pvlih4yrS2Z5g75tq7Ri9LMcTE2S7Iz4U8iCURlk1Z+6b2b+HK7VVHxl6NThMi/fplMKEk
m7l8IHk6r7EFOxiAQ/LCP6kgEHkYOHnyxGadClk8EgatLPayzzSqtF319Pa9ZSfMSs/N9pejnglX
PQwypc43kH+KhnAdGh8Go1kp3TdJJs4lXghUt/KOzKcP+CeN0rZlSpSxJdDyyC7CMLOLjnlb65Cp
9eT2Yhfyr3CTaw6ArynbTte2f4HksXCnjKavXPSkK13al6SGr0AtYSfDNbthkdBJHYbkDJTjEaEh
eWsA9P7Ne07kfVSWhdlSEsKSbEt6+cChvq2bfWdeBlP/tr9iwtDPrho+SzG3+nFww7YNDPgGGk6j
fhYQgu6/AjH+EMqgQSEAMY5O2lAJqIfEjQVE3NqDb5H6ro4mAgvcXjuoQ1aFgtyCjs/QJdos+qIe
iFPM8IoqI+r59IcwO//gzWVWtLvhjehYA+gLu2Zh16I+wE9fi69VTXHI6FoT3DeqF9FjdJc9LADj
TfHCp823dEnQzNOhBFQzuMNE7b6mtAHteuAs56OjUHa3FuXo3C2zMRITB9nLQNh7NTD+NYXkBVqE
XHNEcQVbRPHMVoXFS7mayPC1lvsu8ky4Oel4YA8yQ2G0Q+/Ku050PYKANSfjiDY+yVL+UPumvLMC
isLxvXWBZstpQXMjueKLFvHfyEx+413+vAaufSP1sN23PY6xRL131rAxnvJOzPomMHIGDXV9OEG9
BJ94tcP+92CRs56peTXCpWc+PnU/1n3vqm8n6X6KzgvBxRjFOeZSjaNdanhLHgw+noUArZUBGtAo
yTOugtJIKp5Q9xOOsEy5Vq00EyACHUMViFst+trT7vuBxT0miAPo4pudrbEGV/sq3mFkrsy/YmIf
+gduuvFA4vUuBNSRooEMwFAnfvrgdh4EmiFWABlhztn5UyQs3VclSvm7cp8GbKceoT3BlXqvWNHX
S5CwINV2D6Z1Q2aBjbpzhrCDMhuI7iMrrQZFA4TB2z3e4Sp8v8A5gRai9XDHDWFnFxsw8TIZOWkE
R+iYz63uY4wOnpsuiWFmTKmrdDJkgOVb35OqhhNacY4ASYLAFjoZ7QM9MN3bXCXyAhTzSFrl5Cie
rwXOVymVjJoLVebyKhjhjn2IgwpFzw0kIWbKucMp82s9/7VR0Kue11lxSUbGetVAhULPchXUv5a5
GDxvZNjRH9kb4HQEhe+lXgIBbqxZ0paYdl0Be4Nq0bFtbQdQfXFG6PMJHGEmNqSeQz0UqBc0lj6K
+RDlVbwMZtIOMxDq097qHCSerHVRzT3OUKSq9hn3uX52X5YAlEQbdjgImJIytt3O93NNTnkxr/kN
t3HsM7KWtEb21UPvvumH7zhq5ILz1mVXyQ1a6/u6/0/lwP6g/tbzXu2QIlh6a0j2wP2CEJxa26fm
mIs//mdc3SITR1oPw+grDW2nfPU99O9dNuqBnjZMppldCbMYh/07x/HlR7ya/RfeDrsbVJHG8Eu6
+/hBQ/RPpE2vl4HOV2W5D125mumI2EQpz5y7oGPg4wGVaHKsPfWT1E0HihqpYWQDNrDj7z66A+eO
+M8xuKwU6l/sW8R2O38nviVXisATHrUvce5VcTgK5HekhRM4hM9AHgVrOuI4INFGApUYbv+5XJnY
re24Ac9Nb4cvIN+K0H2t9Qhvqv4Od4UcjoRzzbbQFeP0pbuEeMSkw3NApxtDh0tGk5ifmY1gVVjQ
i3gauyHWJJgXlmuLQdPONMoXh7XoB4HhED4p00PWCjUq4l87/Olysotj+vlt5B3eGZNAd2kDRsHK
8uR1eUFZ1MNkLa3C6mEUlsJXuBeX1VUwvmaYHxP15MDP+HpWVjylSs+pEGOVZwcnkGJgaanfkBm6
LikAYuP/NZc2d1v4sXcqF4oCrxWs4gKCUTYbMfTJ6DKmRJmRLAIVOSrmQ7ssy4nTPXnaJWezYYw1
+gEBwxTkihnsRE17srlOEhGEcBNsob79lPnK3Q1VQgOE78g5eLT54V1x7qrB3n+71KmKUrIhqAXG
RmdCERseIFJbh7WUapb06BOb6DaHC7whOJhFKaQZ6NWkhMsXwspKdCEWzpMR4Q7AUNV58NbsQKRT
Q14Evj5rhvgYXx8R7zIQk2q9MlVZ7jmQmwZF6uHv39qWS/KuahcK8qsetA+VSDD/DoMbviV24rWx
zUxKUtpd/327Qk8r/SZYelxioq9PBvcsmqhDjcZJnjWBo1Qu1UvV/H/WiZ1VKWqDpeNbVsuIL0fN
AjbmPEKpm7CfjFr++9o/NzGnADL0bAg8daN2bSnx01eQQGM8pW9d+yzCfyW+Gw4nVDiXQYK2MbGL
NtganzWayfbDoCgAORJIRye3lbvZhsvwyCmiNn8g6zB3oJMlcHYmVawVDxxjjvKL0KMbd2lOaJMi
Z0SPRvkc/MelAhARHVKRRTf8y+FW3PQt2oit+GhgyRDBpv76HRza2eWGx9ugEj72EhK9qhTqjvoz
zMB6vlApsIhNQL5HNfXSfhEmgPM2jkrCIa+EfsiMowk5Cj8pgHgmRkkauo1bNYaYyaze0cx/ukMv
OWHznykbr8oQlsFp0tpIUgyugYipgWGoKa5QiM4NI2956kGE8WuGJuUlkTwhOzxoFoJZ5+0ArNwk
uMtyNQBX6+mvdz5qgsQelxVTTfw59i1sKHiSskz3R96euQ+VyB7G78hnITHyS02wrMfYYXmI1oOh
pTub3PMypY0GvcWF8x/ceEbFrpHPrnMt0e3vII5gKHU/IFMNE5PnU7DJajcanyBN/coNWNj08uVY
jkSWGHB3+NFHEQSBEbTytt6bmmQ0wD0Un+XsKIoj+VHz6LE86SknYFEWEdpmAkDbxIxPXtH9Pfjv
oRCjY7jcyk+BcLD7sTh/8Yx5YYYqCDHe+Z2skFEgSGQJcL5J5wKzwzrMjxbtZLOYDbRj7oSMOZp7
AFp6wp2Tu7+7HoAIua4LC6SsII7MatL//P3FIc1FOBh4kaozslYeI/iQy1PxBvnGGRR2JGxHGMLD
St5Bf3KHsJAeT7fqwU4tGWTIKW1gNdH/EMiG79iiJLi0zSm54BjSN7zqd0ScgJHql4e5p8ztfdJO
VdwMLEbWfGJblxZrQxi7fj2mo6p0pIVS56dr1Bgn8RJz+CvniaSEv6P6ANgDsPMvCHqrrazkWm7b
PZ+KyAFzdlLo4oBPei/nzunyy3E8mxmsNqad00LXhv+cP4QMZGl1NvzPLOBlc7OaVAlIkijE9AfF
4v6exM0KY+v1JjQyPaUMAo+05wZu0LkCVlFr8CALnA4XD5aoTPuFbGCpxAZhapCksnZxKMcDCD8q
Ih2h7cNrCnp73W9lWg581ojOxhgyjB/Pu5/kTkQxeKcMPoDSfFq9hB6cNV4t/7Eytv+rvDLb67hp
MnmGSAjFzGQleK/VV/5X60PQfoQKWTXaCnP1DaQeiLP5ch9SVqc+fVC/VhWIk8W2i19plfgzUBaX
dPtFZniJejJurysXgwN5O0Xt97aeB/q075HVFLuLJBiFfwPSmKxE5bj9ZRf+RjdhObT2ahUxiFdq
Zivg9JbERO1uA+Xd2xfKzOdmMRUKvM4pJWxbFIR/3PQnl3s3dxdkhB1cvoCmR/lUlctLJpAVWg1r
W89KRefiWB9bHeIDCLN3NF1o6nYnk+5eYaWiLHNXlKEsopJFU+OBW03DeDocXUl+1063jWiAJlEz
Ux2HQjaS48hwJdnAPn1bDPDBi100dx54Wt5mWwZCeawgtrMcJK3lMMTmTaxRG3uY2+o0bOmouqn1
BP1Z+JKuWoFMF6wBUfvQYYtmzN7WIy2/0uApO9iWfeBv/cWGqxYgzChcAjhmCaxhlwYfERI56ncL
G/kFppMgwkaJat6O/zveJoKB72kQ4BoOV0mqvuHE+5aPOiP2iGoTooHLjvXL0jYWEyb3H4y85i9B
hyKPml9S6lBynKP1mb0jRAoSHXhjDDLiJGHKPjBelDOC2vMwTQ9bOOlTk2Jf/dT5hoDSxAUCWbuT
uMlqRufSSotFkHFSIYdfplIKrqwy5VGChfRk9qES60WFNi7vUlvojvFENJAWOAisaOj2AILAqt3Y
t56tTAXOCbiWlilhffIzW9NR6++8lsQOOTt3bMAZrjo1bWUe+VGUg5U2mNYHGJrHris+9MnqfAvF
jQ12n2Sv8JEPazXKkfDiDbyUflcsz3TNJazqjzWJxsRKSxBVyqDqgpkYwQmoCRyfuN6wkPvOU6Tu
r+BpozVfM7ckZgoHYm5wPQgwsELZ7tkSSUcOdEjN9HCz6VhOi9BLeq1OoGMAdueXxMWepvLqLfe0
4B3EGFhk3rh69sIuyp8/6OhmvTyozN1YBzsAOOZBNttZgp6yxaLk725wv97pIBTo63Sx5VmeJGKn
xEj+mAEW4niB5LBG5kYcfQWYPBeMDjRwv0PhjV4hru/eqiQQTlGs3Ky/amHVP3ZQVrwJr0Gz50fS
gFaHPfSwvm/xANtQDz7xo4p4RpIHxEK+4GUeZor/shBnBbWnEdR3KEc3ZrkQvYil+eGULW8C7zzO
51awbrYTIqrQWZfL8zXWYbQ+X9g3YVJ+CBWbs9k1n8ZzRfZ3y5LTfX9oM2LW6OEhrl8gtI2LX7JN
qNKiYAMqglOpGCKJcerE7i6dmSSOLjIZYD65LGp8JPX78kp/wztzi52h6KDfc7zH/ZIxvpSsv4yA
OOm2hz9K8/U6asj9yO0UKQEtDcJZvuAb60Wtu0md91ST8EFxVZr9Kj2hev1JuUlPWd8U8nUQYih3
gTKJIimRY/y5GXtYukYmNpmqTA5RDm7QCodhdq3LhjEjAkhE0mOE/HZA2dJOOIQnx4GnejXg/HhV
beaM5BiDZFnnvZF0771ybLjWLtLvl+C0SmP6Uj3N6uzYJR6FIbhV3gkuGLBy9yNkgQBtA+INys03
MkCpiwvslOtAFYKDnIrmULNlmkguoKOqRpCCNfM38LDhsbpsNlM2R1osI/zowDkHIUWQJZGRZ7US
eUKXzeZZK2iHUUXFA0bjTQuWRrCaHXgeQ2TsMdzzgyJsSZw8pIDsQA4IhJlVZykrWmftP3KZjIjU
pXNCMVHhPV7vlVGT0lp+p8xtyA1HxAzdKfQrtXrLkENAMZ9tnZI79m9sWKKZflupiczNyV5+fRpf
nosuQX9l3OQiyqzclxhLNCIDpHiyAH866Fp5eGsWMq1msoO/oOpmupWL7eE3Z8gX9hvnpwR1FWpm
VNnky+pyRTQZ+3REHu1PMKIRZb8BQKPylZEl7BgH4lJRB1zIZJ0pc+f87fAdLVZi2oinbV9UIgBy
k7+4l9A6QuTD5r97YYqwOirNiJRH9MqdTdxqUZ71EyLTRBhl5AJRn+jIGUdVzUUa/Xnbp26jUXnw
tQ2OFcUjsfDwPa49fSOSDJtLVGTGPzTyWgf9xnu1QNB1Ry5PTlPfG8ntoc6RsmlLAnQBzvzUExOv
AeS1CgPjaSXu+fe5eMxWre+yZm9o970oph0vs5/453qr6VMze3O9H+QSLPVVPdrjVbMj4arrApGQ
8TwYqaXOR+9+8X39bsH6vum3LFAzvuEmxVaMTmTuu0t1bCDcCkupRBo5PtOELxGTbjlQ++PCuYfq
bsgRmMHgFrVL/XFcAzKzwH67ism5Py45EJuYZm6MwJFy3RR6/SeNuEkJa9HBzluDA/BiQ/GNQklP
tVvsAD/6t200aUhr2RiRs1aF7TTzc599hllBwVnF5te8wzOsQJ3DTKtZgLKIfuGKf69ZcapLfGFy
z6Afihlq2Sx1mDTm4rvh3zVlZAJyaSUL7ioHru/6AV33DURiRIPmxPbffTP2zv6PSty4s+pbmnwm
4yp8mjouvJPx+g6UM0MYmPdl1GGq+n9h9MLEnjo3rXX64Vf/fmdwJ7szEqVOlgnk+qebwqW+U27c
en8k1SAQJgJLFZboYYYF1rS/7D9uQFDngWexu9/s/AX9DBWrZquhmbzo+OXuVV5uE1HtBceSO55O
5HBp9NzjKlvMmz0yk8AoEN4Qjw/K54T5GvtE4QH7StxcKDuXV784oajeCLp0+XQW67Okm5Ltp9z6
y7Rr9InxqRyd6A+P4gZdienUk8P6ewA/e/WatYXS2KDNzeylLtWNl19PGAfSe/GqytgEJQtfeaRe
rLgVp4pirRceW2+P/T7a4UVot+bM9IXc2r4JfsjBA5wIsttZsH4drYvhL8lnzGHJiM5TkkwnVY0m
OYVosESq5C2JBDlY9UmxOmngMoi/b0C4CrbWb3dbVw86IHycyNURqL2WOE0Rtxg+JJwGZpd1dT33
jBhN5nGYWXbGEmaw5ACEx9jOBPaQW1bp33RbgBWWcde6V4nAlLAUweO1f0bnKh5cvHo5JND1v5D3
w54sVn+C5jPzUL/ujoE/vJwFkkitdH8YAEwXxaKeyUL6F+5yaXBUZVMCYit8LevgIN6qqVW4Bvey
fDisAs2d6qVg1+3B/tVtJ4Dhyx+kbyExRwmyHICXzW5n7NqAauChTUaH9Pchj7WgsseeA9N+8B4v
sRQ/hGQ+vJmwbXHCq5H6WrLC4BjpVuv9xGPiP+eu5SBGSqA3J5FLJOj8oa/t/fHdABszRtojh5Vp
P0waasDIjJWWIHe6IH1jvi9xDNaQRimc9B5RirEIMH1iIhiQfxRGDA/W8Bm9p/8JkjJEy9q9zxPY
apO2yPM9/JgDY296Z0NU2SFIQK6RUYFETfmaBoDf9/tZ4vQrlg9RijaP7q/DQpzH/idrE9/+RrgS
Os66360/eljpF+Yw3pifZvW0PJVpgqDQd0GRHRNfvDwwfqC12G6EjxCA6CpimB+NAAu6FJMmPQww
00ABVzfFqMPbmptgH6t82g4qeaqh2V1ff+O9h8VjMOXVHyn2y0SUJqKRheSc+Pxy5Gs1OXvGZjd8
RJVfdYxHc0vouO9ARFBWfiMpxt/DZqH9SD32CrH2NWsA54AloPmpa5guqSZtwmti4Xvdnwe3XnBp
Q0/81S1JF22OPVZIjT94ZAHcFlLoLQJnJfNbCG8XyXLHE4CcoYZ1b3e1TkuPJzvqkL1UYaRx6mV5
6/3dHx95zcEBV6E1ZoAPqAcH+LIid0EDi/X+WGcqklV35ueoFVQpKD7BYWAF7LO/cjZgdSzvXqsn
7OsiDpnU6Fohoudd50VCFwH/B3WAROd+zeHT7OaAipcn4n2w3ijPTHPeV7v+c70ZaYUasPkyPr26
1Appq6MUQCFl+tjdM/IggogrjBnihnHPG0k4sy1J/sCbefYyk7A9+CFk48ZkNcUv2rLMJm5wwiqo
8rMBdyrCjzEe5lgH2YYiMmKZkRS8IfaAC476eOj952XLehad0HWOk5RhgQJG7fqTSZMcbGdewaM4
OsWUTml+xV1QWRgr7A2UOHUqG6OXcHSRcM5PFEPJk1YCrE3hwv8XI0wyhBwNgv6BEl9gVsZ7Vtau
vsxQBJ77F1H3wk3FV3heT/ozt0762rNB76IbUGhr72ra6aWYIAbES3tvjzkn2nwPZQYCKeHjuBQ4
/jXJDI+E2svue71Qo61OrG/HmzPWs1pIEuP2JuDVDcjumKIcP4+J6BDVl1AkFpxhBMvnOJwMIcEH
QdXQpQszpX+zX2lxVSqfeIGzXWNe+2eqP3vj+LzNG7HxLcG89513hsfrLkwyABuW8gEkBP787k4T
Ac3bHx9jrIo2qiJojHDVyI9IUD5fNCQfzE/gW6I1bd/Xlu9RpreJ1c8LXVvQQg4TebsLAKFU/X9l
gjXaMh5St7ZEEtgwWuO0TgsfAB5C38iRt2dcjSEsMQt15L68AVMLBMVVcMxqsl4lCIkAQwmO/w2d
EVKJj+MNBy0GfKT9MxF0uslplRBUMenyzMdbIgLeeZ4C35qOsLYUUKC59B1FwlUa8wg6EEx96Tv+
RixqYsXY2UB8C4V6rlwDdGxbO3PSsN9nrL1NioHLSi0yirHyPQReryUqDVeT6/nvYFYpNzcd8URv
SEB/y0E06fNUqTJT9l0u+e22Hjkz0oHzrou8SQ3/3JC3MYSORZOlqrRF4fad18U2myBg4UyXmxqC
12efZXS55BHW9T3hllJONAg+mgYmQYiFHzGVMflEgHyHt1xzDp7MGIT5llaYbZZeAkinpHQAVVap
QBQHt7CqxVel9l6mEAFNiKT+VfHq8GS6Yn4HqkSD0R6alXgiI4GTvZ1iG2wRsaNurRsHTFohQmrs
8U1LST/hGA+OPFD+t3XNtS6Gk58RjwdENaDmONZhHui2RC2viE8o5mJV89gO0kcmO/eKFtDErKEz
pRRzV1cUs8Q9EXWpVPWTj7o9Apx3ptXQ6m5uF/AwLs3VUu/rPNzq3Xp0yIr4NN3JhgNlsreItvT0
2XZ7MOc9nAERkdzhYxnzc5o1CLqznMzUkdGWiy+8GaIptjwa8xxcHEfcKB4H6f9nZ8/4/RFtvuu3
rqdhdm4Aqk1qK01+jWU3YV7TYa8LYyb8Q0UJwllmWHp0GDWfrNGaMovZjUncVaUKqmj+b7Y3Vj77
MXTxn1KxzfjljxV1O2yPH1sv8vwm2cxwMq/i4SoWKZoTcmkzyCKU43hpsAzaDwzgaJBW/SxY5C8H
NdZBVOyuIxI70GkuMQ8y2hFIJxH+c212c8lLVPsUi0tms2MHeDC5XATA3RtNuK9J7E3qKTbnzjDZ
y3NVDmvBcmlDK8BYx4WRGYKkgXzVfOiIaCtU51MCeZ2YL9Y1d/I3Qpj+rLco1+LZ9jYD0xIpc8uA
pXU69RR6zKmmr10YujC2euzxWTdBVMf7DyNvM1ZqEZLaphE89A3Xd5hrOS7Vm+EVabVE1uNgc7qv
Wuzv8UsyReQWIdDym2/tL7pmE0Bui3YFUHauiLwucQiO3iXgpxFh5mWPlYdpQMyuv3W+a1y53FIy
P4cIAKbXrYjVqEnUGiVdK2sQPDC6pF5yv0rwW5aa///cyQ8K0g2tc7SJugAh9cCuPO/BvLIyaMHA
qKbATdd2f7BYCbOfQ/26FPoQ+ScVFs17vtGUxCGFBKotCg4KCc0YsF0iz+/ITf1aJfB3kI8V3dUv
asRaJXC8k6dqKpN+6PpColV4TRaCore2RX68WGArnj+j+aZ97MAG7eG1zszB+wzvg1GQflf5g+I7
MA7RZ8gzzQDpULLdvhmKluHB2lkgxgqrDO04CdKpaJJeEd///o982qqBzB1wRb+eLI2mE8Kvdvhf
tWNgFRnh/Pfg1er5Ym+fKVl+GxKb3VyDiZmZSAHwgM6PMt0Tv2MJXljr2XGPBzW6XL4H1gjKXkGc
afFjmC39r1sjnOrdPjVq4IE1i20mLIfp0FBmmUI1ijc0xS44/6H9ediI+4T2kFH6yeObK6F/eMOJ
OGJOu4Sxf7vD/RY2zz+OquO8cuRM35vs7N7DWgL4+L3o2IbIghSPRdUxeGXQ3YGhs7Q0diYm1Si4
PtJhoj+j8oW/D2QQkwu50xWWV9ACIbRvd6dzjS4SQne0tV/dFCCtHGj+iWbWlIfMOSbM23usrr3R
P9gjb5kfznU2LxHMvBBzwg4afqphHBMytkOebSax1LIY8u5tIf/5kS9kwtgLH+wnTKpgd7dDsqK4
LuB9gJK7svjvETonl2C0tCA/MImtCfGJRQJpIvrYjHQlnWgXxZvTRY9XXG7N5BdfHZ2PvYpqMBsf
d+x4En/xjbPufjhj1nUb2L3SUKeN5XJ1ILOoSHDaszfKszWw8GNpvyAFBP4izrv68SlYfu4VCJWs
1SOlRXr9vVjKb8ewrKqRRVgBRQRCOsj7J60qxiZXOA9xvrcPpwQ6KZxtyyfoqrLGcoAvoo427bGj
iryCKnEq4pChe2gQcJmp4hsguSn/rX4t4xQCdd8mQ6b7sHXInpLvCKYZnTtN4UrNGRpUCsnK2qjo
zHHPjtjfru1rvWTDpH9Y/woaDsa3K7F5iRdok8uB3toenbkFlArj2EaBMxOf9uKAQNBZkMwO6vQe
upkH9l1s6+cwWHDqrhTDkrbJu6MEtq6A8uC7GmTv4xFpmVUmGw6T5ECFpxr3nm15TMQDlnhh6wC0
21tybodt2ox+aYb5AE9q87O7I3S3+jpMmdZAQN4gHsEla9d6NFUystqPQzhgav9f333ziK1s8UG/
4XftNnC89ySaSX8bqRCsmf87KqL6GGqnnztHS7A4CQp/aXc2o+nZaa2q2QhzoaEEalUiS9pCtSx1
nqEFslxvMh9eCQFYnQ1pEsPPHDIT3nqKl3kPN/84te5VXDdEAgTY8EhDrliW8JyJ40V2/pT4o9qn
BCW9chvemGqpsq8dY1l0VxHe98nLiIuN49gn1PIwzkrc1gQN/dO831iZl6c0Fnjyocbiu/nmZrvZ
ZtD5xQVQPRX1+5wgKO1Nz8dB4Pm7Iy1RtLZk5sStKmcaKgOdPAqQJ/m/pVJzGk+xa4XxkZVo/ZMu
k/ZTbJ95bquyT9AjDK4vc2ZPu+wPzacmJ4cNNRfxMS50FDLH8W4DzN+F0YA40QSio3klSFC1Lc0S
tyGnP4r4jXcisPWR7ocUVMVF6GT43vPq/8VyZXAINtRiBsLcWUIgjW3GUdcU6vqyc630KHsMnCAp
E2enZNIJwlJ6rli70qZVO6hpXxieK6/UAHuEqHTBjrLQ7DcLfNrXCBuc67tLsxRfwsZDQyZZvXbS
NOS1lb7nC+JlMNX4M+z5kuBAisw4tCR8VYWoOzphJIyoxNu6NVrcWtYk/nZlp/e/pZ5LIcn8iAaC
jcx8gNhIapth/tmH65GzF49WyVBJlUrqAEK+9DCgEdtImizoEB82QQUYkGG4BIUVUft/U0fc9zuZ
9Ddb8triw2NQiB7rxA/QUyP/N6KnQQCKTeDAsMWzhZ0UurLNVGIZyPzjbAU5EJrlPUVUqk9HTPKw
6p1DJ3b0bIbXeBXa18kuwfPUrU/KJjCxNpvIYtJy98Zkw5b9ncqxZxKHQx0j3/sOtzrJY0PISVBx
Zeoht7VBNHpWUtlz2h5EqGLPdbdVNiZlgW7dUo0m0bL1oWrOzIgtoY8M4i/GA6m8NU5gQFWzkl4x
orgGMG7wilvHo7DYT1NmOXkHKDbs4pe28zJO9s0stCZo/Ryz39Mf5v5sR8Rz4bca3xcK5zbHpXpl
axbwFD/KTUh1B7hoLgAFf23lL+KfMWf4cWlGaVfUZaO8WnuUhliAAezbMCUKyiN0HV6uO2BLxkHu
0qT5apBpqSldbm275QYp1LBPyNiU4u1gEKPhrUvdGeP7+2Xu1vmRyxA5kv+bxJlk6gZBngKW8no7
9Pb2JWSMUs+LmDYvOTb1jvfy43nrkQZDeng3tL8hR8uGMB8U0k+10DLbW1t+AVIvoygnFMtSv/wT
IAQSIvYsZBm1+fij1J4ezPTjumErIt0QInvRdCeWpEbfzboyEegXXWwWaVBeggob93mwg8OvLkt/
q1OFJcpXeIYuGiDGXnnIWwl7x5HgRyb+k86gfyIQaYzqEg287pWZW6Ymqkl9/V51+02tpQY6oswC
3VJDTGe5/ChqnYZdTc2TjdR4w0i7aPlNNrcxRZNmZRMv5a96/VSK6oScqRI+2trmERlDbhUlZmma
n01bAzCoGmg2u/ba+KTbRBP3eIhnU5QSlXF2r6RVxLtAo7FkorQHtrMo9YDSh6GDKEou5LZ8t6pN
rBVZso/b04oms3IO3skSymGDhC9cpfHp+T2+r1tOecBB9ZNoolV9dWjfWQ3DMwePUPTYF3QKl9jm
D5aU5ACAFbtIqy1blf2+Yy73Zf5yVi0BPcY6/VC8xxPBZezkVVakloXQ+vs6KoBU3k+Ukz4OhSy2
nGmlvaTeirKMLCE8DDjP++DoLfwsZNyVWC46HId9AMUDYD+C4vok8WtzKbxKU2iDvi/uMeMWyX0y
e5iKx94cI6PzCWqi6UkGemyeYFH2vzGr+8CHinmf3LCJcKyCL2A9enGZz1VzBATQb2SNq5pxHsJA
pBuV84HXf6JIgKZmIBhDV3pmN6iCYFcwuukB5I2PiJE3x+GHXkWLL5cXIbtUa3MrzBpQs9Qgb/OX
14ZV3UA3ijyo4h5gnnshdPd7GO8E6zmK/biROaOy5RVoSEx2RLj3A2bTnuBfUT5xtKlNA0tD9i7O
gC3SF4ttKOEwtn8v4T96wTkE2haba8R1ykB0F/2ssmSScRrhy+iT2rBGmsQI1M2Ql35t+CnKS313
iuQoV1dKESZB64V68vbXBdOvkZUpt3Tv9CpG2wwtUwZLhmdQNQHuZxcU6aGMqMX9Kcg8cAIjgJkf
y65QjabPDaFjFeCuWeAQfnAoEUhmWbvPvUjFGKDQnf7R11QZJSU/lqOyLl4vy8qmFlhdZPZFl0MD
I+bkq18BSUClTiUnu39I+73gMwBq9Gb4RoScU2tyE/0V/lpWZu2XPKcL7LMruZj05obnnaL4+YQ7
ApQqUDLW0wGOzS2NwM72EKKmPoB9bt/o/sI28LacOrfqh3NzraXJzu1rmlhRmSMzo3s2FEGB5Wkx
FdC38PDwBaLsYjLMKQHpp5qBO5Ad2SRPfQ4w2052r/HlfhXJ5N8e8DhSEus+8Yv7CoBc/5kWi0ge
9RVhWbCOO09WINqRoC8VcuYuf6cohEc0Oi3QbiPVbH+5LXSA7875h9nyGOflB1tMkbzR/3iwFTB8
vR5xRZffzEAGxDPvpbAkiFRXlU9JfhJv85y5SIB5D+ltrwS+yyd1YxNGPXMN6U362PUJXudKtuZe
Eyy7K/gE+QtTomH2fCkSLcvCqqm7LNzU0jZ9wI7ZmlL5PiCmwA6o6O/t07A8WNgWTQ7CN8xFL5aj
S9OicbKuxlkVx7EdIb7EjZfLj2G2QiP8qzp2wtChzNh5doeXhbMKljS3zh3AIhfTTvDpqZ8kdfqQ
R+oo7e5/ErNLat51trEqFMpnn73KEerij6dvPPUBiUwcr+J6NOmYbxt6kWlmTYoKRkn7afZPi8K5
j7hJ1CtMCUh1g7ZQuNAHjhvBmZvdoVMNTkLgKDJylNh5xzS1jnbWPb6ZfxyXgX7rwonCiXZbGbcN
Jigji6DE7uNIqvESsJbJDRiwt24VnS1bQIdpa6pk6x/kOnh9NNY/0SQuqSa4ZRlRSzUhwrbKjbUc
u5OggCbIyCcxcizmA8Ns/NDFR74WJBxX5bWBl88TDKcU0TXLpMkmDqQh1TsW81KM4XuBVmL2bNj2
IHzekmJr0eQ+dsRkOys7zB/i0iIodXoJEBeIWaYZ4r0ws2Ssnv78jyuf6CxjGSPyi9hhHwn5mzvr
X3f07ZqVpZ7ymoZZeih8wqlP/giaiim4CcMYlcBUBih5mgFjb9Jq6dkDQLNFXFYhruX+JkYAAfg3
R957zaKrhaxAMjKoEviZJ8Q2b0SkxFREPKuQCFLqvOjsgckLjyBAI/8DoSIsYSw1W+SrYYOVJn6u
16I1UVo7cE8kY+FESwA9Vzpj5hD67xksTbfgphbTguYCXfD/rxKc3nDPczG5kEL9tCL2jGx2/HI9
KpMp6fzD5m20DC3VqMd8RxjrdjTr90E0wDdHaPPG+tatYUV67LIF0SmpSjmdgUpPT7jaoCdkuGcb
yK2vEdzq0b/2o2pR+2mdNxMYJumRwxn94MUcj0eVx2Ob7lWphlDJh8tY9hj2Th6qzNWx7v6sypB+
K12z+4RJZbA7GFuV8ZhFGjS7RCMU4IK82WIgga1PS9WvtA7X0jWl+P/5L2WmOxxZCgYRX7RkDU8v
pqI1f3rSecCBzNKWpY4ClrpHptapF/xgflbHeo5x8HgG71KsSxFh28uMM2lETQr0KJvo8dhNuUba
VqG8IUSDRPeS4lMQCnpZdetV7ylvb58D/4c7aRUB9F9ZRZG07JTzgjmbvV0ibhSOXqY3MIXbPLaa
OdjHH6IlI5cJHR6/lOZdeniLELvEzqsRN84hmcOlzNZ2S622GGZANNiPWtKdITUPlHarOtvlK6Li
v0UzmsfyD6WEuOsjRRQW6C990rzCW/qZQzWFmqP2R0LCiz7nlJXv+gKnkMt8qXsh5TZCdV38kgex
BD3+4j+knlK02z8ZjcH5iQonHZhIjj6bBLuTr2mVGRFPB/ibuFT1NqXqtKqoz1Cwz76hT/uHPira
Fc/I+Tw7ocuksYu2mzxKCwPJisMlT3PMQ09MHQkSdGzer+q3xQ7Jiw5ZU14aakDIqTFa6RAcuNQJ
ozkrWiqolVzndbaOGTPqkOm4kxYVdN+mVeWaV4bU2SbwAYLy/3BptHrcpMmKxm7JHX8IOKBl/uSR
TmGHxCU3bANPLGmcPPuWdw81aD093zitinu+styo0iFgO1SyYp/qC6e8fCkmJCruAayaUGaU8FU6
dum+AGKnca6dsa1W1sR1R6Y4kNESttFVzxXFgBXm99mO1Z7N/QoFTxaNISbgSueGuFQZpZuWYSW4
a6269lZ1G0xuea422N+UVc3H0/RpM9M2pf6gi7irbFx8NnxUoqARGSdIsIn8r5LPaXgkqwst522W
wJNX3pHtTPQic4P0TB+fIss2C50klbCRMVpsuQ7S4cY8fR337vqyzptQb2ziYJYXbBO6qRYEipx/
bW7v6Cde/V5cQAjdSrXsCD/c3/FUWcfPUL1MguLw3Yrntm3gRdffbtikvz2twse41GjjiPHuadoe
N2pbk7yVfOJtpUCxtNwrhPToe3/GJwKQ73Hg9xgbeA6FbEn/T74qzqM6qnLzTYU0pgD/bhV+T/HR
ViR2UDkDxT7UjkUKsqNJ5VE2/YjJj/HnianAvL8iw4zGWpofFul1dwDVwLIy/I14VgfHgEBvJNJ1
TlRM4JqKkIqFcxPsCR70s2sZcF7yhyzmIaj409hrtqidjr1QJlFY7IjJ9iq3iJlYi198AwINOlAZ
1tvsA7FcSevyqKHLHrg7Cn0DNfQorfx5ThKdSWBKRA8qfGcdDlvIUsEgVBeHQRB/pOBJzJDAA/X7
qocTAvGaxf8srhYDiWI1/7dHfdz75xBBI6Ox+OqCbhSIXZfJJ/IsszGgiyiM/JSGnBlA31eML0X9
5ohtfmCRg4yoipbc3BSO5PWqjCjFnK+ylbjyhRnYdzvmBg/WrDI/ZI4unvWi/3P+yb38VaFuD39H
zIgpVoPwfdGYGCFs98JJ4gPTD0vIrcF5trOm4cYYQcCVgJTC3h9M6NTifC0ldlLR+HqC0xcks46z
HW3zh1L7v4ACYJ8YGbWhuRxNE/OsuBCIR/ladaElb75saYVg2CJ7WHNbmeCtKcfNGunWg6DWBH8y
iIFoeXGAxe0KIoINdNtk/BZGnIa6i7Hws4Ym0HFusVT0EZO+akk8qAaccZNjIjIT6WeHw886cRwc
vi83UURpFNQG8tcUEu8nuOgI6rA2U1SS8IyU7MdqAqOxrwSdNKFov/cj6Vg35w3eh/PbLPc69jfF
CMyzJR9CH+XQDwCmtWIMpGU2QQiC8nd9rgk/y0Qtjt8Ct7a9Ku5KGVWakMBjYlmb7uO+FXLzoxX6
ugjwKCvRS9LoYFw+Lw3bI+Q7X5ZtEioKsIHrh7VFLs4+C84jZwjHrTQefpEZWE9gCDV8RzAOSsVw
V/ksoE1WTr9fE0i3r9zgb+ReY2aTmseA1038LPC7PBf/z3cPgoSct+OXQeJnMOhinXw/H3LF1j3C
qPcWVkISTzlzLAGvWSxUKmLVictqYpEmP+uwAahasUPDQerqUum18B4oQ8yJKxtJEWgMepNSOfgS
gMcicnXMApGC+eIPk1+iakm3j1IsJhHhOTQo/jJJRESSbEN5ZsOmKchlVmfAkCo4p/LrsrfLyPZC
4lGef/Wak2BfbCb3R+ngt4vsjT1znXzD2ZqE3f+eHBvCEWr/kDdtp8LXjz+Z6u/a00gVklBNsi4l
l66Q5NdITiWIpLGaSjd3hipP+mdtXWrRjgdXHq7D7XFLr1tNzhjTKhB5yGMrtZ7Dhor4pPFTCLfD
9MyxRo9wpxD9Jjf6cgPP/gz+9ySI37sBz37a7IoSf51pub+7bRF9we4Ei45S2q2p580uArV42yGi
ISUKM3kk7c1eIhoZDGkVtR5HZFc9DdUGSckUKK+3EPeoHMhRl+GrLc5VUjqGsiB8vQcr7dMJ4Y9C
qQ8To5uBlws5Fa2jzWf4U1o4qxA3BZlbxrnlPo39OC8Oov8mVxKkZdeZqnm2IwsDGsPIKGrsFDGr
RJU/pLMt3u5ckco8rRn1IL7XZt3eavvTuTl6DW7mA9mv8i84r+J2DE8f4zgoiFNsOaEX/5j3AtPU
X/2+8upiZ0uKV7DF0OraHpOtl81jr6TgG4+TJUPj/xFH6YkSrBJ/9zIEwR6W1L3oXj4ASdMDCmtl
jDHkv6z23Ep0Bvfq4aGoRzJQfzjZfxc54HtrlOXAM4U9prxROiLYFEj/hjdnojDFK5cIG17ENG4V
mPxY7XLOWA2vKoh+lOv8EEI4xMFFikxel1BJCetjOaP/9KkHHTKu8xhttYkSWDSPDsUGPyYR0uJ5
e3IQZtBdUAQTuT9/YoPV8NcL5+41mrVqf3pjCNV+/0JoPHda1BAL7UY1tnAWYvarCCGLgBXQ/H8C
TuXx0FNwOCpf56lFV9CGaTXwM700TrDDfFLty2NCWYUtp2SmgPMgYVupej2TM/b/JeRGFc+BwQp3
p9jhbvcj37O4YD/Wnwz1WQI9ycHtORIpZA8N0SCAEPrrmdoxpm8X1C2jWy+4gF21vww41F+xCJxj
3RHThrVx565IZCs9wx3n4irP25B1lEhu3EXZ5vbQ0/9yAxMjFGtXdpnxiWzGe1ZqEuQUyUcmgARZ
H5GQ/hk0wXxtcN4Kw1RGraUWyklo7/DBCm8E6z/Fm4N4zNEE+IY+pOtFr4iZIHaQtdQD9LwSCopB
OLEcoARfE4pBS3c8hB5UvK3TF7QS9IPrIahUjpNw3PIvxPsU1DW4VRzbt7sKil4cn0tmrBeJu692
DV6I/no3fAoyJuS3so2nLu+YOqrQDCIr5WMKvlpVTtVJ73SXxJTvywY59NXeKlsEzOVP0pY64Vdh
EX1yGKl+ko4FlmybR1yN32aS/grEs+GPvM04SgYft4BQK+iMTjN+ZRtGIRuegpwDH1Thcux+ehMQ
iUlVbBhbOUXalGX0+BeiGRazusARHDrgizvyYWUbzEoIBoDBjFcRdrCIdcHfeMyLT42dqGb82LgR
vj+ia7oEQ6krfUJtYBQyFgWByk3EPTPIJpwyHmGxUXq6oI59o+7WE3KZH5ekMimLe5ZVzl5DTMLd
IC/r8bwHZ4e21ugjjkUEVAKGgSkCFX5Ym0T616PFoz8h6fsO04Sh7HmBpy7s6sjK9jyK5kJtvhHg
cFUmx13SzKtAX5vHKctarjypPx0YoDhqawgDUyt3q0b7WFMRdw+UaoraPDw3zLvEYe0wWMoaMVc8
2z3ApK1YSnCGoCU0tn2vxsz7SCLumU4UllsRvQUsTn+zkd5olVa0dNQqA2cjJhLqfDti4jmTfj2x
whLxKFC78Ate7oaSBx9F97dPH2GWnuUyal0o02dFSpPHodear/KJyvfJNClLyCwwNORpPW8Cf8Fj
qfjCKx04jbQ4GbIzQsqiJ8/WpTfM4AC5gmQpJrhDcQZxJIgeQTDPCPBnTUomsnE3YVicwd9Qttkg
oKcgDf1lAi8Hx6TJc+oO3bdomb32llMVJMIvIEim+alOKa+dXlIOrg2aISbN9Jc2CH3p4DV2u+44
yHqG4KUKzOiKRFwrX8q0qFKPDD3W/kwMeZpa9kqYCchbN36/glx23aJ1BBfAxZ4RwuYXm8VFBXeH
4ghjUR7RQzkJgreML3cyC4kO9YRP7xBJuLEkDuk2AJJCFnN2PufjdAK+CN3+cJbRFJndM0sz9BiT
7Rj4aDEQzOvRDwSx9hmpBSZpVLpWjTb82eK456N6XXJggWFTvfOKXGU8g4DMBg5X1BebXlanmgwV
ok73A5a2UY+z3QLC2dsEf5AzZBKRe3bFc5n0SfBS268ho5yMsYRKCmLSSvK+h9QSWJo8SH0dkPtf
gZqijBpZwnAdmqJ3jSk6MxCn86y4p5kcid9EI+MO3w9KjWaXMo8OtDSZeYYiy+/rwsJzdydAqmfO
z9i8rNFpWO7adLgbKA6g6C6JeCtJn0d8ZuPu3P6Xh0oIAHHLMHxJWEbt+zhGNOwR4NnJIS8mZ3SE
X4DaUeaKSw4XGsx3Ab6RPkMbMy+379bDWwiezZ/mvVwBG1b+cL46NVmlR4uFsg9SI25c+niLA+wH
uXAlRxPnddRczREX/4XI1Qg1wXv0BXmX14DSZOpFvn88YE+hy4CTncxzm0G+yHrjGNjuawClkVbU
fe0Sn9P6bgY9qkBu3b1M060KwGCWmSnVTNB5HowVkivkhC9i9h2EqELKxTpqMMzRK5zdWfLKcBnE
vpZKsiqqp2cFj90Q4mLkkKi/kl44FOfx/JZ5xgMxGiF20IK2P6tUlx7R2Ppi+tNS/pcdcYnTOVgH
AK5zjvn/VKEjluHdG3Hxt1gddGv3EhHFY4ZPX4kO+gwpINAN4MbpYQujBYOq/35jf1l2TC8pD4cK
fEEHyGg3Km0TTCll3TK+BfajxLPmuL5flSExJR4bWkJUndORkE5OnbMMcO5agcdAnddIB7Igz2/s
LZOwgMcO0X5OsOwsQU0NX/Uowq/U6BDlMtfBmF3blkZZ2LfpX0r5096gCXkTUjD++q+bOCMq+MeU
X7Ng10/p5N5sR36udXrNQ68YHc6I1ATUfVXegYmIy6nXOVgVqNPrwKUXi64XtnskqltcXAJuKcg1
ipG4MU2V/ZxtWa+y0KkkM4s+N5y0XoYHjUZA78wkQbwzsIxccRj29iAYIpfLxiTX4ozvxAmbteGG
QI+Gf5yPuh/cYGRJs/EHSt3DcRvQz56X4XlHYtwpPahaq6Q4tnzgKagN/eqm3wSydiLH8d8lvmxp
UsqnAL0SFt5NBNCRMDRdotqzXTIKTBMvOOxzjT+1rU29neSIhzyRVH8olOnB0o6fFNWZFIjd5/TJ
iEZs9B9/vzz9FlOVf6bzyInLk/JO4X6mEoI4FND/bBFQtDb6L4JHNcbvsXOKkAUSk8Z0Ikb08Yhp
mPee/EgYlyAc1fPxNKiIH7PsCjb1xWQaAkcC/aFJmg+r4eo96VZ+5yR18FtyI/eV3VZSEkpmNxsD
cZ5s/4HsUeNDnmMy66Ud2pn0zx8bJNyWMgkA3aZBi2Nd+ufy8iNz9Qs8kT5rggjC9qQocG8oAfE9
x/dnlDV5KiSKwVLN+FC9u6sCvPvzRQ27F4AmoezF07++w9AssEXNGn2zu8IVmUqzhn430f1Eg3lb
FmOFJ1IRozDx8TvoduKmIz8fzlB5/7NfLPSGA2wUscQSEFV1vD+7GUjuAl/NJ8Flj6LAeR1B973l
n/pDYo5G7EVV3T4KepuwGp92xMer8Yc8QWYSKqR1TIsLCnwfU+PQOTGemzgbHN72g5Ng2uWdy+EV
Rq2uXi/DiUzX+xqIpSmPQCnNPDjFnvP2hCyS+K7mXGrtaIdAfTc1TQ1ATrktwBHZUBMogGxDsYtG
JO4PPaX/PEbvGKMsGIBL83pvkna22kMzLU+IqvwTKUvG5ZzQQewaWFllUoly7BNa6CRRmce+Fgd8
YITlqHICqp3Ol8MXFPhXOGPbhqnPL5CiR6QK9ZJ/5zRITyUEpYogV/FrviS1K+3HmPg5zitMgaic
5Q7ue3GhIy8GnXAkFXmDpB06L30C9irDfEQP6mAPJHON5+zvjORxop4KsuXUg9LiCuPAQyEIst2j
ELleWW9u3mIt6Q1n75q6iKcbX2CPGQihSxpNz/ORdlQQvhBzRgZnU78fODr7p3xai5hgaZasVkkK
VvxNLapZv7GguaxhaA9/dJdUZOR5goGmtmZjGU6wjBz2ypvBbAVCkbsIEaxpzUEnsST+EBl/Bzys
g8XHLVhEjqlYyk3LBsuDK1y8bgxN8cJGhisyT7yub5nEnErCs+jHokmawAlLXcF9MtR62QD9nmuo
pnw9+BjJ0KOTKNoEdd1FrmRw12aiIHqCSPtS798Xt8JTq+NvFo55u7lUvxNdqYa4/Pug1c7B92CF
C2VpN7N0cZ1o+D1+rixsmT7+7mjNAgqFe4/qQ1KEGF4DiY4f6wBISA+V7t/BcAZqPh3uLcG9h5Le
TcOvxJmuSE4C2s+8L1xP430TOOyQXMFxLPKHViI5zLsPONSF8kEAGIwl3nP6l2kQStaPuNCY0agE
fRH0E+1AuzuvcpHydJzrl9GLQpvj7s4Oja3Ai1upu7JiQ4sXD9a7mBB8dlIgJQAbFqIslM2ugHYy
PbAUL2MWvnPZA8TBpPH6x4+FqohQQoH6Ud4zXoREnczxnDpHY5IccRXaHUY6i2qLe5gKJWSWsuts
jPO3CF7YsGNgtJStodio2tS5q1x8du8RUVsufk2hqqS27XMVgrBFPQbczIPte2Fljfl9NQGlH57i
LPKuM1OiGFQACV/vg6Hpgn6VdMG7SJC2XMDRMTY+DkrfRzGSmUeDRf4paJo5xLdJczpBovlslu5L
zuOmoh+ITZI0IKloBnZTtAUBZrDwAtL77kBmL293BViUOfdRPc1qUnOqt+91EzSuEpPRzOU9D0n6
App9L+cBTdlnVXGEUX65ogYYPxM2n33EUGkaYCvbEbxBtKcBV8IUE6fO5TchvuR1pkc/es5APY26
ydtZoxlfPbv9maMaTHibdIwOA4Du/o7dvlHfYuQq290FQ8/lDaIhSje8LPqilgSn6Y9LPaYDvb0S
pwpzqXdmYp9PK1UTB7c9+piRNI3RYfBuRFQ4S7U0+m70JJEh/IRR644Y4EJ6NhvZsZ6aLcz+Mcw3
NfbI1PPayz8a0RwZchc3plS4RHUFtrkFKKP5GwSCFVSfBgsYGxSZpqli+5lLCjxY/qpb4O0jcU3h
51Zj58BwGPECZquz5uudZbcrDU8CKqKK37VOm3cMTBiQudn1JF6EJZoneNwayEq2oqfhMnO2yP2M
+tdXMPYGbGN9xIbNRVp1y8lr9z54TKwLPNTYbxHFJXEOn/aRO3wBNIZ41jo8J5RoSmCISVntHFjP
YNMbzzTsaVpCyXvV2YeUJVix00F+GBDPXFTRqihYWSU5Wn92SyAXxo7X06hNRT2ApfmMTRukCDxF
lqNbyzcOc8hOfYUMqXOY9whx4x8ZKDd5RXOB5dgRU083ev+qmkXm32htFsdC22XhBzd4Yn/ViJG2
QIQaaOOBA3MasSNPRVNZDmhAreIKuFwNxQDqdOPCbX565Ck05+UIHA2O8mh/cET0gSQL+diNvpgI
TUOUG1uHI94MHQTQbkpxJeKLQiSwYqZtdaHK1sldRJbQ0Km4MrF4VduMtVZc43tA2s8H74wuY677
wJt+XmuKF3cNfhWBPYMbciZV7jfKh7obF752FVFgt7t5V6I89ft9uesvQWbp2nftlPii0AnM9+ut
D+IuMyM7Kb0+I5Rd7zPMti5Ed2Bc3+ZoXr3MWfUjQQnawVtS1MMKMD7BtvBVbWdUd2pj8+vurCLH
kT0iWYOO0nNq2XK/OK5MQ9Ht7XNKPEaMQWskL21i7wwfgGCHdUXzxNua3dT+tHUwqOc4fKlyH8P/
PfLhtkkEQiiEAEcWmQXnsRnR8WkRnqPtEmyt/6kIzvFXyu8UA0PsbWo02mmAATVpAAdOB0jOF7M6
82yTnOdAy1vGcDMg4eUVo+0XlB9xTHUfFOuAFFtEbXJLarNiGi0XHFNDKHktTLBVyhkPogiBH6iO
GP+S3XMhW/J0Edqt16aperFPcPFi9i+ibxTm+BChEyrnKAKDc5+EwmHu6uR0wttU+17Vsc20p51l
rM86TMKXGoXCFA+nXtlsi2DUxGcZ0HOxfqZ70yRyjdARvtKW7I7PK6eOfy9tMLXzsJuFMh2rQ6n+
77Nc0oroXpXK5bdoVoJtji91RLv917CHdA7HlAz2b0syylAokI7M354FKc6fnOGdafA7m5s5MrrB
9h4JgUpP4bUxDgmz5SwQpm+8fekwbT//AltK/MCKAq0rfR75EswkD2tB3wHbaFB5cp9i+KfwIq3U
2N/9Hq53mh2y8FeU3JffBxMwp+6Eoh13DsLTnVUiqWRIbaQRUTWOAr22nck3SowZx/5TVaRRy+Qm
hWuTagWpX0qpsVCUg+RowMt5rqlBX5Nm9i1VTRwD7DGDsJvSfilhHdYZFcetg5MIYjvLgkXLDTxg
bMyTkg4fvlpLKmM6AnhK3fy7eDIX9you4dVcoF64xIkrb7vpzW2Qjs3yyHC6tm2mLdCQbeYYMP7L
lXTNb+5tfQH7lV9bGJ81a9aSjIF5ZlmB7iYzoEfQ8+o2KsZh5l6paJeM7Jm5IfhVYC+1w0gAWmj9
sHHNBE3a8VbkQy3i/V+YVuk1uNmBX61joTdVDJbUKFlXa2hS9YbVk7B2Hn1y+joBTEsdtPV02HVr
DNiRCZrtwnI7T27XlI7uJbWRbNc8cFOo+Sk9uhZqvhUWXtqubL4lpucR8MpOUIO+C6PLlm0j++m4
/qHaXkQaaTjLvevorFL7DSe3kUDIvnmrGIzhlBME0aMLMW4fUPlhkHpf6EQwoO3h7wlxX3CAZSfJ
TedCM9kYSx0gQeEs2OVLxpGM1jkT9KBoOu290T90iIAmVMbrQnTaTiHeFYTjNK8ioH5+3BgYvxT9
9+BqtJUo+w9Mca7/KhnxjCPaGtaL5oxVN8wSMJP92gA8JYOcfIsfZPD6xKfox3b25EDn98hHXWIQ
yH1dVn0UsUEJKO8rjvDI2P0qqIYGZN2CZvn2Ww0ghzZkOpNjL27AxA2vw1f//2K5xI1k3ws2w9qS
g8SbgKu7vyQrXMPbxpnutDuP2GQLMCgP3wampNVYnuQc/PK21cpLU52TQB/idTmVPqz4bEh0hHJU
b/Pq/p02PGhAT42K8guOr6t7kPl59cRugR24bfrTlA4xIIflbpEIzspte825oIuawIygOs19MpoY
DNtKCP1Xbj3IkZK/kGw0dOkKyYGJBLIagJ3XaRh7mp4Mo6z6yPORUAxewGltbgpu6/qLG3ilHwYY
sIQmcgip3C0xhjzGmuuOyH4vbvhfFtVyKPtsLpa97GepITAQL6YBoMV2C/GnJjpmWVgqBpxk2LsB
rmEgHTHyu3QyzOBDhwmBfwuC4WZzLvutXlZXHQj9Zv41qsH309h1TDnqgsWLxp5ayWWaR7DJC8Um
N0v7RH480HCwb5QX5A4PlSKHSyyCvmgj9zYRMleHAW8N1BCQVKXBrkjh4Fjc7sBrL0mqoBKYq37J
WIUn8FJcZQWIDeoO04EKKTnWeoibDBKI480VRZ2MLsoNNauCTPN3gkvCQv3dL1um626cctwzyK0F
XPtVkF3SDghc7l5B0bATN83uxkod/T2AIOK5IgOQzMcCKGEeHFpZp+EyoEfPccXOUlskj95fIBLe
27zinJ2R4ER7WrRJYCeYUiD+Q3D+2r4qKFFmTk7aImjqshuOWWDQPczKrDp9tf1R0ZwLWSPjDhh9
nWWh8ccx32LvsgAxt7bZixfiRlXB10xOizS5WIDVU+rmYeM5kEKDMt1UD6WURVhOxrDBw0BDl7Um
PZ520/z94qSlNLduoXUjbOypVNHgxtDBHo3aeUxJEQ/Q75S2QQ/V+YsWUtZHFd7rzNYfwBeM3Eza
oK31729Wifj0barXMzZ1GkMMjfGzFWu1MA/m3F8gO2cHq1WjUp6OiVrZ09OqnQK8hNkAl8O8SpKv
nm2OSnCOh1nGFUTMAVgeR4JpduOzQ4uSc/BuJwCuSYfQ0WQ1xlh1GWUxYIR2dAUqLwN3dWY4YdEh
Qaae/MgDMcgsMbxypYzY4ewcymUkavryvrw3zuDZab9Qo9lgdcIQMvMs5ZSm45oGT697eKn8yGEB
F6hdquScW0FnTJsl+AXNSeWVblvKFwNUwxgwBKOcUPYhxlFRphmr0p21vc+5WTANzdbfO5kuMAL3
LR2sfsdXdhaVnuejwBF82nnq1oq8n0m/BV7xz0lcaSmnxAxa6vflYP95wK+U9DFp6Ki4z75O4jY4
7sj6Tc71d8mN8QIK0L8tBU0eLNAbCt8YtAHeC2QnHVbgwp6ZJUfOc1QjNkux4aBGwGIqy9E5lPi1
2pzeNYU7iN6PVG2ADXbiqVIcbPMeXN8VSrTHjvLEmdiiunN1HvDi4jAAJQ1MKlWKkZy+JnxLgt0h
ZNScVhWAwsrH57/fp8WTeTMvsdMIn6GmtVlpWClWC4RsiR/rfjqg5Ltlfvst81uQJohjtk0VDHS5
qRFR7bU2dXX8fccDXoLwKtoI3giJEyOQSq1OIbBZSKONfd2n+ys0alI9duQLzGDmkoAEg8mn7Hm4
c71ATpMGXtx/B0R2Bg7a0YW1tgoZ8nUSU0FcoMzo/R32X+1s9eV0KjsC70o/oLOfIViz5wmVMgPT
YCu9dV6DbYK6ZgyNTNTWfIAPd4XNWIeM4w3u0i6qzT9lqJ8fHWmilBHHRXbskAC79eGG7dw+tdsN
jWo/1o8A6HHEUZSUD2yQHVYVc8m3RpqrnuZBofhmrWwuTiPgmCytFarRrW7qNf6knugRSaycoQvW
p0fSr++3qTlnS8IhYtjcRxGT0HIgut0hRhVWlRArDApqbjV8AzbE3IyDg7DxHsdu+f02BNnQMqiz
ecYRU3XuU15htS4KOJITw3IlmCnOBmvxkT4BvCqsfXWKa/JHnHkBM/LoFEZug+5qYRrcHXaYtbp7
FVNFVGY8lMWxczUQNTgiqUXm7td/zIkZW/I9U4TIFu9bsvy9pmMeYriHP0htqheRLziknNU355YM
knWuUOlWlKOOERG6BpfLt7HP4ZquN29/ZJ0bl45zxLetxkPQdbfT1O045ZCsgHfK4GGFawydUEng
wSSX6a1zDA4CLPwYroM2dSmfKPChJpYvjk/QUS7fathLIbhrUJ5g95v8Hba3tcKxeAvouSd67HN0
GHYdIbOEPK6gZitJbxAiHGRNn1CdojnBE9lzKH64v3GcSeWKwMhqwDfGGvY7zf9nvaHs03xpwBze
2L8dD8KETYIaOeV4A5O6dmQmaUXhCkeT6OGijz3+zYjzEnymNNIvGYEhBoORGh5ODz5MUmIIwP9R
Y5kkwM2qxGuz6qmvR8Nij6bfOr7gCkpkapTVawrtFOT9Jp+kxfjj7Y3oEFEuCLwCG/IPPEaJEQmm
rZWUrSzWQ+CzA9iZ9sPpEYhJwsm6IF3rZvlxybdmbW+5JybnXaQGJRi2oAzHGmJENaS70kOMGCK0
hGYj6Ta8/SkW9QH6uxDLQaO0t1hwsS58CmNGGZhYynlwfSJTclKRZV7Oc41NFinSxwkQyVi44nXF
vqspE17yrA6KQGyd4P3aIIc1C6Q/rbjZXCSwxPfpUa3UkD9oYmDJcPamrykSky2dUpV4VXTkimbg
Wnmn3pp5SY2oJ+I39j+OBmfPTFk5u7PKp2A++C7SLlbZ1zJ5K+uB70w2uagjDunrJ6qxsnnQIdJ5
FLXU7sXH+ioPpo/twFrYUcpGYyVyr/6WpmgCCasvH5RLCtCaCjBQ5ZIaJGFNer00NvJ7pu4goo0I
cYPxq6Z/O5aFFRVJkbFNNadn8e1SSfL7uRjS10VuE0MWFjxGfCqwAG8w7I4M+Y53vKhRpW/XQSnt
/TItMEMpgRRI9aVZ43urlGhG9/UL07urygtrvRuNpnLnLI6rRipk3nUt54vRykH7bBXktuaZCgGr
pXgA8/tMYKTTTko4FHSGQ9Cyi3Jx4X03VewUNIbKbCmrkgsQR4rAQfoIOYN1JZ61d+hYe94Nq60u
JCwUiklenJ9sDuipWTnym0guLX3DsmHpYwPqKsvpTgmSZtYzz0RNyuJDFjLF7gdFh3ltSUKgvJUC
OBXgso2+2n3pgSIFw/EIKY1Pe1YNuhMPA7xyp/QA3ea6k6MS8ILSe7XZBc/6G+juyIbjhMXove4d
x/XXwDi8hOHsUwzjzTboQ2j6g5jAFrZo8zFFzEKCKrBJJmTIbZK3xPXe0GodUha4vO+L6SlWIBcD
eaPSXeFD723rFu8uU4GhaYcvFrraDGyVPPOJ1wegDwd9LH4SW0ApTvIbJD3dZl74WpaedEHPYgEx
Ejj+dlZh8zRlEaNCH6cCEvfJIPHbQ6SMZ5WP0pPtDxLtgpMojf8rlCciDpbYMlkiZVQS01qd4SPM
NFxY6AaaNFDhI+4r8F4lVlH5RPjsxqnQw+J1w4uQ3XBmsyoJW7SquhCvmMc+h5D89vySRrm/rTML
nnfRLWLTlgDxMcJtgl5dpjzP8JScn/NriJn6lbOGpH+3O4GCxeqAJXhNgggB3kkwAJx31T0v92hS
k+4R3rNmWRSeFq3JcaCbEPXBflMSW13kmH4JbAWIS28ztL0e1mllqi7yCJx7N0QQOiO3VB4K0yEU
jHRxOLHasuLBtVGF21WdqdY6uZfo1S40LsvlMpCeqDRHbNG4lyehG+UgHM4NRHcVxlAZ9spTzZ6c
xrQ96sdfBRI+x5SqTrrX55K6OhagaWyhInAKZCUfZ6JNBx0in0NheIM7f6osP5JRZVcV82s9V0g0
Lty4H07kzEwU74FIJRyf0Q7omGuetY3jBJg0KKSLO1EN6Jnbe9qqz/25enwAOHxgGDzUGE7R0rzG
3uVFZt+ERS4NF6TNqYJ1P/ZeB0aFv55ZNlVb50w1MSqhs2OCtq59fxCSFJFI7oeYFL2nIySu2/lu
zYH9oSxpAg95Hc/vSwDEHy5/LgsaRNPCm5JCMQQCpRkqMj0E6Ze6YqPQZrA/lBbLziP3EhhUv/IV
mykCcpDV6E+dBb/DXxH9aMKChA/rE++FDvMeimS7DpgG1+ID2OSmV1DHnkIYKEl1JiWstvq6wzVS
Las6lWk4uJTx0Mer5wIy/ZEzZJXN0OOWWjDiQIsO1qz4AJ8WyL/ZO9Kft/L4r/tPflJ4gFl7QrVT
sjvaXLf+8WA1bs9H8xSrYyZQum4KskEwPMzXiNsCfYXIomqp60NAWWAyhPGNr+Ud8FCYhlVUD6KQ
tFWC7CKtuvt/hirGGcEPiZQzh4PEjFKuH7sSOl5H4zZG80loeLXDG3dUCBesReVXlaBWTCcWYEsl
u2LjoFWYCQK73VKM6YgaOTYr4HFsrmQIoBCGVkAoTa3zuFi11lzylXDWwJKMr+NtIycimNIDnlXm
VW/m3EeUsdpmk7LRAK8M1Xfo2IQnihbRU386fBV/+ee58MhKMq4rw4TwWp4ic+nkCKg8o7FB5Uqs
uLLAW7nsiNEPXMpV4FC6/nX2bPIWoB8Ch0+mdAATM7Vl1VrwGkWxRVwmUcow6oKoqr5piXMjfEm5
u7OhOxdm2398eiOttnHgDNyYZHt7YcU1drmUOX0oGRu05RL70PjWlb9al+RHIJdPJMK9nZqYLXng
EtZ1jusHiAwqflvMx1FXvMVFKcTu9MTQpRZLmiJmGuoYv86mUaAX787jEOaMweLnbncvKToZOzup
t8ATeRkNJEOSEezOxJ2wxCYJN9q5uum+SbN2V3fwYoD7UxM2H2B6YnkMM8h72GqD8ZUpmN/zA7JG
lHofD4B10otvuY5lLthhVWR6SoqvheBBLliu8yq2x0R/rhG9PllKw8llQz94k7Nl8ez+yyBYnlE8
WznbVrH86VSIXuOdzvGvly+GmoOo/5sqZEJ49jRm82Dm3qtCo8XUWudOUI0a/pgcKeXss5GpUp5A
+gEmEYR9YSQJk5aFo1WCmfPbImCD8IEyyBlwbzwHhy9vTymArMUP2VFkYmWomWNq3uQ98U4JP+B6
/zZ4N1GRD9ZkAD7Vl6T0VActJeGxbBoylvMBlS+jBA/kTPlqAzkZbnKkMX0KuI06u2ffIhl+PfLF
ANVdHDH4uZfG0Y3wgIK+s3FD5WqeCX8T343fD/S4liBn4wkfgK7uqR3WsadAQS79IAsmyOe4Bll+
qMq6csqe4L8ccuzstGmaY5HQc40AiRWJNMpbzWZ7FoAD588Rr3VKAVbMwrLPndSY+qS/q92KUgJX
IgsB8+nBLAqzU61llXAr5io5iVDqLx5Qy/0cCOcTO7as7A1RohiHcHA9vkD1kvwfCAJd+fQUN/2v
Ilq7otLUwfRb12q4pIVRug2zVK511q8CVNxZC88PFWwiWdVIdnGshUSaz7vqLa9xJqU6IX7HYtTt
CuBQKTsYxiok+ZcLC2RocrnmKGKworo2QBETqQxU6zNAFRT4qIKZGThEwrcIrFmOpii9smX+aloP
QlEl4BsQR0IbxGdwzWXauwF3qfgfcPbMPC79jhNdUVM4PbuhouRUWFaH2TvYOHmBmrK6ateL3FcC
jB8g5Ga4WINDhVZ6XenjsqpLkM62nIkz936eVdrZoHwMQbPA2udTYE7hhFRc0eL3vateT0JaB2+L
yRcXICvHhVn5mRRh6OqRG+XiyA4R30prTTZW5QZFX68Kxx1Ud1fXhF7VDm8p4HU/DxUYE4lREtol
z6nANmSTu2fzoXvAUGPqaDJlGDWGQmqpTbkWMzdn/3eD3jh28VfRAzSwXMSW1A4+vPRDje8ZxCmE
+Ve+p1/vXjU32XKzghazV4u0Pf39IOw7rTvkPVPuAKRXqfechNT6cNAWZ/xa0wH74oxOtRXWO8lr
fu/atNoFngpU0IgXPAu6GjS2tdXfnEe4erxOreusP10QkvKrws5xlEwYeonP79PleNHbsyNHfr9J
OgLzlc67fNYejJm/ZZFwa5XIxepUBxa4j3RvbCAG5BNYMnDDpOH3KRAtobEzhmhusb+eNmgFOCyT
PCqHvb8alL2C/wypWYXMS/WX67znxDIgrfq9Kfrhc34Z1mGl5PeBmPvMCoLu6/3O1sTqEL3NpAVa
coYibS0MH30C/3vqmeWH9uz/L+rUQTHyUeWQ37hFy1J/K0+AEOX554Tz0fPnN9Mb2IFLlRr3G9Y6
/Foo1q4LX7Jq20y8GXck2BAzwYOd6/e9N8UBBB9WcEMRUsK+jOj83Xy/DUKG7wOHUZiT2r1y5lwW
sT/gHmJWyqyyXUiZ8kPiatJihH1OkJeTSc1nFTabu3jeRGpYrcbXcmT/HiChprvIYJCsVaRslEYD
ssF7hdK2hDVOJyHgostavM1L2Uz/QtCSVRe1Dyjx7vPKXFounP8oUgvJD+OJ6Y1i2WiwLWdZA63+
7PWVLgQ9necV0Sa3jvIJZsiScAygFn2cNk44zFWqkhY7Lq7rA31y8lUlVUsoPJ2T2fqyVHeTyLtB
W/4ebAIEA+SKWk5pi9ZH/8/c2V32zgUproOp1y7wzdqmcHALhrzkMIqrIqkp2cQzL3PDMmD3ndLi
StZXfOH00Mhq3U2b/tCFlzZI/9lHEZIQurtIJeO1BB+0qWWPogZLR2PsrRbMNagSKsa4cuACP5Bl
RHrf7U6IxL50ep2ZHZY+UPjQYgn1I4qCVgCFpq9oRDuHp5VWuGkWNyC9ctsLutsE/McQph0WLS6I
AKkxlPdEAmGrkiinQvUZ1GrnCNhxGboYec2USt6rvVgorlDjsmrE8QocEAkzHx4+30pYyWeZ4n3d
ehXuIt3Zy9cfGiJsT0xuaWydh4lMk7pDoj22o+ayIoPVD2yrNBeHe7vcHpRH6F4WSLQP1x6092iO
7bb8q9G9lx+myfitVk+kL6as5xMw+wZT3BmxjzjHDSc4Yuu3Cn6TAerQUDCZM8RYTrGfEr8adVru
a6i6wUnHW2qFmyv5PTZbg+TFTw3SUn+Cg0j9ke5MAysFyOj1/IYbeQxDmumUthf5xozsTCu/PJJO
Q5i/6qOmKGqCBVQ8bOYmpWkd4twSnaaO9A8f84Dkhu8tLFPjw0tzoBO5qXoF9VfEf76rNddvGuO4
iWygvKmM7MLg5WZOK0PDAppMTkRbgvHW6/U5iEBzhUDSyiWJ4Jvw5iOfaMKyvxlLNN9irLQ7/hpg
gl4ttQ4h6SUdAZJ1A264ensS+uUMXlk2tVoh3dORmiDNL2hkkOWX5N06+R07qoZz4tmFtn0RRs+9
NPnJYPeLvl84nnbYpMxK1FJc3uRmlJx7JasE2eHjcbAVIWF/VM6YX7U8mykDPwA8TSIMFWHnX7FS
PWxB8MtnSqUEbhHpGh6ZYh62OzdxIXodNAuq4rQJoPVqBqd0sVFbTje1/stvXY6GNMFbihoB+pLN
iFCANq3KADeWAddvKoBF1gsU+PUEXvJc8cpyZ5e2nJ4BP792yOBqm1TafQ7qlw9qZMPEBfjjJjEy
WIaczhWwuvnvm0RO4K3oJSWsu9G3wq72nocAS5+GeZZqGGVOZk94XmIadUNsVRNM06sMzzVhvhdI
IvnKdo5+Tutfie/o+MlBOJM4raOWeD5mS8dit6X83vufkcmojGaNYrUQrtBq4kNbU+SqGFLl6AI+
JogOBv2xLs9m2oZdyGGzMC+Nw8eIogX2SpWRBvWtBccj7ZTUGUDb/JaYjmbmaqRPgR/Qv7Io3tuA
S22v8koNJcKHtvSB+H3WFNOarZ7V8PX+FhXd2LqcK2VGQpx8zn4FCl0vK0xkyjT/yQuc9WhN0NYG
FiLfIKBJhYky1cRLofr20PZlXpr9caG08ixz+68jnvfCihOJzlfOMmZulMpUfvaa3mo4K03/oN4s
N5hpQ8I+UmghBlPpim3WH10ki0X/ioFI82QJ1S6QXVuF8Krnh226FDDsSfZ96qTCw0UH9bIsY7Bt
GahBRoFyKz4qAZ+x3KcYgy7dB3UfsHZjfETZsIzbiw+kXB9zAHL/ijXG/zIJKqPaAf1O6IDIsgYR
dTh64UJpviYHcipRyKgutrAwV0OcDxrcnvAXqfuJAb+qIHxLT/H8NT7NUhVLUUjBIX51CyLy1Juj
xkWF3yBQ5nRE+qQnOD6BPN3/SeH68T41WU61bmDbPFb5rysVK6ZQUWHwhP+E25eYt/LAepxoATP8
KI4fSUi8Tnsk+BotT8qUdJNEo0cRAPOpE9Gz8YLROMHMOD2xI4+lW15YQN2hxZPXB2WmukcoZQMm
fSKQWUolVvyxUBEjoKxNZejEUQyyKvUvOwpT6GmQJUd5pEpU6qf36Uu5Pu9ULFI5oDkapccJjP4t
UpXXw8t+l1X57SXQupDuBf/mxH7JAx99WRqw3jEcw9kvDpQw7tEfq4Tm0RKCbBvxotTvPjRxG+rd
++mDPrBszvpvlc+nTB2EG9WXuXYJB9Ztdqvbk2V9U9RezvLFQEZWB1fETSdxo65vkw/GJEpnCGU/
h8tJVXSexOKDD/TWOuBhjUitBrQ4JvfWnOh5261zAQSRjKm0ARu1JKDxoCiMSyd44l1EgyfNe+Do
rpo4e/4EYXQDLzeqaJ+YMdp4NE7k9OrL6iKCd/OKE913CTAFrACVksxRC+qbPGn9Arm4WL95YTk6
xLHBWCkpaHB5uFn8lM4HJ59Yy2YJsMyxONsjDXyd0BUuiDe4Py4ae0FS9PesB/J54rjRcdI+k05y
oiVtALA4q/hAtWEiN7RQCQmrsXbhvISExeoPt5hB3iOluYuruYkWoiaLxWZ3eEdLO1SE7uMzWXVx
gY7FNjO/MALumQYmflKs6ofi4XCNiIRQ02REqj4xTUD52LtJMJnbWYXe9g9FRIC8mJdS3cNjOyEt
6FfubMBctQfD2oWXctOGxWOfQJGrL2LhOjayLp8ApDL99tQJL/wBeBwdFsj0MBr316ys+NFlnwWo
3lndKJG9kmh8sTRtfsY951NwMc1kI3rCfQ8HOizg02yPzuRet9ueA4sIQZsJXTQKhPvhFbxGzMc8
SnDKbPQkWNc+uiZs2rmBkU3cXDu9wuHUXw5t7JLKT9mc3h3aotHwQb4eUa5OB082B35I3IdjJkij
YaZSSoOl4UAbINAzcKn5MBm7S6DvvvXK+OXFohEL8SFAbY7sLUWXlfnBBc4yLL8lFHrGGhHzUsCY
a2xABiXgnNYezqyIxT0PWQzHJqlGhvfiwSKQiFWmzoN6f6tb4gpsqxV0e2UJigUtjSBXp4GzOVio
X40RHhxJhz03+S85k2BXt8Hv58z2Mk7g/nUqdBMmP6rSRSm8uDcw2IpSMEb0OcdyR9LiMTZQWwL2
Soetlf+IYE+GjiwUPw1beIGVDbYSgN6as53C73RDpb8oCOC8fgrSAbH9wTiRLKqmdfB9Y+GckgxT
N4jY1Ae7zHztfKYKehX6KIKYDA5qHndIq8P4QUcGh9wRg3aA3g/28b5+rJxxt2UX+5cJy/sWbrty
DkyrBfYbVo6J3FX7uPJrDHmy4CkiES3jc+DhzYj45FtbElATwOb8YNBNXmWJGW6PsFsCU210Tq+e
QtRseUUXxCc2iLCyt+xbTtIDpbEEGmRt0fu2YTJrGyCVGypg133TeoRm8WIB8x+FU1HPBzh23kpB
F+JrnRhYkUyH7R4pda3QcAvIODNr7YnUz/y/xR4JEtM9bJ5Kl5rcMfmMLYHzmXwXLDl3m70hYlrJ
zGO3Z/XL0m3+LSd7Yvx+3YZv1mg1e3WviNxUDVXQor2bUX+N5zFxB9iZ55I1I+HwYjUKnwA13B72
Oj7BQT/daNIASydHtrrKlSr5ejVx28unb2Eu3YyD2UAlky6+irDZlKKQK+zkOlPO/iapuU4vvPHP
WnIYy3SctEfwjSdVev7RVqh3p2hT3o7spgenUy+2AuYH9covt0oBG6JAjpYqG2pxowRy2gJuZToX
QS77vxpN1xUoxwWRTaooyQ/i4MGpSUsDjr/FfuiFDiFCE3ZK975a6nXCD3eq6mhl4xcC+4HIwbOt
EoK03HMDSXSQeRE4VoyqsHkcGXsdpcWrK51kdzWjSGCrfuB7hM/TedaMm268oMzbq7/IW7u3z0eS
X9iGFIoFQ5Ohe4nefwDQhCtGpXStwUoaa1AoPcgFCTBCNWqWr4ARhDwQx2qw4LUImQVpqmOrK9PS
C9xRzIFDk0tQF4uEHZUVdvVKj3BikLYUoR6DXcuKaqwaDD3uL3WnjYTRVBDZ0lAK8wrqkeOMC5/6
Qbnj1+XjhHz4aoEFNsaiVfpfokYb9ZMFLUCbG3EKmhTwH+CXHZ+MAGE8mU8zwoaRZ0K3BtfFyWC/
NoE6vs2/6wGMjHiXOuyKZ8/mvMi8ZLo8BSOHr4qUBIVX5qh8LG1BZcnVpYf/DqCwBiABsDDE37O7
L+l4ax6Ptsbh/pQndcpnH7q+yJnTnFeEVjCmU9P1WRlH6cQM0sY59d4SkZNE+FBZrYRCwnFIYTkn
76RNv2/krfQhPlO+/1LQyk+AjC0bRccKmszZAS9kPq4EQv4NWITaIYUACmbZIG4CkwR5YmG+xj+e
ugRmVe22F752Q6WUr5h8pg2GRvrOEQCb0iYjJTSZ/7mm7gp1FXJ/EHiWr9miz1ORrnwh2a+75KLW
RbB5fhzCND5kKB7Zxge6xgZbPnN6kC/k5/5cJP39pDD/MLwgdDQsIwx10uQDbzAVkp/tFJLMreWs
sum/+4Awbrruuz4SDcs+6Ez9Tsf/IRpl/Ej+N18imcncAgjwxFkqSI+aCnY6pXJgbpn/YQiWEm5U
RdEe8OC2H8OC+BrKoS+ChUN5gyIsJlCZSH9r+RqYjOOVjIpN7h+RqB4vITE+in6naiwwEqlzdFfZ
DiUeeHYDpbv2Jis4U91XsitiJKb+rZsS9kfMjzt7+dnVoZ1ARK4JCYGJTT9lzn9ApvZIU3LUs/Y9
TSeHSpyfZMmJnSRJV0wBktyLCyZ8wVabzBscvZr38IwK/EgH7dCJ+9JuIF8Au/jmt4Z12yKVrfY4
hJStOsFlIe6q2r4GggF4jvyjToJteKFFZb6xcigBT7JI+klbUHGlNYH46yT2wXFxVKeQkTLz2NG4
ELYQ0OncGD/61msEvK1rzIpdI31+23qNEpSOpMX55ljNh0SicwmXAQ30N3x4uV50UnFyx2FcODPD
VgSOF2gDI2KQiONvFsGSW/1LYeK7JhdSeQPVjD6rMBP+eurFrJ7aevzTFsL/tEUl07VrU/RLxpIQ
zKOxulxWxgbBlVTE4ejPfmC7p6819yO17h3mNU9JznIrBVpBcAR3gayAn9o4RV+KgwG/DhtpBVD6
RHarsIj7TOyI9Dg0mejiYD7CH3TJ85ApaxEUNZYQ2XaaE7u/HKFFpPo/akPASl3HNkILlp6SAi1l
AL3kFkwSJP55C9fHkViHrNkZFDqJP71DfVjReurg6GsUzY5TYna+UC/EIUBJu09ZuD7qqkCmGz9y
up6EdIVZYElCAlIxhdeFi8pxj6HQ+/Frj59z6KWW3eW/umfewCCNekX82kT2FcPQtMCizf1bVzFJ
qQAvcdjOpWJ6thE0Aec5zs2n64I2K2mA15wtUPnVyvSZXl5riEhurpVNYTc5zIPrERZLcpT8KppB
gVrdQAQ8vbbQoMHB+IvNwfd4F4SbgkmSu3TiThY6c5z6E2x6lF+TikR+Y0Mv5dTF8ZICmW7A+HOe
MNKZQJeg54FWwQEPMkywfF/+Zhofa6RNRcy7PE2qYvOhbniomV831oaDe2sVSVqOqWsbHeuz4oK1
q1xjtQAcoCyYHx2+ZWwULhcR++q7G/EJvv9ByCgpmhQWFI36BVeb2+SYKAXkx/5qOXev1Kt6+4sK
o4fPUCzz+vbq1umrVUK8zp6wYwLuHO4GfPEVHBa42eKybTPWRaxHB8tN/8Nxp3ahpJ4Q6g4EJVUt
3M5L/KIEWXSDVkBXkFPyQOt2qvxc3xHxgZ8xQrYNS0KueF5pISwSsZpsfFyNZX2CoazR8JPRHrQf
U8wy5pguQVr5rrxdTos4wp1/LPv7psjBjSe7wz4r6jtJLCaoLgmgju7pc4Z4CdQcDdoyUo6PIBKQ
CmclO4/nps9djZqDRY2G/vVEwe5AyhFFm56oOjIPW6Ad6KmMOH1Tkh31r5wcq+KdUsA2iPlOHrCU
0Bb9nO5F2LcHeqBvabMRIdsW2UPoRk8YW+yADKLCuaV2nYak8Mp+ar/KDUIGTrCP5OEYKAEkVkA9
zJJl/lBv3Eu79ss6foyurq7WYrQByhpI2P3EwNJ4C1crlW/3RzplGEwM386RtJfymF0tYZzv5K6e
Vrwn1kPNUbsu4/w3u0uIgF42t/ZOUd7FT5sJi/hlxJwSvhKTGS+1Gcv4ZIOjOj2nNPLNlAdhlMQT
piDK+fX++3P5wp7xPERz2MeHi8WiMyr24v65Y8THPhsEKGqGadmkTPRkmjd57vb3zweEcS/ZFXUe
j5VOfCG0uI7FHk6FtMbRHnKTGNqmkYFMUQLRFeuFhZYt3cRD7jzuQaCJVBnGxN3EQBzetZSpxV5x
GJ9Wkyyt9RJZjIJAeFpnJgZsFMI/SQCAjks/IwEUImboL3U2aKFcZnSp6/wpn1pokPFBkC70SL6t
3N50aSQDqF5r+0pewEQEjXjF9D+q51jvfYiSWPDuNDq9juWKTqwWtPggdEkYGubskBKf8dPwoajU
7w9RhX0gkj7qfDqKq8sfr89IAkhEnPoehPPGuHBhTzzgv0cXr27TWifRVVZLv8jl6Q3cOwSfEb6m
Ra9vWOZQVLlySOU1ZHVM3rXMEa7cq0X4oRm76vVy5hnUMmahvwwsT2m3VGjcOJKGNMgsxqg1HlDZ
RoC8RodmE3DtjQk9fsm2o3AtLJJa08cYvrnXeOgZQTi79khVJOl4U9bbB8Xxj8cjligEkjAg8DNk
k6UPPs6y2YwVf27YakLoJCwvZ15knIjJ71QjuMnritWh1pxlhMQHriiHdxP3T5Y9FNImBcEwdGsJ
Tg+pmjwmTtYek/aL4jeTfNphv0AYV7IoVR3+EWK8aO0zZdSfOy+Nmu10hudChJt+y0aYWWNiG0Pa
mW+yaTFYdZD7LH+M8OjlzHoUA/FwVZUyZuRxyNcsUZbZo9h0i5j2x0Pfg5BtS0Vh0HrWL7Bj0nYC
nvq+823jCXIVNQnQZRFfNppqawxPEZdX6Cq1N9PzwYbxzdVLOMf13jNbe/P+9TjwN1qHJ2dABddx
1vf1OBn4mShEGFxjIbZ4t57owYG1GYdM59n3INgwToqoLwp25YknBuAQ8f7ZFCLkikbAhKqX4qYQ
gfGg8wXSlP34VFW6TzxD+OVLei6ritumx6kjEuKwMAdErDeYVKG7sAIMrQ74p2WU7zcP6lZh9wow
IZvu2TivQdffa09eUekaDckR6zTUpw0oKSSY1eCd+WhUCk+mAF2PoSLkC4W4Ojo5GO/s4E598dVl
4uTAKBsDvMJzQ0gZVv15SaodYG7EzILtjKD1wg0Xvsii4gKc5HdY3vZMTrmBscJqBdXzb0QtMVrn
2e0TKaVjRKH7xEBTQml1vDEd/TLJaLWNoVQ44to8b9rVJbp8EqU7oV1bFBjGYs6f3Cwz2uiXJhDw
zZXLjLB6Os/TGeqUdL7YJpu6oetEsLRHgbFVVrB6d93bxGBbyxN4w9Xs382LaXUgXLnu5q2l92HE
xal5TTDAHeYmqkLiRJEATJjqllLr5/m0/+NiLIWrK0X6xzki2z57NRgs0GMpWCSHysROgaZM4WLg
T0ncKNJYYofkdtAsVlBuDf9o3qC7YYf6gK++61V24I4eWWn9WUkbpus26bcEQJUN2rqGVtWDLZCc
EpZaqjFo969cKU8VTA3LoLF0/gx4sfLTOcraIpZ6VvyyA4e1aNcvCHdShzPl7jferZkWo4qNVYPl
rHE8ZzVPPKDO/p4iPhcXyIrY136ycVX+nk5iaLc8Xqul/Jv9008XYbBS85c6sC6EIC9PCwIcbAH3
vhvy1ybLs91Y4FfQtIs57XFhy+0diY4VmCfgT94yoi1SayPS4vzUWjnalmxmogCUfAygp705M16b
Hu1QC2QNr6+eT/09G4CEkpTNWzYkb7qs3+62z6Gmx4UHv8VbIZZ71YnSqygduVULofRDysDgOOYV
ElD/2gsqX8ZjahgF4VN54eR07B5J7xjoZge0V09HC1Ta3/ZTVYTqFCwX7oul19Uh5skbl1A7oNQK
SFep4GCIGI9ZZXnGK8B44oBW6dE3ShaTlaNz0vLsmnkculbCkqVEQxGvrx3H9Yd68xFur8NUv/Cs
7IBRpqTghK/r2RKk7aSkQSYhkZFMY245iFDnk+0/XbUDF9RKXeuxvmAvHQu8jbYt8arDVKLpwknz
+SInFVEBLxGOw55EdQ5hTsMPBTn9RzvbI1Kg2gsQZMVtAxmTEX2t3C3OxYUCDPbcm0Ei4ojlvXQJ
l4DObPK9SvYn8JhXeUlTVMMjwWZM47LIdksFg/es73qMrKRw2pB8962tDBrxE2Vz5lGWHg6lXGTh
hk13/OAnBeOtnOWsuU9LAI4WRedq9eh6FO1371OqBhx4HL7dCyLnRLF4L0+wjYTKCLeXcQ/S8+67
b5fyLiGD6mi5VNmUyaOPfQcDtu18wkMVQd6GagcEPiDH/R7eUBwAKjGDWSuaxIbA1+i1HC4T1Nrr
RDV04xuKJKf+Qda+pnQxLydBapQ1B6+KVT/CFenIvzF1fKfKT+HA+LzvXH1AoqLcq9gAIyFNbjV5
wMaQSepjvQs77iZD65vCKWXR6tLVEIGLhlx1HczyyYEZvkr3GSuV4hrc1BfMR5x0ulXfwSQFZr16
wXFqH56TmI3wc9keZP7o7rpc201GwMgA2QVRTv/IKYg8tzfvfEOewK2cHWlQ8QgabgB1DNkKUkNz
oqgGs3bfkXeJbgsTwWfDaaYR0kUQWRBm5d/pppPT3SOmTaCPQwUNpqMfdymhB12IYjChCKys66eQ
q/IwsuEFt2rI63GUft0wQQphZ3x4l2tTwusIx7ZnQnKdGHE698RVLayZ8AX+quzqRGTV9kj0WNVg
bcIYl91EBLM1fjg4+ohWpwSzxJNwBriN7kYxtm9bR19NLw+ZW+u58lWbLgb5TrFi5E9MqaaHjF5I
/0pe1vkM2zv4O1gsm4lvARNGXDlrVPUlwcvwzABfl/zfa8zg4OIC8xYgALZTpqlAIDkK05QbwQfg
Hen1NKg+bM1djL/AOXOpdjEvReJffbxLEoCc1I1QhUjpV1eA6sL3dLmMrQ5TjS0X7OTjmwZl7v8W
oWd4/JzEc28F7AMwiJvPpGjiR91l2dkHTaVop4XrXElgIg5uni/lswiXqD5kMKmQTwgtPNumZg8T
WVQzgwnv8QXfa0D7kmT9RSFxyQEif4+hbuNW/WUTEh1Kk2HB+VYsfWooQQ1+c1TLuXe+LdP2OJlz
6G8wbWT9SZD+T5V+dMz3E82KhW+a7gZBvivKBWsiVIUECc+aNUA476cQlcyMC1FBqVf9cMHZMq0D
YKcmhmOY7Vs6qrC71NHavvHXSysCN8n2BBDYWCtcu6EJJUYvpBBrSWVVzcs2W0wOYtObcmAlDtz1
JsHijWnUPLeY/RY7vHzUOZSyi0SLQch4rzzn231UtLhRNuh/clba6286U6I/BogDma0+Q79cxNOf
t/toDRQhQMltvZYUz8+37t5oBqq+C48Cc4CMOy7E17lH8sb6kUOZtKANx9Z+LOjdPrIcsVzVLOfT
V/QkEA4gOnZbyPGT2nKhYlXJod0UnUUm3YZidbQnyyGpiMvnpwWiKaClmPDH7KF7Lo4IF83pFAq1
Yh1uUDsBGsBNSMjvExP0XHRb6J7g/6x1+b360O7VMClklOy11syVl5l/4EQrdVMa4MpUiYeVTgYI
5Eq1drkTMRGbluYcM9Ix/8G62LYhPTsU/xLPpWgbmER36aIazDpVzBkzgcnG0AizPP+UOUVlO5Pd
4C7LUBDGgf6mOcdB6Fo1okxiAIjkVFAbFIflf4eWOWA0Qr6d18pUyTIX/qKwyVtTDUMW4Elkxhh2
Ok7mz+JstAcVkQ/qMtGP8AQ/OJhzG7jsI4x3DP4R/TUpgLqapvTZsOs47kjFvIKl7M2fVtfodXy9
W/xd1hL3Y9J8vnAk/JjKan+FVGGuoxGpdUpzjVl9QB6uNfM3fcMyuKoj3OuhwzEqSp5F/Zizk6gv
XXE35dWljgVwQTjZWeTgabYSEWnNuo1HuDjMYMbR5tG5GVquUdP8myRoEVS5KCkLshBW92lgeC43
Cw/dTWUsGnjVkXG8oo+RgikOjqeClaS8S8uUvPt/STHzqMiryP4lns+Iw5c/cvEXJqUnvALYed81
THLxxVblTCeDkxZ8epqmVo/rO4yOHgqpPmKEIEzO/O+qk+e1s+Sc9AUt2Nk/u7FvMY9yuTMw7vBy
ADic5FfHVMjY1YGVSbDKiwcp/cjcdJvaWx3rkEQTxyr4gCSHapvGS6GWhxbbLhR6KVDzWrc7NMcE
YOl5CPJnOfAJnHJfro5Igc+pIoOhleFsBXvZEAekC4icfD31PHxJYXg5G2EiCYD6T5QLqnJkUYCS
f3SXCnYHravV7C2ChHhdmEHqxkwcFYXrzoP3VxBGnvqLnsk+C2D+Kmk5ok/pdjtbRfJgsxr6ViqP
dHB/rJKTtct7bcrqFSyj7IOiV9TmuuiyhNUjqy5b34THX46acYUE5IElHtg19fNfsE4cNN8m64XM
YlECLfCrChr5zBgJoi1qiOLIa34yGpZfEFTKGuXxCsgnTTTa9U81gcv8syn9xcKzGjoQEx55jm+m
hu1BdvUJc0+bDfbMDzXLphFHGzfMN2caXdOFRI5Kjqrq+tgGNFWlJ7nBQfA4iUH2hhxduoGZ5BP7
KF+Etb9XK8PTakjPuaq5kUDA5+8pbK94Mbfeu4pi+mzrb+u+O1tBT06O6Z0S8Cwg4cn3+O+ANT3U
XYVh0q5FnVLNQxz4cv4U5HpYZ8N9/E7Qvilhm4sOLz/3Yex2AIyePZjIRROUP+b68PlmsFrrhZFw
rG5bWp182/wP8bHkSWzhiUAbIbe+dnSdrxVm58jlyaEqNOmgjQgcmBjxO++JBqnWtoWVqm9vSiZw
WsGkO6MVpxByliGR1FLWXAfMShTEsqkZ7MudxCWI/htUSGP11YSOfji6AQuCENpC2ir6YMECInCg
7hsk7w7rC68mTuabvOkx6+zoFFcmlqlFKmO2kCuJ67J3Pk90GA7vyElMw1ZAfqAvjmMRIgAxGG8S
XVP7L1VUj5fCzk1eGer17ofIwAlyKICMISrXpoUmh6V9cicn/tkyaWOKHnE2OBfCIXpt/XbdDpDM
QIJ+zYVxBMvnc/fb0TYzcEnrV8xCK13VCgxI3oZ+gNA4S6vGAVa2cbkkRPYwJdQyDpQTolY9AnqP
htF+Cf4yXT0Sx2dRpQFCRchdwZcc9Lgffl2dVL0rFsi7+XMcD+OLcq1AtaL1MGqGQ2UASVvJqDcn
FTlrjEMNKzHDTi94BrSVgDEYPAowuHA0xUDBCPklt4tw4M3mkG8iWMZd1QuDPr/qmvGkahDrzawP
Bos77ZZk8UcvHhjDjJbeg2Ad29Xl3TKtw/MneeiT5mzb2eulXv0kZcOyE28xq1Cn/bafez7j35ma
GDjfnoeTyMM+pvxhcQ7OTQ8LHteYpzWBArzIenqYJbjJ5ohhTp9vvomwkIFhBVlWR1F4khgC8p9D
nt7VRKZqVODd7LWnoR5da4vfIUkqToag7nxBEWA1jcNRJ+pEbm9AGvbm6Izw4K7QYkqZtIphzhxt
nyV4kjxkSqIaYqlxnPHlasj7umt0a/9dPXgcnoHot96Ij2LjoSy5rTAFudWxnIKBeJqm7nk29h4x
Frdk4HvTdg5OkxZYcYaUPNzbJJUdMrzeedPa8ZTBNZkgw9MDI3i81oAia4Dn1QIMbr0QZr29lRvK
AL3awLqfNVRAotJ33qSgLhr6St012sMequuUS2k6ApHmBBmizpWKc90wxNRlnJyp+52ku7ZdS4MV
4jfaxDIRpn8/M3CVn50ILSO53FKEcX5Ct9pglSniFu3/Rde/VRUeH8k2GGh+RrRCrl49IecB3Kgu
VejCDOltEAYSuM5TmJX0f55LQtqTfKuQlSEl/9n0l9VWLmEQiRSKi8Pq5eebAAjprtL4eQhp2y3a
7F/y34NqwXE5ltyIaS0zPUgA7rPoouDjKBl4hwJAzEj0nMW6I2pLYd8UbekLnSZW3QOvQQD2k+6M
sGc/ue/NOBWlE5bFq5eZLUQZbrUi7W2RNcarYKpgAr3wPFwBZIzwEZSrUBRC2CChC+SqBcDM71av
Prz0xW7pRFKpe0ubMl+x9taNJ95HVAEOkCfYtJZqoK3MVYc3IMeIQS98kc8JSDuwElCuw5xvMT34
GkHgB3yZVdLYi0JQGlLnB1fgrGR5IZgwFpntzmU1i9Z92TpVpXSe2ayDjbSAbx5LxDqlSoveOlEo
M4zfsTs28+wvRBNCJA1jUhDfJz/KFtsk8cbrvV1MYwWdNpuVIJcxsO3uPTBHE0kJbzg1af9hZmGK
whD/tYQIZWISHN6XtNoCqT2KMxc5HrGLVWKNt2lVry6KyskNNrKkhxstl+tUJ7KenS7kdflPguuQ
/oFJlrNnxfoBsDsV9TXJpy7OQzjok0dGjW7fiz53DMnAJpsDiCptQEcvSwadx8Xr15AdoCGG+X5J
eOcsLbuVws+m4+sTzkPw4fUSl5NLbgP8ErwwvXiXm3+nTtT03A9ELcZLagm83yREDQ4ZbTJ+eN6M
vhqtgBmk/hsLHK7TUbXVPb3JLw6HF42HTJX3kWwZKFLsh/SYXgIa+PVzErdHgnIgTtBft47gw3wX
uNEulkDeuCzmfIRKJw7FM07yO9WqeLHLrYfy+SQ+Cg3Ka42+Es1+2unaooatakxtIf8EBjxAqal3
gMGT58tjwZaqH8JSIk9AikgR/ZsoDgY/QNtlEq7taqc8Rhdp5cZqmp/NW1L0JD2JHbXxfmZBKjJ2
QQblPuO+RFPkG9aBZAspKvsxYJz6WIe1Lf3gx86WfKpoXKR2RMDwj/TuLs2ZlTabhSaIHpnqvqBn
ZCAGdEtcXpTKkWF4gP0DK4F2diVJiBYA8Wco2qsq5VCRywDNZhbjB02gYcgDufyjT8mfGrCUxhQ7
zih8QC3Gn9tr5S2ZDl4Ta0rPD40ypnpqR6TTj71y9u9+mX4zfphxR/IEGx2k6jEff7RJlQwwKd0/
qhpXOg3vysI+GOHxr2C909j5lWAY9DeGiiebSc5FSEbtHwuJUvnfe/RNuRgkuA4IccGJMtpCBWEz
JNPgw50/EJyLr0MZwc0pV5gj/HN0O/KIAim+n1jqAQrwTTYhRFNsmthZoH0J1QKMl5V2gnN+tTYb
4f4O12jt9mTMUv9+ApRSx3c2h/cXLfK2ZSAGNh6vfPJ/wxgd2ilxdsr4Jk/EFT5cOh1CBt0e6kh8
tPxsFd61eO/KgzXz243WmseJLz37iQXVfBk0keLXyrc5fSK4pdpXJqkp3tuY1yuS16GBpHkMC+Ca
3/SE4ITOdfkvROI+Eq0EzfYUF0/j/XtvTJE5NFgaQiUkJNG+3ECNtLGbGYUH8rMdwpSzQCX2BHcj
xuT4b+W8SV0tu8JCRxZjvbDi0h8gJsOqyZAGMfn+wBIdK2bzOjV5txGGpTXt4AgV/AwmVKdfwIW2
nQYVjqW6qbzDyv0ASgbqJC8DinuzN/Gb7s6w9yUGA9V63vFhtQ512nkQRCQRq1yBdewV/hDpHAjR
zvadFfuuxZQMWjcECQ7dCwmsBgiEEAv1bmJj4k3V0LTLqS6vIxUkVBmtzyqEje4TRdF+LUuBV1dd
j1iPQhOnC5TmkOLNn6KvGsh3xSwSa3gRo+Sq/INbdszWcjwHdKu3JNo8WOs9yM8CcNtksU+y2y9P
Knxbs9WM+7WC8pDbDbzrghAAzdO2btVuJ82x0IbFKMpssHzx/qx2Syzj6YndJsiQbigybdiKEg+Y
kmFetbkl6+axa09XDGz6nGV1a3ICWm8aeRIWvSHQkW43jqAU5DO1D87gsi78jp5VHiCwWNqW5bcy
sv6dsVTVniG1vYIcH+K0tpgVqqom5sqK56ZhwhUlIiURdfw2YXMOKdc+5PssaTMJUZV8kcuM+72O
CdCMUSh/KmDPzRAfFNHWL5EdftiaOAiuGO8Y26f4qormWl2MHOsoJ/YJzqqTJZ2AUDR/5XSwE8TV
SmDnDFHO6pDadSqa2Z5GPvqdn0W+4bagyJXHyyQWt8yIwKEO2R5ns7Y4ya3SU7m65hGNCrhHdhHI
BKGWcMz3Qi1ZmOHffwtNHFd67+J+6ntbq0ix8X2WSrriRx5UfiiTolEzPyxwnq3BQZjOxPCViiMe
Fd7YQ0no5g4xX5R4eUNdH3oTgr2R5zKLVhaAH6ll0CrJO5DsxvYo7lxxx0Y3LplZdHoyzll6uvkg
CdHPQ0zlAXxfEGhiDQKDcpp1H35vHu0RuNZLj/a3lhU7gPklw1dsi8sprs4fMmABgQFOrwaqwmtI
Lw/txHhE+qexftfqHGyjc1svm7zCO8UVpyE5SglE9Iz1nk63DvKg7xtwAWlyOtjOeOGxSiru55bl
ZAfJfe9sOXhGJQZOY9oKDiWQ08L6Kr0gCVa2eJq3c8+C4LWC7mS3QrNE2Dzlpp5aDz3CD5Is6DgK
0GXaibyUTzMoSCiFQ8yectiteljxB+zrQ1P0hsPvMP3VHuhFuhxSTLKSskwTPWr5nHy97zXSW3jW
WCK3kN8puKu8ll/F05UkNlF3XbgvZd/Vnm39FoFdyPk+eQDC3BVLgaE8tmWxSwnTmyhDdRxQt2iv
UywiM7TIAO51iJQBeFVh3T+AhjxbMHRLmwbnkaqFufGpsr7TtlSB9UnlL5HS490HXb15zrH6BggU
YagdOIGzUzPOR2rFeZk3p+ElJOgyfiyiEl2YxuZLQRalitC1PhJKw5xKPk3QrGDRD6frQDDMwWR+
QJUdDHBqy5DXn3rZiCUPOctMRMz1Y7j5xomG8RTwEdrQYgHEtFKSRmXtVQHJ9eMCR8x22nvnLck/
XT522EtdhKQBrFZt5SS0tTmHxKpFCBHlqO7yttvbZPrlL6gom75cYijFfmdmoOO6V/KMWS31kCuv
KkUWMWpeIr3a6WuqZkSA6Ru8e039MJEDqED8W/dcDmBVk5ukNLAXRY6dO8FUKUzNasi77ilSOlQR
e+qqPTk4t6+LrCMn8hhsFpp6kiHdXpjmN53oEBKIcnIcaObabIGrdkkT4/YPHBsL7yEezGckChjp
QU57ngd4uBafj1Q1pLFr8nDBl9P6cqF72Ty4aTeCWulR2p4k6yYJePVBWcYae7snjxQnbl2CJAsb
QNkKRqX4NvdfY35kBaEyXKH/TR6MfhMfXg0SX1JCjSZ/WL/NRpGyrfcRr+u+T41n8iEOggs3zxL9
2rpuWcWwoD/FfzKBT5FLkNlKeAVdFUa19CQrXb4Vudklav4RrPAclVEHMOWsxmviyFt/PA38VKZB
Dv+2gUCQ2hNQhyJmvXBHS0UGSYLC2ACCd/b0xtvINLZJSaVFbqy1+BsRPcyxDbb4SE4Y8Tqprklg
Y7pBNGry6iTL2GcT3jE5QM9ukh4PZvPll4oB18rqWkX2XAI4h/k6vwU+GPU2B7AOfswPpjXtphQV
EWTzJUA47S/Ne8AHp5r4lp7W/2O+KHn757BiII0OvuAzHERguawIMI3SfPheT2MElMmmtIVzCY86
+PKc499LI+fb+bRxWJC2X9SR2++0aAsvR2Hld6fiExq47II9Xtemck9s0zgyL9aOf7oDa0dRcS84
cZKpaLZeF4pnzgYC5Y6qK/VFy1CdbvksCDEt3MWdztJOy1xbq9rvF3CWJa3SaigIp/rsZivokcbI
wB8SfCJFboSUHVyKea7fXRBEFnvQq7DmJ310/uw0tSaZGovlGbaLE/obaoDReQwHQ7zInwU0pVUh
VzRvT7+ROs9tMJr9f0KOlijEan1pYLPG7YQz01SDKE1O5KHLtndhG317wjQ/9MKs5vX/g0Vqza0T
jlANEgziNTkkmSaLFRWep0EyHROiNRNqsohKJZCSbkAfMYhce8IQEWGqJiifHJTcJGIvPzvHD+2w
HHgsnlbFTJzUU8sxU5hQKKycBUmzJRp6Qe45D11MUrI7H9nqe1pdlpaPIQRGQtMiDZBYNY1jV3/E
A3KOT4Fw+ZKdrjWL0NdzaDyDfZ9zL9tlO0MRjoh+YR2EgIv66Lo02KlmH3aVwhE6zHfQlD47bWgh
DC5GHZ6YPnrZlgPJt8/TIAQ4J4AovdG4OpisMRq7O0BIZCjzRCjd614OmDLYOHR7Wg6C1usa9bHv
tIrGLM0W/uhhItZ+OU8uGf00vb70aTWOzfsbnSzAQt2qWsWSrFK1smHn9X/bKXf20lvpanaq0gM8
r0MzYAIWw6Na+F69oBFBiHChbb21jVaSFOJSWW090LjA+qGMzIObbPJHLN5adzYJJXkOrCA0ABZ5
4ssQIel/2KVYJF9NjQBEgGy0+rRPfK2UQLRvW9v3ddhjAI7lbkOHdt3LZQO+IL86s8ZIP6amnBkF
wH6ov05VbOjL2DVh+wSliDE8M27R/CmvYccraDsIwF9xYTACx3LEELyVSASn/kHpLcWTcYesfT27
jlCVTu3+mmAx1GM626pkvuTdG0RCwS6vIZPU+xvCP0NevtKU60fVoUN8fh6jbGXugwUJZ0BzAf8o
esm9QJlvTcQGOfviNUl6yzFAjp3eeBWJ8mbL5fycGfapyA4KyaICQc0AW82s8maCoRkdMKadj4EK
hTGOq1VmfxyRII+k//KhssuAIjoQfE87NnqvYUUy2fuizcMuhrYllrateewIgEdPt0L/h8l4erCd
qyYd3jgBsAdoVd9pM85v+gNcj32wVNkWnSuDIbolvq4rJZ5drtF4f+8jZecfLE1NAX+zJIEIcXel
Z8OX+3g61uZ+D2RrdalStmI3dPWTDvs3kl+z8HPU2ows2DCwzy7Vkwk84FRkdlK4QLQRckYZe7Ve
aoFsKt5tjzLkU03BxokiVUuLgD6MR8mEIYxsQBouD2TNWuTHvEPQ9EDF3w7J5O0cOs+aY31ljgnD
oYAwcfns+Bx9AwiZ8EBEIvFeWxq3aYaNP6YOhnVtF/p9QaPwrb+r+24ppD09SS11J+phcM/w0is9
76sJ0nMxwy4buykbIDcsQqhYcFbS0PYp3YVA5Kb4zJuY9bCNvA+hrk3Ex92++F+xzJ5DYyaGnqfB
b/N8L7H1YePIruUOOw3tO1g8+GsEcz4BQUePRNs8BaWMQJhjiZzTrBrCjZpbw+eW7eKOUmBGyVKV
gZozldObZuJMIbEUQ0Kx0TM66P1Yh1xvR6YHlCiXmGVYtK9R9WhzCtwtyt8kNSfv6s4VTsm67d89
GK6zsNFmg28cEQwTOfDndiVIfVd8QNEcB/dVlKHFGdl4zzfEbpL0r1l37JZs2Mh6PW1mbgtT3cQB
mmVaDLiCCtOTBK3mCC2QAjL79pJibFTS3JScUB/tazGhGSvCGlUD5Qsh8qo+7KeNpDyHI67NVI86
fG4xeTtqI7gXj+XyA8BNGOpByVemc4yUbnMJE4y0Aa4G+h2yOQpBOUJnGNHevmBOMmhvv4ui7kBd
Txs5eMSQ876HEJpD1UBj7giOY/vdttFCEP2k1qe3I+8WxbKQSWOHARhcSnapF+UgJ2piD2guk3gJ
tS9XKpG88FD50heiEGqArN06u/t3YMxRweFNDUpAtgMw8v7zfjt8Xu1lJtoyVRifWvs+S0j+WDTU
M/ILnw5uDgwP/vQOAFVgOtHYWi9817qqnaV1/TAsFDtbeOJ/be+VsR8NPGeIjNOvOgNU7QhNkXtE
7CtiBWwuq4stN9LZ9WMfvgi/6xkm72yY1I86ZLjUdg57fAvz7MlEXBNXiP9EY3CCMgNBs0oasLIX
R7mgkb9Ybg4c4MjC9xBimLDIIOm9xR80t6sE5ENcl+Mc6Wj5M61odwzn3wErtlb6vSlwgKUldqtw
fUOxg9OlSAqEroYznWrW07lW3OFRaNWFrnobecHSAaCBzaAv3+OKrhu80a3RFl6/F1xI/3WFYNNu
AT4aYHhH8J4k63yq0MEE9Dipsc615DJOwDYG4A++nWQXrTkaTJB4MWBbPPfcbBM9Y8/0aARQOndW
kXcmijZlJaxFiCMJRxKcHREPEKcRZ2xbbnoxKguvOzJFE4QuHu4mN3LR5WHiYUO7yPiWv7gg1EKJ
E+mS3k8H7Wt0aLOMuqhiPshlBTayaTQaw4TPG4goWhjBqfyH+kIguRCm9C/+nSXU8qdQ9j/IDboG
ibJzepO7J6r6CvJv5ywg3/pvbE4Xb9DZrNZM534ue/54iCM2g0QiIDXpWrURG38bqLQkx81NXO4i
NiRbKy2Z9lOQqglrnNl2gogJoCG0UL3TLZM3S9fb5rmVARpLaGrnIVBlqgUZbjHGWkyVE3HnOljv
bhB7LTJTNJbfJmfes4gPj/M7pEAQ8bQA9xWFkjCcxACd1FE93y5PiZULzC4Ek4imR/AVvEv+2OFP
ObN/jvPJveiEfCiuE53DHtcuSOuJhItJQzojvoNBPkvDHuk4SPoSne17aWUCqT7dorol919m5f14
HAx6Ky7YciosNPt/NBxTskGabDTwu2bnr3sQBYlEvS7INa2dovpwj78KlObIJXB/9RtpWCdPMk5w
ZNQmYgUFLccU35iPlKTGLz9jz8sQpbPtKthAusza5Y+HCViYC6LVQ+aoun3S7M1+ZapuvADVKvQx
3zlEG2YGg98I34Bvb7DW8ZwuJBgZ6NfBg/M+5SZALfliT0EwIW3+god8mKt8wI2gxCf3xEfydzDz
x8I9gAkS60n+/gghqvDPyZXdSWiqPdhRUeNlmscLp4E2CTEUmNyOERiePRcqW8KjotpVqtbgsDz9
3QjPrPwYS1wYdVsSzXbb08qT2u/pPxjsX9MhhPC2wOdmkWolRguJS1Yb6UmD1IcBfGkSN9Os63K1
5XzaVqgLlbfru3Q4efHeGyxfqnirvSMT7fiqH5aHI59gge1UVdouMugJ7I+D/1JpG3ud46ZRmZlx
MrX3ZHkEtQ6qdgCB1uGDbpeOKnBlYqeMHkECRZAB2TLc6yfDN1FQmQyKL+lCZzPBcM1wDnT3n4vi
YZzJVEzEe4+uJ5/fPBQOXzv+UGm6DGrNgiRSrEVHxlrIL1ePhONSIPz3ynL2mJQzAoXe6lb1Sn7u
UnZdF7SDL8JCYU6ZtBF8hE1O8GRxz5zk/lHhWSxfKDJY668unXJ4EDdcVuoqcx4LsFb0iEmWSBR3
oRNtIsd6RBZ/iwUyZCuSxHOI3zKfnxlIwThOVh/K6P6xLf1rXsDsOFk4EYrhd7oQyKkRHBvoN0X+
BSzK8IETRUvISOE0aGgxMWrCcn3yS2ZATmraqHqPQZPbrmcHFdvZQ4tWq2t1HwryKrG7S2N1kSSK
XmRkE4FReRd14idOlAixJLFu0Qvz56rIYMHF+fpQH5wABSa/yPzYhpk7bsItlgCq2dXiDBoQ9QHm
ezdQK5yxZomgEOLcUpc0vcuO3pd8Ty8xgrzpf1521Fp7TqT5UJq2XxHUj2v9eK1dxFl9F8bi1lg2
mF1hDnNytF9H8sKRL1FcSV+ysNVTZpuIdv4r90jmKTCJsX+e8Hpkkn8wX+T671xUdqOWofVgka0u
lKiOG9GrB/x+6nAEsthsBnImzyZmSWPM/P7Z7hxfHDxaAmX2l4CdDtAp9LfokTOvlHp2k0c5MkrU
8+RMNt9xcCql7ziqHmt+WzLI+xVYURBWkDJEZ+xdV5IXsDzG42xghDm5h7R/kaGj9AZ63YTIjYcs
yp5nJO/JNhxwsLAwd9hiBcCcbsSfkbS8aGvgeRM/+8lurojURKWs+LOZjgMz+NOQIAFNA0XJhtV4
8yuxR32yeCJmQ30lD/aYI6cq3nXfypvyiesFGli+uznNMEx9artIyhyIHvX7PdlNaXNTSmh1mJ7S
EcAFNoFUVR/H/7V4ej5LSXot4Wd9F+XL6dhWi31q9vb0iEiW+8XKAeQkdnXVltKBcpcZwg34ZNgo
sb6CKWosl4S+Rreyw9sLZacBypfH3o5eqqZPahuOwHscoNvPz/gNR1bqICNL6MtihuACa5uSb9zY
8T/tkgfz7d6ive8Mb21QMsef/mtdzyzQ0rengF2b6M6dv/aXLKde2ZFca07KNAw7MNuCzoY95aBy
yhkdcNmBrq8N6+C9Fu6gzMsmWTRNV2iDc5xRXHl1IO5VkI6ybESIbxnHTcGqfXLpZlhWf5ZVS3YP
zGIOH41trQbZ8uTzU4S+ZzhLoaa7h/aHNKTUXR5jS2NNf6AN4egNzI8N9c5hBMrmGBYOXJsQ80fc
vpv7AgMQAg/97NNytOVhMmGpBZ6yozXx+3Mp+ffUIvjEL4k3qkrhLjSsQb23BaGbDNGDhu8fzpXD
cSPyoQI7Vej40kvSqZwXTbo9lGtoZ73oZblVpw7/3QhcGjERNMymo7N9UDGYT3CJXS9h5F1LncOM
ho+z+jmITGQGhE2qoB8GljuFjP4YDFu6X78rBEQOt6AqdZLlVHDPMcVM74Oc5BNQdmxRq2w3hagp
83fDFgqz+6xKTrbdHjWbVxXYWF380iQUq1DrYJNS2gmjWX2C/dRDa6lexXqrXlBOAE9xpU+Dp0SX
nGjgW1gZ3YMw8+qYOr7FDDYqeKiMQ7zZ2lPg03ECwAAFHt2SZ324EY5mKOV+WdfOLZ6/twfzZyLt
3pAAMMPLPL+hveET41TqlIC4SXskTymzmW51Gkybp1fYSrP8amZHSSSDK5U5aN3xkNhjMNZ1u5Tr
07mb0PirsVzIs4E01BwxV4JYufRqX+j/9YjtNHs4/KFDT5fPsio15yCTGAJnTkg1iBlEoghGgQWq
rujiSfxZSWeLO/oFFec2Dx6WFpxoa5fFlOXnGSwKUVoh7jFGsJBi8wPHge8ceidSilSLgWsulUuU
eDUAOlEUH4z2coJGkyfmKlbKMoJ7Zp+lSdRIrrfeDgRpxdc7foVlslsDHw9Q2ynGhRrao2hXwLmE
dHaunJ+O/GeTSsjPSsywTeScZ5lE41QdwtZVYVQ/s3VaYJZv8PocDoOZkLyr3VQsipE2WaZ3DsL0
X55okpAbe5bG1jU9g792uoYUgPEFLEvqjAV4bmwd7muA+DKstgjIvrgCV7+tpN2qJqzmDHe93vIA
4vyds84CzxukycgncJH6zTYvmYfGXLJ9q61j0wGn8kyrfzCbHVzKLLEmvN90Ro5Cd93xYJcJpQ6C
91se9eXCah3ilGJfWMFRHqS19T+WZUO2l4BA54FFHeXNFTUbnWaD4qTErgVu7Tn8um/3k27KkYfe
Rdpc3NuFwnSd9NP9dqRpb9JNte0vejMDQ/tfqGBR1i6diksaqOiQqQIiK7U+bhm+Aj2euUVfF4dK
emFqdRAtnDN3CM0gQBbm7LqmMXCsMzSzK+9oRH0J9lbX4PilEeGwdvnCUrOf142NxH303+0i2qdV
X9k2rS5EpG1NEVeDXHBN+Uxk/MTJDPvou2yJNsKt0iaXEFvbBEArMJFaq6dhfMvAPLSfyhWwvdDf
nCU5J7hPgvIRZ02U/py4eIzegDK4/EBsp2zVavcz3J1AmCf0bOunvdQXL76L5Qxh7ww0VdGpfqWY
1rLLySAsP08cfr3BNGlYp1GWOISJC8n2YX7FH2KJti9VkLveh8JZX3DMrWUBo8IuJRxnCEi4di+i
zeUsUAH0z3N94kGylP/pLmpMaVeLXz8RqaRI+o5J0Crnbmf/3QJxW21cidYmta33FxQuAnxTqSTD
J0Lwtx7Tn1NQv/lL0LWr+M54roAMCc5ndELKBoW0g0h8gUdms2b0/sow56eil9kXNAWxIac9WoEo
LJcAud/PsKfCSaYei2cU9ymg4HRg6ocEq5wHuNSYGKx+xXhO6q4bwg4ko+y+sM1+/5G+qq/U+0cw
HOrLIxRu1iuLp6DhWDY7ulNRLpHCR0IpBKxANSyRtjZkSq6HwngfDQuCEpgEfIlqwmm4N6WlXJQB
X7dP9mXgN8z31fA4y/t5xp5CYAiSQO39WQjtNEhh+mykuHlH0VNCs4PEPmxJZNLxDzZpipCn5uY1
/QFaeV2H05DHNizvsEF8T6KtPtq+cNlEHbLGsZ4uFDk4oZ5qLiZNMsMwU8mMAvUCK6JLmz89h+E9
cig1JHsGAWwZsTYXgplZiNwU0gBqeHXKBdcwnuPISiGxgaK+VFCe0A3oOi0dkeyR5GkmPtnTW/cm
DbK2t6RRYOF8EwBcNGO+82lbj9UN417JvR8VBg9Tf3O2uuuUve0wWFFfP/PU5RAsqhd+by1QhVVd
wN+65h9JyXW2ITnjn2emhHxugJajJdAisnhzT5jdBWsHiBIRUy/RPZL5PfFQrZQtPwsdx8zO4FdV
NbxRP+wdspdqo0zJ4Uh+muDCIZZpPRNDOhKx/6fiJ3aYoPlG0SqmAHDhRdysGHMdL5PhoMuU4qth
ecCZVWHdrmEbE1T7CmMpJ3JiQeAsZ0kVB1hKbBArQtUTc0nhzZbkgrDD3xSVKXqlZNpmQd6blkGJ
kUNy84bWXdPOsqC+U3ToEOqjTuFql1XwPFNxmYgHl7GEEYOoPR3blXSixDmEFe2FCugGR2vClGFs
64VeXbXKpt6DIJu98amFIeJmMusALpRZjwsBCkP2cAxzZ/S/MYpcQvfivswSCxLOjFrfDj50+laB
Dba9oo5yze9nCabZhbM021aETk/IyOOCaPbJOfhRA5CcBCapKlo0U+qWyAvqLyF4yHeB7ZkbeiL7
JaM7ZmbGcSmtasdJbOwAoMulEjK9uWeE3Y6hbbJVRSnPQQWH89W4Ihtg1fHEAyGVuIY+BsPZyR7i
dv2swVjLm0HRT4cgiDi4pTbkK6V28v/YJx5Ia855mzEkT0txOYoG/aAZmS+ceg7c4TZq/qP5bVfH
ngMwKJ+bWn1L7da98/5QAPLKhfqFB5Eg1n28qcx7MyxBbc5iRcv0OQnDglvAcDldPX/DdthIRoUz
Wr3HuSOAj9ApTY1FBrEEPr3FUnVT1P+U9JIF7kdCQZ8CKx8t+iWK1G+RYBEwI9I38A41cTbRbWx6
kvOIE9+y077lEVOMMbBlUhcTOzeNV+cCgVl7iScXrzy8GHjB18v9pEhQgT2kWvqDK495d61PLkln
Tk5y4ljMtzFcwQyhXH4WVCBox8SrONlgNZhNqK4e0X2KqhD0XDYG86iAkJQq6CcziKqzkWP/o576
TLZnJNoEKAABTXlCNDBnXrXYyBAp55X0Wlq8eqfLB1vaDQaPgDBsO8RIaoN5lYnEd+Lo1o7VQ6c7
KdgejOOOeyDZATiU+1GbtysOYrv4U9TC6GRZDjpMyycOCpM8dDGourrlyOBVnK61mMv5qWqDDQXt
PXoDd0rtsysGv2uUKnovzJd9TXC1zsjP3cs1qrFViiyAb1kX35298i2mpJHZChf12BsaLNHvjQeY
a6petS3SRr1q+Shjm8zsO7WaRV4f70lF8aJ+0oo9Ud+pfGywqtNrZfPpI0Ugd0bKfagdcdp3X/iA
er2q9b4cTmFet3YiMuRPSxImT7comw6brzobLl6ig05s0JEviLKPuYNP0twL95gfHWJPp/yzWN7G
RfcVto5sQHSEcwAzPFMN0TJMaiYUMviat2SvJDDDYeEHRigNb0wxD7U2CL7Kw9QhADiZE8r0SoVx
cT3YxJ8TUW5wMiEJ+nWMMew3AByz43gPmnH9bwYc9MHxcjPJgOzeVcM/vPPJrLfE7wa2R9HB15Dn
szvfrokYrNTMFSI4DvQ6mcBxY8LAopokxb5t8T3EISjQ6A+Bp6AOEoXIyAo1ZTJZf2GJpbJmA1hd
lVG1H/WYZcsSt7LU1PkFJTVhmVvjc1+B8IlwtPrFy7ujnJySQ0Fowwea6TKdjKaGA3KcyUc5VFSi
CIEpblOZX0Ur23rsrhRGAunjdHSvifxtSOOkK5RV/7Wclhd3aLnGPE8DntamwOMO7iVHzrUXN6qe
98j84DIY/a53K0RdET6XzDQeye+fzt3YcaSqZNdo3EpCBT0JIEIJDlRbfUb6zU2OLAahi8Wf7iha
by6mVEBOS7XOozLZsuAtdI7PYxh2tpFYd5pwjM3vjoGyHoLxO2/fUk7jAmB0c1n0HLEjykuIbPm+
nhv5uBwJ6mDxb7umSchGhlE5l8eboNPlNfX42e35x9i1NRqid9zIRWowXOzCFh0tcva9n6wua1zc
0+4nBlF17EuxktRmeH83x+lvi1EHmIZ5pmA3JpG/N10FeSHKFTnCjWGPsSgsNTGkdyfjxXmGDt+l
fDqgo9S0wLSRaH0kXuIXg8GkMwg5NCpp9z0fSyOgedSsWtj9jaQTfSyGhb3rcIV2z0SPU5cPLJml
9lqbEKl7wRvnyx8NWBmyyTCl7OrHGfJIlDlsRi3G5KcphuGa0NwOWjZFPg12SnphGf75WBrzwcEH
PNo0Qj56XvpNlRByYbHEeGLo9cZl1ohjxpVET9YYzCr5/mIZ+477jRP/UYiDPuYv7XbrK9hkfPGb
WdMdzBth6UXo87szrLMTLGTWsHMBhOabnSwZDSwOTe/6Xmss+BFJhPOlDsGqTXzs9AI4eC++B8EH
sk+u2+QpossuSlK5yx3sJ1hAjq6faErcpyjkxpp3eb3Cu84DAepwFtWg651R1D3egtcGkptNIs5l
5CMRPXx7KS1h+GNf1yY5mSqd5+yf3W7A3OWCzZwZkgAhPlcHF83GVUhJIulEla/l9yUrJC4fTUjE
7TKgNNjTzp85IAHhDuucO0rx4AtJu+xEEuVq3I//bR1powu0re3QPfQs0ixqwGvOsrdSRz8lXtmm
8NIKyvkmJYNUeMXHb6pPLC4X2vRcK1jD4AJRXPeT2DDA39etd0AVCGSRds4fbK6uYe1xQeyQaDQR
5b84PX9nZyqis3xmwaKVyIXjqjvV83W8FSGa05XtNXKMu271ZZ+p90cpiZkYAxUCLqhnmYDF1fTv
6YRz3jNaVCltmdcYPXgwrNkSvWXWdrLnyByG44rhoroOz3BPTntfYpS8BdZrS3ajk60gFg3HP/LT
Qqgu5TJ2pmsgXOC6y8IFqB8T+J+phLpYqYpf1SrKuc5GE4OGx/8teYLVMICN3yGAIlB4tScUKTNg
uC8hwER0nMDdgGuHH8vrqKFCDc9fXrtqIr9T7cBAxgutKY2rUSFe4oeHiGJm9h53jmcyfx9DAvq4
F7Q9b0Nu2HU93Zi1oX3poiKQwvbDZLyguxxhC/FjOgIM3cdLFaTraq/zkvRcozV8wUt2y5bZHrxM
meEFK3cQ04utFaHzSPkW0KV7QlZqhlOAL0n0G+wfvecM5h6ywLySRrYNoZ4Z7sFxdklMqoXjnTh9
gRiKFd+T6uXY+SQUURl4ev+3Y8Ks48cFR/3afYRoiaIo6H+KB/4KsLBekEJipMPkciqCJ7Fp+b3J
EDFPdemVHudrDg99ro12vUBQLQhmSVBbf2zw5joCwXGJX87E9BnJXGnChR57CdI9lIztbY5nRZ0S
sj9lAekLEw8/5TydAFCXrlltVbl+6D7eXUILmPvwgvZBfUKlr6NWiE/jUWZNmeQ2XDhF7R1oL939
eVoTppjjUyc451MRmlvtiUJS1aasOpfXrWibyZ9UpqqW1QwbZAbYqwBz7od1YWr+LRcFQGooSC19
R7+L+aMJzlDEiAIACBI3xb8cjVpuSCgHqH+2UrasBIEWDbRDy0FoXBPwuEVXQHDFeZdLDHJhOYo0
kw+nnK9PTIzURjzrqTUcuurXWzsONAi/VrOtizYXUHBQCGxMXywXDlnzldJPsc88Bt+kqDVbpSZT
V3zdCgkJwXAe/DNdxCHzjSJO/+D6gprVo88eZms+7gbynkr46UMTxz9xkoYhkp09KBA6WJE6Ohpk
ODYc10PS5hDOptmC5mJa2IAoQZdY/m5pGRbyosKiABN/YMEGqEmnNa2ItGOKiM23ZgoTnTwNg0RT
6/HNnQLcNq5M01cjDU20GjjlIELBg8Ihwvxri1hyYLtOLi9w26khM57ccfd7qeMS5V5VChK+m9Ij
Oydn5jTMC8/FSEdW5JjSVH6/RQ4rNXMjBjqmqeS6U1Eyc5Cfn35yIXv1ez9zYbJafPWNrup0q9UJ
YZhQLWJxkdHgKRoIqvmXNzW3zovPleda+fGKLMN+Kgu/iB6nW4PFlT1fsP4dDQ8GVUD6ycGPSkCj
X0e9k3/MCXQTzXMRidukXC70JogYUM8fidR+TwFIMtpN8Nmg7cOei+03ETzIhR3ZSVItPaytwvE4
JzL6ih3rQnPbACDzX0eQIDDN0pJiVwOOaSFSCDkGi965ioTxJrXrnyo3TqI9uTCiWuQj0W9l+uXG
pZ/GnZgTSgzuLucE/MVV2Epp8Gmt/vi+IoCr/cX3mMkfxDcSrXO8wB0EL/DZkqWnA0WX6/EHq/xS
pRiS5a9n+hy0w83bw5rcHU+7AR88RinJYg5iLVL3NQaG3+UwNEJfOJ9MUP/SHE4eeG+vI7CWrGPz
ifQWbmfBNuktLXqU6cNRhpUG6ZpmVT2WmiRDheJcz2uaPWKkWJEK2sskIIObcai5Tsk+b+ZDZl1Q
Rl0FBcSCjqufvEgdfbNMNJjYN1SjJX0qlFDPz6tj0BuFINyN03RvJ1tg+YgncpxFvGMCql6hAcFl
IyN3jcZSMkYYrDn3qp1VTE1VdHTTAR6gaxQyy7PwKH5ApU0MUNJYIvd2lU/5XF3maLpOW8muXB4u
lJ+ISkZA9it3X5qlK2se9Yj3QAgLFHL6aPIlOaDrAzfs1onOvHecCzQIy7v7neYZ8C5jnXvkG4vt
oZNi5Pg67DsC9MDgsKloV/Go8uvt9zy+XVUw/5socsHLcFJvNDF+1c0wfzwQo5OrOOT33vu3ZXbY
73XpfiSJiBE7WCl9IwOJqgQycoS4nI1NwIhOfFdP0UIRb0T/AneO1xPjGkjeCOTnIQBOG4EREO/w
K/igfc0ee3tNByKAS3qsbPjfpQKgn8uu51CVUaFG1xkZoz0c7tj5KNL1MpHEwpakGVK1KhODF+e7
JtF9YX8iMV9wFwx4K7QBGYFAgVPyystgYTcnnOdd7catRzDTpN//S6zGsC5f96mLHmnE4T2hiCAC
6GYTGQsVDDpeaLwrsZrw8UmwuhJ5WZ01b5PWSWTzm994W3gxDIAGG/IOWMXlJ5E6Ozp9RVfuyfIw
NwYURj6ApAXjdyJcNPonh7PRPnQHc2ipKglGRGVWZs16/zFdK3ZoNTl63PzkMUWuor81vcxSh32/
t/GmSIycPE9euSGV08MbM5kfZmjBjskOl/N2c1iS8Ajda8VBbOOaaUW44F8a0E+kZ+Y5bWIy0YnF
vzicDeVeUCZCM1FiTRkLS95CUPv4dLQCOl1/8/gAc5RLNUmmkpG4mukvm5Jq0WJ2OkDy8ApLYRsA
C3xPpJJtxXa4DdBItGgmCVG/7FWVTxgrA4gCTUp/ByAXyFZno5CrYRuG2Gku5M5jAqY21qDvnoMg
vmL3FEGlAdESiomxaCwa4+I/mMhMR2BPaYW2aHRzcjF0Z6iuWp9VNB5wmhRVamB4+bf2/EoLZhNv
qsOAY0PeysyeOxDC0zn7zdleLwYIC+Ajx1BPsSJ+UbOh+fTF7lchP88Fbxs/kmMzoU/MCaczV+ev
k2x0gtoueo159rXnEFqTIuGpAJQyrSGFDEYNp80AkyJD90aA3kDxzE2Ypy0kSKszdUVu6GjUot7/
o1MEAYHHzGKpTiQwtKQiYGCg6E7ZyI2To7E2PTZG96DNnS58Zh4FwcT1Q6ZGkjnldVF/J1n8q2Yt
lwWZn2xwXWXPEeHQvesAyR/jttUYOX3R+LNOYqRjg1x/UJeWvlf5uv+K5uEz2bIin9pxH3/G/8kC
sqYfzy96+Wm59w9YL6GyJAredJBHKo7/OrpF2dmx5LgTRJtPaTCC9dQFTmVHd57MdJ0FwCPNMdAD
+tYXAVEY6T44v/v0Ke7X/NxzuuphT0R8EtTlt3b5RBPJXOjqxUGasNNUbuVwTN32XIXTCcPEx0h2
VZtsLUvESMXlQtqMKlwYzjjtQNYe4tu8zxhw40/eJgJ3M20gkCPZuIto+iP3NlKmEISVm8l3Ywrm
D0QwKH6m1jrgPZLc/5KHiRsfi8lO04c0NgdkIVxfCqzxSySQh8b+7FoNZ4IXvvjnw1BPS8hi7VvG
cgXCLqaI1eHVQSLNypUSSxOScAWGY3m4EsJyXbR2s8LNJX/G8WZKlqy4KObHBeK3JVPGm0bNj3kN
4hd4qaJ/gbM9xq+5BQqVusPE2NjhD9K3lJ5hTZbEdU97Yp5w/lW/C0sq1Sk39yN8xzYu99dcpUKt
3wKqQ5D7k8mL0gCkveJu3xaloHk7xBGgUSxlvjm8YfI0i0vBTt3yYHtn/b7GrQqKBV+tZNcjP5q0
2Z7vlWw8vMNqs/O53DSiQwhhqkeyPd3LI+8hd1Csdl5poVeQectXvb+jVAUMEXjB4ec+7lolYPwL
hPu5f/uzfnCnhLVL+EtHhmQJg/3jZX4lm8EMPahCtvCU2EqAmKUjz4p/5ymiG6xKmCXe07ZHHtOy
O7ZjoeREe7fFXFAlU2y7NIS3E/Y4bzRQ50u+gwyCN+VwFyu3FvQJc9hXw6rihSzuF0bEGSRIcws9
vd/yp+Pvpa8UYPvw+qkVNZlNVHuSiH7iY65X156O9tiuvZzk6Y/GDN8qRfqmZLyjfZ96TtUXwlgC
QjRi/qCLCDF1oQMqovDec552B9p9JHc0kXBCIb3L1fBEkzRWxSpobisCfeHft0wnm3lWLQ4unGk7
xIH6lqHtxPaYUcRHQhwEWcEGXLLNrq35UYwV1FdTJgA8eVWMCSvIFIs0v3hcL9Wz/pr9HUDXvdQ3
ISctnvdWC7hp7G2ntm9geRPyedg/oKAgCog1CDqsLeEgVMnRENZ2fwiqgClo9G+QqIaAL6buPFvq
jPAk0gvoFjQliyCPvHF/jZ3ve1Kx0pf4WW6u/0Gn4FOxmiN69hs06egdHcRllEMnC/q2uYJHxJaG
DBWZ4dApRYj/LqsZ21cnAuzFqDHPKIwQjQgr33PRwW9HjxtQUIgvd/L74A/pTYCtM9IXZ6Y/hQXd
eZ7hbboC+9T9EtJG47LATuYd13lrnJ2Xbt0yUPXIgniWddLCvWuiX4wsTRbCfIPQFv8xh0VCp8rl
Ok5x5zAHvu7FgwW5ryxInOmYH2Od5zxkdwqa8WUmkJfOWsJClRQx15n2yc7Jj3CpAeviRQdeR0vd
c3oL3Juw3NGCDUrjI3cW6x7u6gU2/m2SHp/erzlqOsjhAtnyVqooymTlXr2ie7QCTgrWyUA5NyWR
H11FlAlY5dABnK4phYQKy21dzax3RM+Sy/JMxl2AkxX3czpK+DvkrDB5RWYniH/bJN4SNfBsvAUd
vM6dA6bzd55exuOiWayML0UGdi87MpdpuLDizZOQp116giSxQaaVEUR5/JEGvkZ6+EVW2CQIUglw
vo8sYPkyJEkMYQvBq3OLpG/6YkT2f/XjbMONc9fX93LulIVyYQkwGJAqJKrlqMVCzye3IJszQ3Tj
CBAjmjxeFbobK1pchUZvxMYF9PmmqhIUnuiPdTIRn4cSAI09al6ZTp2ob+GoTA+1nIBf8qNiFE+7
ijbq6yhJ6wFnw/Hna7w918fXdQnGhdRh671+c7B0C57RDYe0SO5tzZ8rEnCyXibwVgIUtBqE5CfP
Y9M8QwkHPqRSF4HozjAXVRA6ZTsaNXUx3X5MjvlGSlzFjIydpg+pVozl7mr5NRSD71PwCuecZ+Am
ypJpX03a07CYcsVEq6wHBB+z4CoMmk4stNoeThYfkDIzgdECP2fyblu9CmEssaPuZxItLXGnahdy
vaUW4TsVGNLCSDwp9UOQjyNuCXu3ppx4836SlQIz86QuSloG2ktks1jFGiT7VhW/girnBPySQXIg
h/n5Od9lmQ4TqfDrFUlao3969vu6UiQ2gsEStYssYBH3bk0B5uPvz1eIhC1C+IkDc9BdogK6B4dH
GgNC6wZzNK5ezOVy8VeZludTLhJ+SfOXdY7c9EfhxE8GRUYBtZaiLjXQOi586Tq/VX5yxRsoULFe
nCRp+JaSL01haaiKIZT8FfYdjBspqj8iroD1n6cYGEbKabsNKGnIGBeIkDSCnI/w+Emd0fVDIr9M
iBdD2SdwSi43c8vZjGL/YJOx3+C3/uWxe86Kbczu/T52pdwfxbKTbk9nDAVmCwaR65HudLX8idyY
kryN1BF/gfU8pkFNnQdGZpVsT/hFBhw5JQRI3hpuxfgER3QclkfdQ66tJtvffsgJ7t7JhyD36YTA
ajYWyc95pp2et85AGNRkB4Q7lb5MtAKFzc14vrOfDECsRR7TrFIEFCJwmMD5DcxmTBmd+KWj93yS
QzwwbjtSJcwIMNxt0/azV6nWwAzVkdtVCzrMAR11jEL45BFLSnNtNExEOwyfrvEgwsGBrrrcqm8U
gI3CTLQsprAcutfZAdty4ksVot+hScRQrP4aWMArkOW6oswiA7q6mK/GUav6vB/DaS2WIEqLMxm7
ZIe4kVbz1kKP0aKbSXabgSfZYl6N8VCoPiyEX5Mz3xW9RFmLCM329Yig4eAzNMEAFyb6F7jDFlkc
TUpMJY4z0Ruj3EHrBP0KrMg74Kf7BzQ5Hv+8qEjLaxc79A8l9v4rdw1rn9qOtUFMceeJbI3Uk0lx
G+WjBt1TGjt+o/AlXtF0BtDuD5jBkO+MqPUMLHYhBBfPx1TenzEy3A+Sg99JSVVZZPmo3m0VvKOt
hzsUsIsi/LJCdZCPze7vra1uZxBjyHIPaaAyz95+vPAKLBEiGWSE698+fIMkaC6fOkxSI2r6qTEq
UGSf4HhlumsVWGhI67k5+AYXy3oRLN4nBW4R6+ZZxgYX1ILelnap0KzK2mVFLMpAkKqG8RvOgWm2
4k8oRz7fEaWps/p/yT3Y8sDLHIVaJxcd7gP7toJ43jzIRuOIWddjahNY6lYF1tH/U2wbgoAdMRNy
g8SV4AuFgng5HoCopNwHRdF0TwUfZEblK1X+1qX+GvzVn+MLXRBqx1J9PuxcwhVKu96aOw/LE8de
auwwHoIZ0A4GDJJj1uaRu2AYMwBRY64xrwTV7ozKLo7r1hYMTbKU2/+hdCBLgZRLEIGvh2bVINhl
93Hg9Byc2EsgbF6YfK7NT9HLOvnELcOQG9KYXKBqhqRABq/aXOB8ygJDklT11Zl9mEARaMF0Ytlz
5H7H8GG7GluMuTVU4dA6Rk5p69p1BlvxYzOmD3n/3fggVRHjsNPpPAADc5AAWmTOjOEFm/J8ODS4
/4F7c7J455vF2+F9y11omJnIL3XeoA7FURwv2af7VMvoWu+9bouXA5nsK0LKN6pyXQDZFAe6E9hs
lpOQKeIVcbDiWY56+mwpVW4fbgMrZlemnfsQfi9j1Pb4a9EiKOw2b0qnUBIJUJIYd0a1dQaZnKFL
yxMt18z8qkSMZRll2WPTzV4ZKvo5Lp/NphR+fOTBEhYDrq/kIRHsRgvWlwLLmv0U5LNdu/w9Vqua
/k2a0OdXzWsVAVCbI1eI9+VJaedgzCoF/uQnKydbSuLPQ+CYYbaOl84I6LKQZF+pt9BynLdzIoGY
LavhYXtexrCdwbrhpakTfMqaoVEogf9Dpzizxb9ZwbwmA3iizOgKbW0jeLI+zAbR4zfNzwoo+EdN
M8iPc7dnEUPjD2VnHWyYyjr735p91vAmt3iGkG1C67VHojx2AD3UvDgDH6eq4J0ykfVRnujiiLXS
R/N8Du4pqikPWQ3zejD1w2np7s7RxjwP2XUetTz3BKto3vInP0wEPwnra+5d+MhOfOfzHOnFj4tT
8JnGSjaSWzaf+rWjQnsH43adyWuemAFjZHUiEmL3KAVnwDUOKUIjK+2q8YuiI19OGSV0ra1MnK/p
S0sjL5XzbxGK5+R1GqsmwKIHA0JiK4sfclpK9S7ZDVwjjMXGmyYuu2eyb77QnV7mr8QwPadwoLby
0Rb2wiMUVhpdfFhz/Kvo2k7fjqVXKnsO6u8PZBwc9L+A5rwn7sgAasYMqQnu7rqRh4SUzTjGhuh7
9ODbNMbZtAYa/jq0wOTDceJ0jPTS/MgwkKFr6WLgHyNF4yVmGDUHhhRvFp0UilqLiVi2iPNTmmyu
2ksoRrS12syFVeNgQsPPbD/T240Fpam/TR1Qfqe+7FOqAsBXmrHUG0WqoE7Q8aUry34pIiG4y1CS
CwNnlZGcvenSCkyuGFc+IhpryrewhHhrop7XdsSk1eUkDt8BKRLBTldT/cvVTlr9UiSy5mREXgf8
UwHJuRs1Xben8X15h6OEdLazHUEEgWdD9bwjVz9l1GcwJ6HC4yuXuR6UEhRZPbnTz+6rZ38iULbW
ABZ2fEyIlVPhUQLa4pwDdoiYStbJNLu8Bw95dt6jcO7uzry2FY+e8om4VmtYR8AWupOf890DFtKh
fy4xKMm5EEUye3b53p8iPzVAxEWHBEx4zto5lrj95sLhT7jft12umqpmUM0f+LO7q4jDRdzcI/7I
UhPSdCzl5AWkQlaMUW2LqOLUSDL115XX0BiQLajPadfNnAe3EIKAZG4dBRJDYPRrbAZAY3AGWNKA
TAK344bvfMSrpMvHBcjkCDgfKQ6q/5ob4Ch9dCoa1gLMgPIBwpeJs998E6tn3Tqosr//xu5DPhrd
7hrEV63zp0XDClPQfUP9iCwMYicAH3HVKfUuyClTlOaguB9/cPEC6WREVjuO2txVgrKzV01Xj12Y
bGajRbZMbW015U8HPLWVcJ+S16WI4Cp9EFJ+OEcP2j3Yl1RVe1KuE/t1g4xuW7T494F0U9FtEPAQ
LSF5UW31n8ty6On7fK8V2E2ujRnuxusPiqHY6qnmNuGFb6gZMD7fWysrfaLnOe8Z0WFHphaLAXJJ
MXwNwS4tAews3cis4FL3dZ/YoKWf2crPr6mUyltpqcTSSKE1v4sHnwUb4nC9i611saSccx6JgR4Y
UxTm/0anBQtdYbHPy4eThAwFunQjY7nVCHyGibxCzlBCU+GvgAtt0WCP6iIb5BeIyz+D+HUwIQi4
59lKY36x9thATeuOhm1tJA/gYR7tPwTxfl8RtQJHOZRx/7UGKO/rPO69uigLMQHSl4QfaH+33uWe
7eo2aSuufuNFmSsNncKHfWse8WeJefh5CRTzB21BwBkRhlf/xfWEEGBv0lfhYV7pq0EPOCAuqK6L
kilbmITHUTSzzO6N4BKRWIf6Mo9kE8WtAdMkQeMPFV99VcewhopukmUp6Pbh6/OoItqRurZDH7a0
nv+54hwGWg47QFcl8cebmNLseBG2Ytk4aoCNCPufmBDb1w+luJty4JvS8bUcRiduAfHEJ5iuqncq
P2/gbGZKiU9eKoMVc1gSB0atyAFYgk6+U9z87OsIdI0Djc9/5JZR1rRcG6g5n2n0Ugsb9KTzdfiN
YEchPet+jxck2Cu8M9sV/8VvRlIBPgaKdqy0mN8p1hF8LQpOwUpbB92PdN1pNxWdCuz4lB/PRswL
6C9BbRtNL5ta8y1a5FaxnGC1vVbQSjjJbhbqwgebfBwF0emPLmVMYB41FMQoGSG+7OwP98x0ou09
X/Gxq2De5SjSI2pi5YzVXPVCPQ8ln8r2m+sYPotsew7XlvVlElQLlqv/6j8UM5tG/jcDX9b5mNdw
LlzH8kpxxMxTbi3QoD5elRRLZQlr7T5fXuVx/OZ7dGcDMeZ1PcpPc7Ax1SwL48JWM0scvjyDZ0BS
yhHEAH5UnfF71kInRiZBbtFowBBUE9c5IJDqwpp7YOcsqfAk1PeMOXdO7vGzNS5yVFyJJ2aY14lP
dC/LlPSCabTTYM9q8ugOHNUh/PNud7tghOq5QlCLFZzSqhaxTzMDm/h/IBerjvqXF87WXEliwhFt
pLDpZ8uR+2O5gmre/6spVzWTBBWormyuDvecQZZDLF7uJJAh5I1oi6O41ZEod8wNFjv9I/qyWsBK
GI4R+1vU2wjJMQrwProOcClCHExqRun6t1ZB8G5rbV7pRZXPKDdFCJNCo7yQLzMuQzltVRdl2z8U
FsbpD9k4bIf5CdJiuTvr596nslNtR2xlNNAfbZzy58ipoAOykjw1ocDcVCJg29bgUziQzYCvYCGB
xQoBjpAfdLvIEclIsHhq+azpWJoh5FIU3pUo97+vodXG0YEbm1r1noBv338s6+bsvcDZx24EVy+f
T5oR87l8BlyPUvrAQI/TWTYrcbE6phNc5Uo/LGDoyxm3JTbr2z/6QmpcE69h9pU0fZLYhTqGi9cO
8zvcY7s2UUVZ1XWCN/NvWJBsEgfHPwBVyxh+uY4wktCJBHDaVOZN2BUq/7fS6JRpcdu5MuIQNkw3
0GSg4p9GXfZpQs+AyBd13TkezbpCedMXASp8UqjGWJ87mCXBmx0KIubOG5V7na/VZxuCH1npxw/X
vNK5f/hQ3UqXwVU9Hbd0FM6p0hoBNNZN4PNfpuASoO0du6YdLJbkgDamVZPTNCc6T4Mslg9703ot
x7pVOGG7gcYDIdyS5nhsIPmjLan3XmJpirhL82U9A8hqYKk4TvBDBFfhqRXuZeGYhVwbIYRtVPUe
Ha0OyeWI1b3mzDfIZBvQaorHLqPL+8I34rR0HanNw6AqXPytWi43N3RKbVFYs6o0FWT+l5IcD/0I
WhgtSLIB2E0SF282gMltXI9HPsibuHGLNNC999yM/ftwhrlx2LNjUfK6WZ28odmsWaLTZpgutfeX
JnUMiDCx6yD5hEsDJNmGtj4GgFRMcglungXWRyc2U94YEqYIyjeYHk0jX9rY8b3uYrRrEE/8SaN2
k/22/Kvr8XKzXEsO31YiSKvryUSOnajchPCsallJOLGfH1THTBrmaTKWqfjmcwM/HKSFHSikcJqV
wknwj+Ekhf8aPBg+to8w2mzDYxGTbcvsqtEVx7k5WPg1XagJUGq5EttIT7XTc8yN2pjio41lpqcV
sy1jVVAEuQOYGtvwzA0POKgoRG7jx3oK+IGg5b4zgjQUn/xuz0bQswW8QQ4LY7VDCnpPJHnhOgbu
mUg4ElG5+yDkZY/yJWfwxmYtluSWbaonKpsnL5Zn1Omy/VbEj//omAQhxp8lc3HtQpwSjUGte4yW
ahK01k6Ss77ocaviLgDbae3tby+fYD94qph86WkVM9B1PLIrooSEiYY8bF+lruhlLHmGHpl7mpYO
IlzngkKia7p7+zg97b49jxaegPvQeNCC2hj+9j23czEL42BId3cMFdrQM7Z3P7WMRNCvNTTVGkam
fX6S95WNkcfo+IOOjuoSZG8A30qF9aNKR7KbCOk406BkVBB8dKXQzTOZFfhLFffhRUBYUZpZyLyV
Z3S0V+U+95LjYq3VRBoeiGmlFH0piZbSnQRgU5bbfv+I/kCPklykDp9hWYazaPG6muBpAUdnEqva
KcW3wYRS54da7zQOcaHL2mcQ+O0JZJREFwgZfP6zDy/oEzfZjbFdRxXc41e0RPoDtJpWiMBerBIc
TQfVrn9K6j15pY/8G1lqH3MAcVhVTedd7UcQDVLC7s2LHT/0aWwCiqQW9lqiafqBBepFmKiris5T
dv+nexFs1JPY/jN0WxkJQvResP/uGDDF/EymjQiu7rF/belY8HeAIz5B4tSL3kejLcEfS6YRxFam
Cf8SwHSPCiSeVlXG00hAfOK0HlZOjRbTM9iwYrqUjwehnUZMc10fWjRcmvgg7gclqyL5ubDijXZ2
EiUALcFuA984uPGGdaRu3vpJ7fwcNYvE1HE3XmgBJglXek3yIHwuAipPv9GymDnKDtaZgQ8bchlg
bszoh60ckK/V1epgh0n+gt9NNvlNpsLrOhJBBjY1Jru0IljeBnxAVPalsdWlx//QnyaHh+Q3+0KM
eO+Z5tqMn22LKQkRIBbOpR6/HYcOtfecMHtkUCn/98bnHrF1/K5yCAa+BvTW6TnzBB0z9PI8Y24M
H4MQ4++txVM+67GZWmXswGgBMTlvhS6faZ1xFDy1SpgB2IShi6NntayQjsAcssLj5/KhmXER6rbL
4V7rW0c7nvKudRZVuNNEmOvQ2FT6eilWfSpd0It/hhZX2G55zxx0pOYfsaLBMrxkxYfBd5pqECFA
LTxs6a22ABM+yfaelmsSUTfZmFqRSWbLcLyuSDwvIbf42xxIdubSv66c2v2NflKURDcrcXAvljaq
dyV7H6djgrLHLy5qYisQh55RY2dzmht7ms9FB6Kf+ocEJfCrpkEtFLBILCTbbNXW8aY1GggakwWG
S/5LMQHIAvCaglmJPTm65+b/9jBPk7XjX8bP5OJbkHaXgJDFDeB7ATzICaol2hutEp0ejjLtoyNW
RdF8BKReWbtuaCwc/TaJeFfqjPG+0k1cOvuCIQL8ioNCAH4tzVae7terI2wjNkWUAHGA5PScJ2G4
p5DmxiMw7NN0bhDjIsYLzuj7iHxqIEItWZZbFH9cTYhA50DBtjePwI9imSo2FVRMPa1otZmWpAJX
XCaKwERpPijduEfPF6U0eq0RJ6x9vB4IBI2+Ry8FWbwvYHhOTgiUYHhnpzo2WzA3CW0Qm/Wdd3qD
njNPCbWjqAuFG2mxl860TUyuI1RzIkTkAK5eaL0wcVwWAR4PutR27q1oQJ+1p+O+iGiiVK+QZLqD
D6wbB2jXBwf7+uxT550sS9uKkeMup4tVcmlDW2Zj0L9D1622Hh3u+S0sBsu/6KusEcIS8k4V9p8g
H/xiH5xgbhchOXZISAr4l+7KBxJ1jIikzL88oGP0HmkxeIb9s5eBDtLr/C3K5emFppDGejmhW8Cz
VCuD4l5HUs2hJIw+eYfmy2UVTxUpMpKBERIY1/zYO/h63Rwp1ODiRpKClF0fRPJWmcx2w712Iui4
uvDCSzDiaQ17+3HrvdT5isupx1TwOITBQUXX/DK1qAmqs6WskOQPsQ97XvPbzEEE4aPHrGGeOyv9
nR1THYNNf+5unTlcafDs/3qD7beS/w92ThH3DdSrbW/kNuDlcyw3Id3Nn1ijRQ1L9VkcRHvfrGb1
C3LLGaiArjMvQgBHNNaJk8h8zETC5PIcnbhRvVyy7SriwVPNY8N9ziRMIg4fHrG7qiUzCNDbPUp1
rzqJAdw6XyLxVfTxmFqjafV40iYBi9cTVPf61CE4eVQo7WooZGn7+qSORrQK9EoKnRSlgTiBQSL0
abfTtUGQSn5i9vWxG1XABDBmyWbGwRw3kjFVkqumG1GDF+RhNOOVnNvco0AIlQlE1npTxshUj0WJ
UCJAx0k00t01TzcS5IGqW0HA+Q5YuorarV17ZVQl18glOOw0jUpflv/ZUgVmo8mq+v0RIhlTeslF
B2566fa+ak/z+UtYZ44agHlRJe+awDJJilgSgdePAyxp/iLm8Bc4rr2icK90WRghVIjYYLC8qv5S
Km1rbGqLExhEbFI93LHdvP8Gz/Om8YmEI79pSHbdw4Vrk5f2Z/asinPNse+/ds6zCKa6Yc3ghiza
SDPJr5WrAB179deB5X5ZgP8tn7JgCnu68tfoso4cyf0E79boWrkUg7MIxeOYCuYccDn7l7SSg7XQ
QbAUomVWUmsr1Rc3AXxTc23pfy9WazMyFuG9YlMtXFNlXOTHOSLbuTtWX9ha6pXszqBQmjZmevk2
2o8L+26lENVzVMypYuU8N2Clwm5GBd7JOiIuk9iXTAiCf8tO3urO0bsxlVWPZN1iq9rqwzYAUIIL
cLbX9KYYn4rRepcna0U2XEALqXosiuSLP8AvPLRB3fRdETBBa5RsLypqLaaaTfJisQfDZ9OXKWy8
tkFt+rDeLGpwpO2mCy+teTD8MnITW9uOYXPreFJUPz0V45wIx3ZSTK8hAgDghdDlk+d9jjEGQTYw
mn+YXymCPoX6R9E4THkqBVpfuD9I3h/YSMd1oWbEnRpSmC4p9rDi3hRDTIIsLjpn6FLGaRcyn9xS
Dk1tlFMdoTS+ZA8ezIFStcy4OCwkJYRr4ri8v/96SmcS4QyKegav7WNHmlJ5v45k9wDUYW84JuNL
caMWmjKJ/NIXlnUSqF+P7O0+kurWq60qoLhTw0r190B6kDBoR41ceFia6bY3j3ooeVzK9lUuzF10
/PpZqKWbv+lWYP+6gsDcyliNDUvliUMKBRui+3CchUUuR8+Z6GOYhisuE46bEee+A6VWtiEx88uq
aDKp1Aozqna68IlSe0IbxHQ87gr+ZXUkYHj91HNM2GBsE7mbDR5wkW9JDDYNAfyx+8EjzSwakWjr
WKtAWV2QLUOvnxWCHV8fvzuLXadVVjDyn/9056qAI7gvQH6vV0kbkBV3MJM0mQAiuSWD4L9wq0JF
aKsMgIyTChEfwwGGt+Npw2rTFJ7thx+zmpXWR/mwvYIF4CJT9PB+SWDj+Zzy2XapjwhEVTINy7Sq
rUvW4bXX6PSLmH4DAK/pxsTOog9Xis3FDDH866CphxX1z+d+Ik8R2kzqVm2gYTWpAruqjTeFtsmT
yLgn6OB51egFQ/pvgNvMG2uWvUp2zJQLqgGEQMbcCwI7ZZekD0YOYbZIRvHFTsghktgXlbp0hwy5
EB4wshVHUWxd9um2LYzbiW+Bp1Qqkdi0JHEEd7XUr/ckdb6k92WxRUS8Wx8R/azegLKK2ph7F/tK
A0sq4fb+TSGLtsix/wpg57bjIX7TX2lnpfSiQ/AUtWuSFVpuMdavFov11KcAT/ESwKuzn9zlesxY
UMSS7VJ5MYKw9yfiJikYMMLkCrwK5ADSpUnWFzcIvJesI49SMVH6xt+bRSe5Qe9hKSD4WJUHEIx8
kR8wxqoXcNgf4j6KkbQaVwSseaOVbc9BNRvboDJRZY5xj7AQmT7CeWKuYFPHIRRVI+c4SKhpKau+
2fQOOn2JbMNl1rWV3cUdvVjmIlBZSaS9sbb3BVpsk+wMaAwQ/yAiNNzQcOFwH33fG3POI2VFuQqg
bfKZ9veaHtpox3ek9ZPszGJJu8RzDcr+Zt8INLkvBMtWKkeBmgzJKaj4eqQ3XqfsTLoJ0vJLjYFS
fOXMvP6IhVFzsRnFsxq7ZP37UpOlexnfQxPyhPePPNtmCqHzMI9YVh3aKPNlkRYR1HvDYMgh4yFI
NWkOkQbYuu6S0c8nfScINtShT+upn29ypV6+dDcmnMaQbzgwVkInaCI/9NGHn/YqVo0ZuweTc8hH
6efrxcDPTuM5JfyjPUZTdjPj+s2fNaRLT5Svp6W2xQmwnWdEDdZYoizVYunp5RsAt7MaIdkmHGMu
VhPi2dhcFqsXj3z4L9hlUCj2mHrbN1v/luBm/hRjl9fehj+THadRQtMXan/x//EtgqUvnfGTfhD6
GOR0ymyyYGqMeYRFw8eZlosyOPDc8qbq6GrHwGv/LJgN0wAnWoeFy51MmdHRcsQifiKPp30nv/GF
KV6nPtiN+QE+0wDvD/eeJFqwFdU91UCxm/VJFgSN45jMBTlKkuzEnfgY8MfLqQtFERdrrVBWu1I9
95YUw78g/rINH32IyAp5q/cJUmYmV8mWZnRkUkn5A9gvUXyjPE44mvqV5gqRGrDfGNDbNqOcIOuv
OEiqYpgF3SrZG6OqqrFP+a6xDD9EzzduDk5vlELCrmhPUOIiL98oD+yQu1iQceV9O7vkyb21Fj+A
Q9/wx/2xpI7obpQfage38MqDELV3IH2UIZBK0ZbKGe9dG+RGjczfjyUefeJLyeZZe+SdyOotjK1l
kMRCfGbIAchI43MD0H8PULut7aV4gEesyz5cssWlmLJz+fAAR5EqKIkdEqYvi0vkt5d+K0W7KKmT
J24ROxkK6QNtpxvyOxFqP279YnSaDlHVIjEILCwG1sh4vK/Dh6AOAZI/XDjaLZSZ5wtgf5WTe08f
N98rnaNwPY7udIp1mrr6gHEz9Ig55c+jTuROho+xZwhhYNtjfiEaTRZKJZLEAL7vZaWKfszjTZnP
lO8L/MpTqsj0TysQTh+Q45ch31fBc/BqYCKFXAVONCfq4T/PtESEz/8B1//aqWzeToZbcbhBL5K5
Gi8GYrw95nq2OSr/SKUFKC4C0U0S4DmgicIdGWrDBEkv5mmnMPmnBygijZ0Kwo70U0xKn0MAJ7Ik
Z4bKBXd9Jvk2uNU729axVxe56W5DsIPr9XTRS5btzg1/6h9hiMnzoW/9CyDGfUsEHAAjEbJf9j2e
cBqd0Lv8BS/wKaS8hMYtoCxnlO3yq+SrWOtAUOnT425sYmDsncX2PTMNcMpnqMxWLH8eopeUnlx5
NSmTyL0Cl441GUnQ2t6ZmIN2Ap6PpRR09M9kKanxuh0XCk24VjVex+1JjQ2tXrwK0TbYxzhQbxM4
ZUzOQKtF8I9Lm83BxlX7sfp7Jew9/ENfV4tgn34HJXLPKUrP4V6VP0reW7DFZHrItIAi4Ei1DpJG
KRdRFgT3cimnx7B5babA9VWuJtPxhkwY1BMQ9YW8j+NDL4Rexm9VlgVDU5bzstgp1OH9a0GoqsLY
hAU78t0zQ02ohiS25jXf4VA818sFMNrW2qS6l70IWNvoQQcw+YLtArKaUVnig4g1vjHmo5L8aY/k
/DT/kTPaV4mvracMXn+97Sz3ExyC8UG0mDlznA5r4De/eBvoFnYs3iVtii8X2b4mk6aVyqqTociE
H8MFUXoo14EhzStaCFG08q53bqiK1zgSUlFIRdmFsxsZhUJm+eOPVErGZBGqQBp+rus+lcURnakR
8hrJgcqfCPdT80u9muB0r8CES+TkvMG/vNREO0KJLGoh/x8m1ICYNlgDEPy4a76b0Q6u9bw6xXZZ
yYnDeG4V9pI37F8u/T9gisRgL3VRUE1xB4iWm7W6fmlHKDgGIZYgkccaH8ZuuNIt60Nv5keJb61H
qfHt8B4Na/m6+PW0SEezoAT/Ebb2uk2fBb4a0/7kdkdMZ57MCUYhNm71R9S9HIoW16/8xeM3S53O
EvnQbKUwCviH4jwkNJSaBSE9LQA9lredLO8TrBEPIDmfYdW/UxkoxJzEzz0RiCHE9q5XXcWGRXr8
RMYlKSeaUaQlErNuPs7ypAmC8IQtF4tZLkg/9W/OpP7hRzUu1cCLBw58QrY8YeOT8vXdaoDp3F+7
OfvUE9Dw58rP70hJ6e9dDNMaAfjCin9o414VihRSuqy1wtKBnHlvPNAqrwvuy3ImKsdnI1mduSSL
EUblhr7PZyWY4UZzEzRPYENe4CARHGbdGMBk5E6FZ1qDkAFxgszhkJQN4R4H5nh06ueQokwP2T6C
Xlcp8Ne/u7hAh++aX0BTkM9h1c0qMlfUqte5ueXus1ezeCB03nnM/uYg7FTnVXfxbCqB1nxAqSwZ
ag26LQ+KbIg73kwGR6T2ZAOtgw+CGqicl2xwzLJHrU0nnyL19nQp7c3fPFBc/wfD1C69CZsEno4y
NAB0Nbx+/JWxoxU41NLwzQEMtDMPcymaNg1Hdx2/pNM4Xo3rQPmFG8r+dVcrPIi1RK6bkNHBqA8M
J5/KTwumbE/9aiXrrA7SDRj3Gow4SxTlNf30RtdzK8Hh1IhOVXT3XLizcBUMwbKPPGLwiRS33b5e
eYIAAd3otNO0tThfeu8YhD2kYe0ijGgg9CZMXOIsMOXyEUKG1wxXQjdKelXNlOcujqkPPJyn73pJ
jkG5D/f3J5XEzcqK6BpLIBDtVaYTW+rOk1gSGfqh8yhtAGrOCV/Thl7f3rS14Khdg9pC/4emovTV
UH1PtTGyVeL97ojzkJ8qfnYqbo4ZhPSkl+7QBP+yT60vIAbNprkVfsIb6zYQ/bexL8INMfLkIjew
1KA42N4cnTN/BlLE4hhjnLL8ygza96I70W9s4Co0wXh7OlVpRdoBFrL9fQxPqWIxhjPV/0wgkuFl
J7aFUaxxqyEq8OP+xwvpqd1FDVxnHs5yZUnXXZaBn1ucLCEdmuJFNt2JuP6/TUqjwQJu9lFS/fDZ
38K10ZKiu7TVASAQ7oalxzB2cl6LZCVYtyCeB36aoC5CKM5bNlf7zg7XtxGcYCRG/gNUdTB8ICZS
KK0i8F/LLqtBSI8t/1TfIuxXeL6DnU0h9m7agiqLS1zTmRbWz/jo7l1+bFsW1R05XVc6/TTmyAvy
I2+Evq6vktBrxfvEc1FrsJUry2Ux0dGzgq/GjLhGQ8fzN36EAw22imXlYdvcMDRjTy+WUc9PMXRu
M8+QwGIPDQxHYOfTqW6NyGJpKPmoK5quRc1XdXp1sN4qFGsneQ4hnN6hm3tMVC+IFe3bZDB51J0G
iRHS4Xw5FnDps5gbUW2Yg4TtzfNC263ulqGw1ytZVfWKLRxc3iHjtp1X2GF/uaH49MIZ6sj7falH
7zWb1Zxr4SCKPEcVJEPp0J8zzfJ6iFxO+jXSE/Yz9P/nz2aHUgizXelSURglX9/pWs3r8U8GxqOn
lsKb6Do+T89kL2m5b7rkBRI9KcZhrsag+Guz1b/LBzbX7r2aY7EvWZr+N9KfhOI3PGlbWZno8Fgx
ksiI8Y8ox6C+LSXjv2RLiInWtoNZwY+lSUG9uxQNQLkTrIHAN7X4xyhph5o7KgHnRWDUjAk6q6u2
w8+suriFi1j7p8kL7iEn6SMxKfnwyaGjOiXS9FUb9y/YhPjsdZX9TQq1Bj94v6a5zTXztiMVENYf
iF9Xl9X4hoTbKN8Daee8ngNCKcy04OZbtGGcWecuG6vuQMRt3oBVtLxfHEI2AKO4uFLXWb2ExhHb
4/mIsHmP0MEsdgP0EUOaENLCY/HiDSTJAJTEq4Uc8otDuo74xk1Iac6ow1FpcpQcH1ihcgUmHemJ
nQxGCKgM5OL5q3nnb+dR8+pt4hLssbxqfmh6YP/FIWPMgO2kDFJRrzOhuAtnhBLLwIR8iTtkm+oF
UBbKLDfuifFx668i6boPi0oSR9A7qBMxVBHhdY52fwmswi0lTjlzdvYmlVSEl9L6xJLA++Ddi1Eg
oV73ogne6Z6bvO5HvU0hRVrCnY/jrRQIHlfaA42BuRpARd2UIOsUH3thL6/7f2+gS7FcIx+VBE3S
lfDhLonmdLzrXM48IOcp+7wyexrfUuMoDrh6J9eKS2klM3X32kLda+QP2N0YYs1M4a2h+kIk4I8K
k8TCAABmJb2geZC4KDKhtFF/bseVCvmO1r6bx7ZlwkN/VDFQQXl5ov6ZqFwFeLahDGAH+e9xqQad
IY6hoZZH4UUD4u8I1e/RsBocoFcmr8A5QWVS9b5LSZieKxd1T0JZJQwbwvmzIyFoCmlS1CetRs6G
ET/4WC/8IE5Q0LQ+ula57NM3HK+U4k8aRZoAjEjYBM5gELFIwWlIPX/048lMSFPGdeUeokSjV+mO
Z9JukGo2FZa1euKzCrPVFKP1c0GpBLOlsjQwadkjKnRnSgl1+0Wk8yr4GGdezvq8izkD2X1Ri2bg
dOKclPKEtX29jhTWTsP5uv2zYgQs0ZOtjUHS9mkmVcvFRZxzIcC3T+B/x/lj5S7M5qHI/79cawox
hRYj4YZLSncqe4Nu3xZzzVqZsBpkNoiiqSdEG7mfRU6IzcgeesfKIcLHa/XLbKTX6Oh/JBz8ESw5
WnQtVhjzlUSFU/DCN132Q40VFaNnEQzdKHmcmfl92q2ShS2BWlo1cz1fKFy3Ngc8ukYqALx2pmI4
iCqlUSb4Aw2xZAzXr1TS71sLzf5PNXh8amWw0ROUMgXKTYfmZH4luZPQdHn80RJG1vzKDvvxqduZ
LDaIFrtn1iuST37UIAcuPqJSLOM+BMfpdjQT+0bi1ttitjIH1Q0pmb8vyIiuyAK87I9BDduAAsZA
W2dMSIFTbLh5/ivsENDphftaVHnEs/IsROSxN+qlKVf+o23n43X2pXR13uMjVXoGrzDTAZJHhwCn
U4y2rEjf4whaRymeSAiD8nN5tdMNYI8RRYXUptMyt/vJTQ4GR9KgSct4KbeUwyj6ErmbTuXX9MdO
1GXWux4I+lrL59it+ipgCtozWjwf960I6Ah8RjStL24HXwdsPbjwfYhMj5u8t4CeT1QrPCsDwgZv
FXMm8JjfqrCXGjdRehfgWuqEPSN5WMlwAQbHrVKjTk9VvPVGoq0jbf3k9/LmKIAZPlwZrCN24k6C
Y9Db+vUj0GGg1pxrrm3f2ZCLHWhrSJGxRHHYv2/x04itmw2FqwtWWZrGGqhS+2DwIiN9e55crht3
Fxls9jwGfZUapnPPWeUBoXNSzqhZMkJfw1Mt2D7Ut6RNejgYmk1xrB8G+lsVhPfo0rQTAg1X3hOq
jHy6JCqVuKdaPCCAo3VRLoXj1fWzHL8xDzP0YUX4XvFMGPhYaVl6yrlVJ7/0gPmukkHOmbN4IMlV
I6SMTyrhKAAvOQ9C0mDiWg+rQig5QYAtc2d21YL7ZzZpv3DZeXzGFiffIFZpQheevanMTwgLLBzW
vqvHNH01WE7lykbfGUvsNvXcafFsz9sxdbatH+Wi9yLp4rXeF/4SKhEajEigjRZ8BSh3nsr+JywI
4B3a6UC+Z5njyKc8lat1QBGyiJYXvZIxmJAhexQx+l78C3A/72KuEzRiadaPZJlW3f5k2HX21o/P
NS0PbBrQDhwEusHy48cu2zA4s/IZdrtSrVUi6+ErJsiE1hrsaZj5CGhNXlbSah5LO5NIVP/IWyJG
JGrRrWJuA/LKsm35xgAInvgDIccC4uvDDva2S3Z93tGZagTgtg0AWKKAzvkhyAcQ8BcghHwKsOcu
Vl4Wrd85SFLZ4UKbEEMtOt3yTPEvIXe+tVG9ue+5TDEcNzD6aYsfXOFswDCXL1sprqmqbaVvm9A5
PReUiBJaXCBURZkoHiRhOx6lmBFd9D11ZkZLj9og8pd9yPH0coFU26PiF5+S4l7F1S2RT8sWYcB+
1PFs/uicF45frPsTxbFIjXFBfaPbbinLI7D2Z2AU6dV2H9VMnDznsMnTd0Z+g1f026uiFyAc/Ycc
VwWZqJ47FcfdAYtsM4iW0wx7EK/4nW36GnygG2qaXzNkY4i7eGDrBIP7+iiOjWi9J2o+us8m798y
ES767zHjxPpD30YdquBMZrzA0Ip0NlWpw1q+mpT1vqZXvJ+PHCwYQ6vIA2cve9w4l7ZggKtn8VTc
7f+sHGuQEU7Pur8sUJdN1No6ZDoiZCoWr59BPIk4L1PCHMvsIu/xtn16jBNKtvtPj+9gxuY1epSC
lyP4l5OnYJCJwAb476rd8Dgk4f3HxLCYqlWnFoXe7h/m+In+S1GQ06UAgeuQBPqpfU00Tjny10GU
jxeI6CQNdMUcDxEOyo/jFsMzKECLUWT+9uQ1NqVwdXEIp7twYtUbmhFAf3lcU+EtkxppvQ+IkSTg
DMbxXe6bvkBI5KcS/BPPYZFiFIWY7UnHbMbsxC/FPmzvM7lWbKCHiDxYIM82Dff/eJiqxRFb+yFY
1fv8Pj2yGUoj+bBhiHPNAvztAEdIfOmTnVuT0JF2JqxBwaiZqn7Pn85C2lfaQGdt4LdovqK3F8Cv
x2VE/yNNUJorUrZj5CEzZqi/vOJ7h1Zj721OD//jT/borqETXIPcoWjieNSEBd9xTES+63+anSUh
LlNJlvUB2atZ0jCpin6QU59DeMJkxgFDHTIYKlJvfbv8bJSCpQ/J9y0gtbK+nUssbSaOMni8bW3O
kcqqZig/8VzeyyrbWqaU0MUzCV5QcRuoZ5/YVGtpatXbz6JQh8D6ouxXM5qS5pQ0P+wgBsfv8v5y
Kg2r0ui/c7KCLsgXLSTO+oaR2UGIzMbFhyJbO1n2ltEu4thStsZ597Ud4/B3PBiD8toVDBRyT6fb
78YnhVNucSn8Nr3olfF1leJ3/UGpKsrzN0DZJy8NBfdlKd3K5ZYXqZM72IGBYyQssEI8mU3UOY5i
MWE1nIGmvcK7QD6MPHXXTmDqAYN1HTzSSu9jnpoVPn4d6S4AUq1DdUKDAUZ/qC9GXdlnq5FnTc30
3ktY7mw4ZPIhGqzjLTAkMJzoT7qPltMNghviQeoV4q0em0kKMIdOgeKTpeilmAQzIXuV8ik7KdJ/
T2Vlf81DgBO7JMMtY+4VYm9eZlLp2sSkuLujIhre9sdQjYRICNV1FbhCjFDbSDLe3xbfQGiwK8y9
UGSOgrBUMFuC4i0lNUBwC+IMgEtB4+oUdmaMTebP8onKdikqJLLU9blPrGLS33GBGb2xvEysgGcj
5hNOje8hzdHHfX/7fA3n332+NLMXrvbcQ/g/kG0bb2pitpjun14ZdHera6G7w4+Ut5wMfrtbaJUh
Ht6MiHwIkeMzUps0wxBQ3hIAoxQik9Y6WpHwBPTTzgmial94k/Nw2wE0RSyO7D1Sh2iTjFV0hZXD
P7ExXI4wN5b6uCj4Hnxkjuc7h567wPG02ZFHsVah7AhhskYBPDKS4SR6v10wUph6YEWtsFM0LW9G
xxCbUsk3y5RWmgIOvOlmZtuRQcJDLHxy9QItBE9iQTon1ep3bERq/AlV94YggwYlaERZFrTlg8Mw
Hdvlo2Rqy8LyF/JTT5cHpY8TxCJ/7bG09yUURP01ezjzWuD+RTiSAC4i4dLllvN+K5Qx2F0/QLOV
IlFuTQd0XPxb1r8b3noEiF88nTT4q+qF97Mx+ypMILfXh/+9n9DW7vRFs5hcZdCQJ1+25hIt2ptv
LaRIWbNcp6UT20Ri/DvjXfx4iTFUXQH9RuckX3UaK0y7E3kvmNDbrRi2IIGbYQ6BszL/2HaU+xPS
oX1kiAq9JAWEsQX2BvOqGdd8QB2o3LAE/Fm2wg08PyYlDIyZkQDhPuunNLHj9DeHWVWBgN/0rfl2
mFf3Bcyks0RRWNDEFswwzO2xhgEHFGbvtPzJu4cIeKjtM/GwhiwWulvCMyXQ+75hc9joACT6sWP4
+1gEkVj3Lfw/fbe0exn+d+Z1eC8zhmBO8GnJQ9dsDVpa68O+tCSPiT+Dtp+m46LeJo+5mTXicq1I
+K3hiB8t0g5EFTeboaD1JChKuyT4w98IVK6oLmBOVZRFSxSnUdfNTkh0hdUyrTAS+oWmW5evcNCO
5gyjOuJNtecISvPGgxLS7ozebpD91aYb4SfePkCW0011w6NLgZCBlHHxiwfru7CwSOXUeTUJ76yM
rtTEWdNwG3bnvAHV9djdCSnrsd1dJXuI6NVQIGNecUsVTHIZVydMYff6A29XgBQkAhWsuzKuDzUY
PdNB9GTeSicEtfxVPFDvUCD6jYrBKuThOCWwl//3SOJIMIVg4OcJJ4vBp+j2bcAmFUM4hjgQ7WVE
Ia0pJ7aJmQEHgrBNdUEeGe4RwNQqOcZbPSRMH9spezqqQoSgTGdbHAzmnhaaAfqE4ibOsdmWA4a8
pmmH9OtyNCnp7THdEzClxkPSqEg+eQIBcYUb+yf9jRSksQ7mjpbKE3Nu2HCQDOgX+9HP42y0aZKs
SKTCwUBTGwI0rL0Rr23Av9IenJW0rCA8v3M2YGsxEvNFeCrP2nBon4RD3Ftkq6i4En/Gi6t/jDW4
CKK6ppG4s83sgw0+1FWub6qGENB+kow4jLanxDuu04yJb9CA2JsNfYPY5YR+MFoX/YneYRDKrWVS
3fiTZNDWQ+wR4NyfVEDXMAcdktbLim/xDX5OOW9Oo+AbevUv+rh83ljFVohkDN+JuVrI3UujaRAs
cNzJB4wAXLcUfzWQIc6n57iR7pRJzrZ9XMIWpyjf9gAyNWCgMcwloMJRWyWqRRZ9l5sLTe7SeVFA
5918sjly/vs2nwLw6mz09551UFc26abo1st70Ag82XlswMEoXe94w5vBLcav703kT9fuRpiDGp+J
1Aw+pKJlQ0cSpRWd6JRLOdSuuqlAUK7AgCzd0crVZ3SoznE/68VT4wwXOSmdeawGNdo3Uuv8KU1U
NVRHj4FPpA3gEecHgBDYo1qNT0UvA8GVZrN9/a9o4G/SsupBeYw3QXOBI6F+efzb3Iz2EkShRlOv
Os8URB5SzFMtE3Bdty20eEOuOGgG9ledufUTWMe69kk/XADJP7MAoBevLUrazxzM4dMHRvAoZ7x/
ka3cKVppTpSl7DXwTfL648qP9XP7eGIAx8HoRZ1UqKphqpfTqGd7KeholqM7EktcgJiAY7CDKDUa
w61sZG4bxhwbsWbYpjJBa2ETek5W1NscfWyGZqx/75vFV/Xetjii1AYN888hwCnz0MroBjzOCWSr
4FMpNu1nExJszcq+CV6ilHrFs7SXAaGt6zlpGDDoo/BNA0Gs3YFT1FJWW5KREWSR7R2EEbrIO5pu
+Z3Xq/TaWVr7GF6Fm+fasDqA0v9fifzByLZStako1QJzie89uIhvkuIagniFcBdruaVEIGUX4tli
lioo+8S9IkOnYvMupB7OpbGjrILz3IclcfUxzu3bJcWCbzdH3HVV4iTKX6+AtE6/qhdK5SLc3+P9
wWZAlLnJsOh2fTHwuJWmxWcq71iZ7AZVZgBAmKQxSMI5yMo3JWMXnfrPKItPk1dq54RUWYC1JE2S
mTnsWfkuNRJpOtH/O0PQnCpuBQnA0KUlBnFrxFTAOh9XHSkGVUxwo4Kf7qM1KXZD+eSgCPJ0pTct
MuqLE1eTbu7fNTkn6TZA0AbRC7HlrUImXiZvFv0+cJe0lG/BJlPXjeZk2+uegALMsdQj1jpndEQP
dQsGeXesNzC+6YhTavuAwlB9m4spa2BMNjKb5PzbvxzOAGiY6+YvEAPFbXaBeOW/L3o5WL4ONxYH
dBy4khs2kyIPWzPbDtBLkfRiqTpYngZRbhe53c8LTJJpsZKSlHB2FbOws0XDSDYjbwb7pttWY1wC
raj1v86TtLVr8NWqm3bWqtUdRrWGTkmrQ+Jp09xduKaCZ3Ds+38lbvJuWKJzkz5Z34sxG1tFl7CP
j/7t82xkYTLn6R0OlDX8n+IWAVaL/rbbBxjMqHUliLkK/kkcqN8WlMlJRV6nLxdB5/npt9gEFTLU
kH63OFWqt3HQi0d7J0Kst+TJvRusrav4U+Ax5jGz0N4w15kA1Asfg1az78Obnr64I0r8/AYRO1Qr
AzaQmGq3w6xgLilIoTpbkZ4aEHBdoiIfJvTewDhvnW3IIKjoTfqiwDEV02Q3fC1ZJb4B2s9HKiz/
NIqJctcwVWtp85h+KardijREezMOBlgXYv8zoni8bMJRZkn1ZYhLrXu8TDY1UtfWxmsCf+bTFwIC
+yDTtC2SWhc0bDi/tCXNCC8LItUQ1GZ9I30xDNVRNpf6ch+24i0wMBhN+BIDAUzOZuQC7NyX4a6k
Ywh2TisnbfFUeLF3wyoHiRx4vYm1wFV1osqEfOIrLgKuqVHUb18/RNMvnP/efKYkxa2bY1ktj2Ql
6RGQj7fdE6k7Bi6JzwzPA1PvzLReM2GHxcGuirvbJtk7AIU/q1SfJdlzmZdiIC+rVKgZ9Ggk2XSP
5HOb2UQpBbVuDw27FocjDMqcjJw423OeQYlQD3rBJXCsaN/4v6+37Wkc9TDkM0Io3hkG16/TZJjM
rtVr3c83ncW6eL0uqJhHTFYul4DjzweoO/IPiO2nM7vLrdVayKTecCmM8Lgt+inyF8v/QCbCUe1H
3Y+M+OEVvRgG+/XqxhGZHr1RnmbOw2sgCBmA+MsI1Ydt4nQOPsUmn7rb+U4DFdyFGJvmLfBofSBe
jdfQ6ELUnpOlUQl1Wl596bEKM5+oPJw0yAubfn32HDvmx5hgM67N420H4BSV3rcB1C0D2N7pLcOx
4pnBZSOHYGi4pRZaJoQxfsK0vb7sDwx09v3e3mRHYJqS2sWSnoaixB0oHeGsMjJwCM2mlGp4t9Y8
tUd30rfDezQBkT6LBxQMrlw/ogH5KUHht5QUsnCKi5K8hvYc9aQKGk0ZKe+6TwgE/iqSIJVrTEqK
cqedNPKrN4vl7QpbYa0bMoMRZmE4m/Lg1oAyoDR+zH9aOHsuff/dghvmHutcVEMqxJRWyQ5ZJDFB
dZctuTdUx86pv7mIOX2txSz4wqyZPbhZ2uVYFN7A+1LkcYYrKi1Mdsb1+Jmk0ehsY6tTlJwq5L5/
I3Cg2vQ6J14q1SmeKNL//IrqOm8nGdi50xdO+H4CccQz5B+pzhXvUgZ8cYVwFkgkcFMbmEOt2fG+
cWDO6IQsQZzCf3lamP7fqE0PEDgsfDOTWbFrOyddvku4DH1e2AFc7LzjsMqEVFofpobkwolaDm+C
iPfSN50GAbm+OajQafNSm1VcJPCjOV1Dil9AmLp8yRCgVBMaV/wFStBfM/3sC0/64HduRx57Q7uQ
PKyrf+mx1eOeGDR/f0h634J3SBlGTm0GQmLIUNaOsdZU8Z3UU4X9hPYUVFgutLdgwWvOOGy+c6VR
haI25z2Um7aNGJFiACYtoa3Y38XPqsn7KXUF/kbeKWRjB1Cgido+KdQ0Pw/QZsY3h5KJNgdsStXU
rBAc2v5b5999u5yQey4uvKEEVmBir1Jy7HrM7UDmsxm6o9sAIWpnOCmcmg8FSpSfueKqAlmN0hgZ
iyA/uO8xipX55x3eCMjYeCtKEKVFBYYBKnOusQOb4HPFRZi19l0jCjCvOX+DNessHqrTyuc12xnc
mF1WuN1uMWnriiZAurnheyhhhk9fofr98AiXyVDiCpzTRiYdJoD0u96DoQKWQRP2zSPI+pMrGO+E
6V/g9n6/6ZEva+XmZJWXNFhEcBXCgNsGSUm3oA6wuFYmnUgsQr0SOBLH+68VET2AXB2eEyh1OEcZ
HXD77b4ngMll/TAn63ceJj4gpt63jTtgrU5s/H0eAngEZyvYEcAgeTwJejqNFp9hWVc0ByMSIz6+
hKw4ReJiEbmHkMZqMhqptXmBOnJ/VU+fm3ZDohQESK1HXWBCxiyyf2DE1kZE9BhZFZtAahK/gRQ/
NaJiQyAl2DZD4MQVZNLm4BJwKMV2KwpHQaE9Rf2KLI3GgrHiAXOpdF573fkLcaBfUsGWV5PP+dkm
70+XK2auKE2ntPs60qLfkdBgkydiy+yQrgHzTgy8wE0T8uxHP+2kcGwMrSBGKYGgL3i5eaC8lk1r
t0ZLmf2gaCFlmcnxn1o0UJlxiA/pstbOQipbJpmCSvw4ma/8qWTGEpPWGkgBDVX0OMZw7WtTpPHh
gdCm1ANu4PFjm7MLC8SgmI2JyC4vuFy64sHTUt9iogKCZYhrwsRV+Ilus00KopBvRZdb55KbR8/5
lHZIzLlSiwKzMERc2+tJw6h8OIe4Pwfr3Qlg1qNrutapItuidmqI76d+CKVoZeLvHszYj4KWPv1f
WATv6pNpsXKXKQ5N1l8m7PDRn1yY8K4pyOhofO+AERsQf/D8uX52d7c0UxkgP10NMrNiCXP4ZttI
y8RwyZM3kiOdVOtZm1292+pDIor/3bstiZ7nkpYsoKHOvIwAj35bHze9viDzC/6yUGML5KuzP7MV
QrwRrPUDu0qC1jk38WlrT2i/TUcN+CuvwptnQbVwHphcxTgobDaiKtH7QKCHprJW5OGWMjjvDOWh
vObdxnc/cD3wCNAhllkL9DdtNetjq7w4cGvJWxvhFHTvCfX5uLaUVYJFW7pRaX3sKm75G8tpyPuT
LVV1a2i7Cd19XI066uEqmXEXilQZGzgqFlhzNYAowKX6WmXggRgk9sIpyeQ/+Df6eIztf13rT5i9
WtyCFN+rIc0Hb1kPVSumz0AVDA9KfUy/EpX67zZ4WwMVit/HU6LXTCKnXumZZqfz8wU56eDBRNeX
cic9Fd+Dbg01sG4o3Z4MWvTYJIcq7sqSuTAK31CtCpE/g2YvvxtuKLiKTrIhpCxcFyEPuLuzI8RN
FgAyqZZyVLmTy+cd//Q5ztmsQKFvImZ8JuGLJoUOuw4XC/ptBl4REOPI0n4+aXU5eP2+V5pyOVti
3OyuhbP7s3N+IJFUhsjDzdWkNNS6NMCmW4EdHPzx/FNhkXcC3wa0jjzAUnOWGnnyZBdqRiVkY8no
ZkQ5wG/3V6k6jWPcVYdCP9amxo887YW7tOVQoNrJVbJuUeUWuPQgk6iMOAYMtQ8A8W+tfG/7Fmos
VOph9i8l0bXaVALRWccyYQifqjtO0yGdoyJRoFDHciZOgRD1Gb962q3fiGhncui6S0h8GTqwmN9E
UwFTYvry7oJZ305y5Z/5dYSIwnw8yoSAfP02dRs15QvP0zJtMIOxA6zW5MV9GN1lpM7QmXmdvQuM
pV1CbaGwU4/y8gH95/R0UKIUC6LJ4ZzGPfaDOX+cRNaAnP7H6VeYt2TZxhzIrBrsqs1fe355z6q8
sF7Xt+bp7jIVxi9TL5qi8GDs/6VhtTiOQEDVzDT1u0g6uG4uY0QdBRu9TNdVfTwSx9l41tjse8y2
OO4OGL2wooUjOpJ4fJfzirh3h5pylgTSksBlBPWIjNczjE1LP7YM9d5c9ObWkGNyiNx8t37FE/vg
fC7GDNoYcc/ahvHRPYLfTs4o3D/G9SUHXb9ZS9/CD51n5w8seyw6OH0ubt9npcQAM3txiWf0n+dY
WwByavsG5YiZKaqYlr5RfpVp3R0ClfOiJ//kgNQ44Xhn/XyNC5mnjURUUWxPc3vwOT2n0X4qNKTJ
CwtNVG5kIe9EtSu2ODzoUGkj6xuOpEsri4ojAJvQR9seYOegwOzSVVEf5HKyTM3d8c8QbxwSzJlT
GABj22939C4c+HXlUvDW4+sti8FvOGcv9ymz07ZGKAPDxlskeHWWtTY5MS/L5GNeYxLIMd2GB4J9
T3RyhNWEi55wSkNCvvDgjB9AI5pyuO0RESSNvZLpJryWM47J1c47MP64UspcpINDy1qN/1ETKB18
m2GzEnTjY+s5Z91Mc/a8umKcjlePbnl29R2XtQ6TXF+TWhW4X2Qw8IwiPZA7g6PrcNPccoAfVuFd
QCu0p155LLhoRrUKmWARHy+no/04ibQgcO6RJz3iwdRDzkYSBxHN0dJLzYc4fa9eH71IxUv3LDn/
GOWHUn+xnHRjLluMu6t7Zq5BB9shQqtPsGwfrdwqM8cwEHZl1+sA+3g3JVkExKX7/hy4MD/32KcN
PNUax9LS3aTEZ9iVcN2F61E6mVfesaEA0Xydzb9gPZYGcgvrB9u58CPcEf/Zzb8QigxpW1ZO1WV+
czLJjiwFAKhRUILGcFA5hJxCcSe756RJD6hkzoK3sOGG571KMWmnMrrNaSDRo8JhJ2aZNzBVHAVX
QptIzjAAVH0aFKIiDu9uL8SMwMVHiMbrBfIkT/1TrAI/6cqV7jyi1nZ65VsyZUuwa4NAny/1LEpd
eLU25l0qKAv5wVhTzBAJG+dDxmNUidjbMGACEnsDaeg7jEr3tiyyua6Cr9xbmwLDwliIyhIQa20g
0SU+xy4Uzq0z23h8e0ABEAwvg7+GlwN7ZZdW4jo2WcVo0E1WajpyXCiNHT9t+9OsM0kqs/p3PmQv
2mRtFioh6qhNJTRqR/SVOeTCcgWShpkpYDl4UzrKq3FS65BRBtpEikeAFyFQJZDrkCjDljZhpqf8
ybFDQEfpH3+S36vok1SgjISaSbstwzQc6ljsS8L6f0yua8CzW7FgvdQW8sy2QZB8yGFHX6W/7K4Y
FV+faaU+bV1MTyciHRZmaskB7JXbYaCROcHs/56fdqyPK4U4zul1mnOeptWPAk4d9oYNQWnaMTCm
x3daDBUNU5j53omWarBcIjkPpRPloFLTW9YJBn7CPmGVRgjg0OndOfq+V0mH8FTvt6xerNDn3LYv
rF7SOcZMdtcykD6jfl24TOwfApWjGQ6teBmqjOwifQU8VTKND1HA8cgWRLaK7EHowhihN1brA8ZF
hk2Arqy0LFtsoziFWrfUbAKwOZetVxFmFyecaLxjWqCABdBdxZheSJRDk7vRQpoPbPJ+vO/dDT21
EDCV2/jdUoAAygqNnSl32a6R54F3recKxQhKdolb3cRH1BI/Pi5/qFMtZiX8J32JSrEwkwrTpjko
7iOEiJF/DA9LJCXaWs7YWYbzLVJUPgriyvvDv0jWW1q19jOtbiKbRPsBib1dPxAIO4cWFjfGGSjA
GoO7cG9QCcbFCHs1/YBZclOYKLFztMSk8AZqId6J4T4cdtnUyFCTS+orNjME+zB5PkOJtRwUaptZ
4hn/ADBcFCt6QhDA4GDxOzmoDcOxcDV7VUitQyaK19nO48HW+lpVUddwseB6R6NgcgKHh2TLD9s+
hcyccpsYRWZ1UjcfPYa5/wVnreK5UA6vYo8YfGn3DXo8Yr3JcJy7ET+1q5mi6o/78w93nmCNGqZu
haE8AcL0HJsn7LeK0lGQQvnncXVQqg4ZxBT9fAWNg224BownJZvu47WL/hARj9fafIR20d+6n5SA
xl84rQRdBmWt1TddOI68kT/UZBKpNKFwM7rwejHY3HEBr+oF0DWzF9TC4+tAJiyURHbPPazzQHY6
7YCMI058VhrD7ug+JnatuYsRaV8l6LxfuOrMA3a3VJBH2U/Piy7wqdh2rS+4+woprytHmvXRrLp+
CdUR07DoYmYg7zZKUKAYV40uFxAQSJiR8CcXJ2uaD+FSfM4bwjVn0nNENLW4OLrsHyPR94/ACuQp
LRMXx31wqXM5l/4/tZTZMcAU5jnJM9PePSFiAglxl8zbSZgX3NtCs6tjbrWBWmq15/tt6Ii2lzwy
ATJOMYq2SqrEVo3CceIecTwhROrXj/VINivJHC3EfXIQiN0hXcyqQ9GLndZWbV1fmltmTfa4u7GO
Uf4EtKF9w0rEXpQE7DjXC0V4biehdIHnd/8jCAwhxlTMj2SyROUiV03VUznVhzeBdTlv08JyLhdN
Y3Sl+f2P29PBLktNyMUVJuxf9pqllP0TyRa/0Zy44CWWSSlTPv2qpXFb97rPsTRZLurL/RqkKA4B
3x2RqMyZbSPqlNvnbmYw/n21BpVi1mn3lc5c53HAL6YcrJenFoFY3FMQbJQpXfM8J2pbDUSt4fig
m/gkUR0RZbfIp8HCqyNVd6HHI6CYZ+cVjEbKWXQ/FpC4rKb732OJYqliNBMUb76Nyq3lvhOpUP5e
Nki5LN+w/EFvhZM5J6xj/Dp6FLQP3D07zEoGHvLvJfXZ1aFwtfcB1+8O2YQ60uBrEhkd81lQqmRV
naxJzk/48zfxkmk8SAZe+o0TxAffXdq0FuXDdhgML1K6cn1yXf/qvJD9cfE0tuFwtDxdqIUFC+kA
c3up/7I5JV1kd/DJLauKdDwaLvmRRzK3jtnEHu0sKjmp1pXtxnlKcoH5e+Vcz/K8gjqvG42SkznC
ywjrJM8ZzUOrqSpyGjO+rk2bFTomMP2fGhgUIzRMwTUbktKz+XkJ+YJnC2/gtW8psd4kYYZzhKY6
+9Hchec8ZiDgLvWG1ByHiGB+qXHaANtliyqdqmC3eHqlUs3+4jgKsiyE+AQEWlnY6fSL7hZdXVyL
nHx0JT6LzAqXd/WjddWnzi27E2cPN2cwchywH+VDLVqSBDTl9vNhtgH63RNihAVgd2uCuw5e+lk5
8HGCHXiqVc8vHAVii0WEqcEa73rROvBp1T+AiWn7LtZEDQmxo8ojMmeSXhDlDtXUmVv4a1OzWGao
nXRTUgMk+fuYGSBW96Kc8YVfqTDNnn+mZQ0ZpKaPsQmQp039BseTiZoHSSog0o2h7S5YysPTQEsp
o17Y9C5tnpdx9FLm+7Yx9zPiQ387PGursi+15cyfZ2q9CqUlPooIFVZ1SdMlx3hThVDL4E2DQM+/
o+LbvE7fG9M2Ld+QnGJKKQQKHV9rkcc8xcjq2HiZXV3iwvS/k04yMVOMg6GvvyYiIAJZqZIAD7dP
RS4/eLwzQq0ityGAfOMMlm5uzhCwXDYh0bk3Dzc54lrTtoXmMZW3RpdBdMJOTIqOiMF2ryIdTZzt
54aPZWX1okBmrghPM1RZ0AEPCRFYocj9XbPcSlq1b9sI61iIjHDIBEkyxWoXuBP7wJtrv5LjALc3
422Qoy+td/eYcxMao4witgafeiBxn0gr9lBj3aa6b3wfaCc+5FRUZMPydpfvJSOkb8j8r8JPGtrq
7TRlnYsHzY61NZeZgmXH+4ePgutVK7uQISSmm/9bEwEOQFc9bkUWBZcNuLBobbzqilRtI1apijqu
3BGrJ2IxRTgdlhuVyDIB2oYZMRJ8pwhaEzAVz+dSYrbEWmLgl7iEUl1BJwWXLTOQl7LlrUZTelxM
Oj4mCOsX2zQzybFZgkkFPJKnzM29xyPbBW9sxS3yrjJwLv8J3xRAyBct8RYWLqfoHuzsQCuvLi8E
3HctK7JGs0xfD3BSAUtCJw+BCP5RrOJzVWcEd8Ot63W86gBMekj+FwqpPVLfcPzrA8XdSVYLfNL/
gHWyxPHG8xOzLm6k5vlHmsDALzxppJ+TrYhEc3rjrYGzH1VVBHJwOvK/BccRHcZ6xUgKyg1E1lNw
lTd168KWJPtrWW+MmU2qLtv6vgXspmiLpTbBWq9xiTRATKa/CxBq3pQR7JSPyfC/Ktu883dpztlY
I30NWMmJ/P+ThlGl3obS5xXR6vCuA/ADrHQIzqg2AsG6NTUmlufbJ/YUaK4gw/pqTJI6JX6xmATK
K+BfRIpBpR8jJw/93RtZGgItfWdAekjxO4KUTyKESbcNNJ4KfFmrH2bP4YWlLg9kUBXGyXK4/UTS
FWxGUJF+d2lnboOawgj/nYNX9yPXd3DkT0snkBCIRd2VnH1LHFZ97N05V+1HK3NJ/y8yiWIGEm/B
UnXwGK+NBODMnMoN2ikGeLpxBqkN5UKwDlYGDg4v7/oUxNEUeAGT5iTloGbf72jhf/EK18S4uDW6
qxy8OyKtDp4imv0ODGSKrNbn4CfR82tSRL0QFsyJ3Qs5fCUOVP5WKFafxvutc/rJ45iYsBDVXlw8
gpq+dd75Ix2k77vqhiqLnqNJh6mh9bEQ4mT+a0WH6shxs2Y/wfsTn81nJ6GoPbtrMCEUYydwPyo2
19O+eANxEYKfht2vmp33B7dL9kE2g0i2S//4b8KzTQncO0pKr88DqUMoTaMRRyGjXp4xrXTSF2XF
+EgTh05GxRYoUMbEN0Bo9nq26j40bBsnoVdaL1iJe65yDapVbqoPMuPvFwOif6wbvqpVtiok/Ck0
cetW5w36IObYp52h0UHJurgBSsXYlOWZYh/nXT69cpF6A9TEK2USxAd4iuQUnE6/OD0IKxyDzrIE
SsJMDaDdQ2cVRTaB+EiyxN5dqEt6nbjoJFE0N9F1Dygfw9rTt6gHQ4BqFMa5WAZOml/XQRzubMUK
KfkRMGBDMp3NuuhqQ5Y/5C5JY7MlMlcJZpIZ3+5jMt/NVk7EJmHyREJZt0OJEyBga3m8LU3pF7FH
XfGknaWhzyRKVJRvrBKsDP1DbLhTd3QHeB7WYb1oZM5R+ESDYRjkSS6KVukDRzPLnTv57oyVdTOa
oy/xGoAMxr++jqW9Fwg81E4XteB/YldV0i8ZECSuYTgysS9dQqTkbzI6LepjuXsjOUIo7RGhXEHd
2dN2LzgLhRs2nq1YmwM7lMjujWCXIbcnx64Rh5p/IORKfBVFH/yIW1Kj8Rb6pXE7Pq1yI/y4G4cq
niU1Wlr/WK6Arl9bsXwFU26U8VoO876udcTw+afkAmcCb/SnV9MK6i/zgR4nKzA9wpKmSPPD2T4m
cmzs6hdG112kBZpri24agQN9VKH4JjVux5ffYWa0VRzn/Jwc92YFLnIQCURLOWjE6eXgYZw0qVKW
zSuh9tAH4+K3+TbtRxfaPl1lOWHmVQCp2CWHIDs0hDVbaTCJ5SHk61zmEwu3vV+lkF7vGrRS6qpn
H1BkFPm/1OlEgYMy89pom/HcVg576mKHeQJmCED/4xf/b1bQ5PVuXzFcUnRIXC1VsvtBENkoqJVm
N1g5+ZP4YcnT8leJ+g+qHE+WhIWhOYxciXj/pEgJ7ywD8dIZM0L9HddjbAa+N8DKFHEJsIvZComr
EUHRwPhnIDcdB0Ti1bFdp5xzPB+gdmkc8i4+ADFL+1QyOh9gTJdMEoEvemTrOfdrdUkTWiXuRg5f
1+M0XUKdxCcp4LuC2A3Yj351e5k8KIi7p+weyhNYPHW1YuETNbgvFCmz0Cqwnjm3RDhK3mI2FxFw
w0FQlzn0RcXXixS3JHo0ZjSmIeSnVTtvjG6jK/HAEvOMqnnIUVTMDnT1iLsgtk0dy26+jASgKDn6
k9eZ7aUoIelLLUQcXBt72Xrr6FiwQSluECgL+Z5Uxc33+WypwG1hrQvEHKSmJj52enOxty3UtDyI
22z6EphJSUFa6aODgV9l8BkjY44agoDdVU3+TDDzcu4j1ycC+uESI7A7OCbyNJ9trCcs/i5WiHwv
hflWwi81Mbz0eZ9fqOvpdBihXpT5lclTK9KJuKdewtZKi5dz7bwscq43uKWCJeXtykkttg70VQym
uMJv/OuJK/OXIikL/5b4iYSSDo5NfJfN3wASLHRyrpCYAtRfF8WI7UDVo6+wMERDUTyOvLmKzNXB
4dkwbPMjZgmKNHYJxR/Tu7gDQ7O/nxJMc5Rk7ODIHfWsyuOwadjiHX6kgLQWtcVRvXqySLRfTuVb
Blh0/g63dLh+A7rBmZpb4s9h8ie6o8ejot0syH0sfFHtoxsS64rb+ejXpt75peJ4h/ZZPk1mQVp3
jWJj69R9bR14oa2QN97wgj8oTjxv9lF9xMKxlpxBtYR6228GynbFpWUGKcFIVxTiU+/DXWclmhcS
dAjrBJVBRES0TAmFs17pSjf0MjvyY4olT0cMi4gL9DYAh7dNr3gU2KF0P1Csl55QGgB5yWJ12b2D
GXIeooNuWfbi+KSk5dXNQLLSte5eW1hT+tpySJxfrA1sbxkwtx0NlUGvwpHRbVU9mHlfA1rmIJCZ
KP3yArXJydkrBKWHuy9JXnmsclD9ISzqTW3F4icP9kZ3DxvP/NHsEr7fwVqCjz8pgi25v6D3sCa6
MGFdSHCsJBpnQIysw+SUmjP1coTFPfLLdPR3KWVmuG+V4vGq59h4xRiZwFgZeex5e+wCr0UXZJXq
EEOOC/wyK2snEe45ICy9UpnsXgzGf2tq665aTgGQs+iTXKqFOMjsyQyblUKzD+OwjGBpk+pi6Hzf
JGkn+gxF9tk5h2kSGABNia8wnYGwhCJ9Va3tTEM8dO3Tt6zFPoyeoDoiaI/L3G8Muq5ZbmNrJAYH
FIdoCEUPwzTkRi8kf1P3Y8+elw6boNhQdaii2EMdP2jTeegtODW8UFaVHBTeqcd5M+VXZRQVv+rD
AhDWr+Z6Sj1Fkqq+vp1CubKBiDCmzqB1mjvE+KWci6jwZnGdBJF5nWAlpixPPBCRN7BXXAmlVFJj
m9djLOUne7mHfG+AtQaDtrIhmNJ1EFpwMIc8G+7EaaRE7XjLK7sFpJDCodUKzmyppAQHZEAwbOAW
82/yfU2SYyAs/dcE1J07mSARPAiSqAqxKNDp9qW3Yz0fVowyBG8NVx/dc3Z69GiPW1NgbtK1qInr
ZI76jOSximdTwwux5Htai05RRGPQTVfWFJL2PX3kG950JA/zvyfNw/y0gvwuFIAIv/dzdY0LhE40
bEjp4+iZ3KsxCvWKEUQs1lA/jFboKx8fWUUQlHC4RXRMix7iNWKEOEmxfVTTILlXL0QJXr0iamx0
kabogbC7vaA+lCj4QeYvBmMFcp3wC0afUO3i3IGkGNoArKJNMT9LEkHnF2oSSgByAgOQYHlrDTrQ
hZBeZlZuw75dpFWyQhzOv733cIF1iTSoFszokaZV6KkPlJ5/Fr0hx2oZT/yTIETxh3kyufxuPSce
7yaBKhiNLiVmgegrVQq0VR4AhkGGnwRI2BTM33Oo54e5gZyly4oL0crP85t1x9f5MQ/ZJeqCkXXE
LbXhgTInD9hqeq5NmfTowd2OAGJNcgTPYo9FX7ywzA1DVcqmI8p9K3B0F4+7RsDyloBkUt0RHTIR
axB7hS2uX3zaLIyJYHEjeRpUbbiEAWCmy6e/tbJCVOZGefCZSOCQb5SP+H2epHvomnoXvLiGSzPR
wb1f+RiHN0+qHh+3LwPS1zLrxS6dE81om46/RWSCripCXG+k5JqEx8OMQo5c34EXLg1148nnX6f6
31v4+CYNZ7k5e4/IyqptwkBhbq4Ip9HxAWnEsy6Z5//b2BZm7WcTwUmOnN9kuJ+KQaG7I22fzTVA
jbZTCm4f/kpSrGL9Ck2+7k2FVN8xoXSP1DtDOVUfoSybXsP8VUqGlgVvzHSC2+1taxQL1oLgXYXM
vAmd5Qms+Kow32CMuPEQzhdinyh6ZSjQSydxLfyXoUaTrUYNZ17mGA9WeoOY8S5RDeFt/ZFviDyM
l/5/bgqgaaw4iWRpERMHeAx9aGm4KIQbXF/okJA0E46itnUm5bRKb3aRJCN8RiU19LFgMV5+A1OO
c6+obkNy0eGs7fPQIb6Pa7gTM+8x1rHyi6q5ZwdFyGC6KK7KOCFtyTuOiFaZ8fl74EadoGz/HnVo
wtf+yxyuf7XlJ8tw8pi4ncfqHWIVMxgu5Qg6gaIKcQyq5jSbe/5Pe3To5R6xA7KFuZzBAdasM0EY
MaQLqTRyIEa3/3misUdb/JUTmzfYXVTXmq9QWhDuWapBLFcZMcUrGxKi1g04LZDbDaObY7VnBc3Q
XBEysVVax+SD7PicVHQy7nNhZQPNgmhKQaO6CCBa2TtwpOeNaavyMs5bD9YNOdKgfCOghSSXFxBU
JKH1JPDmg3cwNNH0jbFWE5QL7eEapVK4WmdB5Dg+OEVow1LP+UGvIVwbRHQ/6RsjWOJ+/AKYfxfG
hs7/c+xwZNPMtwBcaKVt0jkBwTT0nt2vjiJ6MZfIOrN7MJBCegWQh45N+XnXBkyAd0F2ACUTyZTQ
LVKWKwVNKc10l2dYZ41axlvifZ2qeec+y9Ixb5XfE7OvZkaHNOLq7j+H3ssJI73pgCNJgdEj3w3M
++kn/5cYeGMdYrsmRWg/Vr8wEhkgH8Z/piYHA3OUJHeW/XeIxNJ7ShC6QCElcdcXlrGm3IdLcktI
uJL5X6S5043i84vJRWCcvYTb3WLVMxWWqXc6JNCv7Mzyxn1gMBfbDd8pboBYV8jbYuzk5rK7Tyyf
NdPMOH78pgjXHSVO72kmKzBNHcP/nkTgEgeb68nqjrv6AJWPfGR69yu9p73gdByy9E3oEunvbAmm
YrrSGoW5p4cNa9aXnGeUK5EKCVsFU1Gl8aYwxoIqAKzcKnxLCN+hCCsQKsy6QYhHZy/GVpB+ex3M
629e2fQ/LM7o+vg5JkkC2JCElODVCNFZnxXB7OCB4OY7ta0oGFhZZ56bwpR9fHw5Q++Iyz6hoXXk
ka4XvNoZKhGmtcWHCWez9PRESvEc6h7ZpHEXFX1lpdshnisxzQ1ypPOFKw+Cvp1c7S34Pm9lW3Yn
4yzAOtJLuS4erpEOoR7A1Uc5HA3YjhiguefZBCqArCNynGIJy8rUsIpnfZwCozl6/jLZNEZXn/On
Xop5qpJifBswxrtxv3Cgl+vlui63toNkZikBYWMlo2J7R2eeTdf3d5l2aQ0NUKOdh9u+kNP51Uvl
sRCwk3aWNuC+sI++rDUZUfIF9ossr+oynS4UQqhJpI5o62kekwcw/YSZxamIX2RiHaLjKJZGFTsd
E1XaAKHoyXxLlki0NiUTgEpQN3wunBP7ESNyWaUYhOaKco21xydk/NX/szxmV+lUAzRR5WSM77n2
AaSSLoNzNkdljwkDXzt78ML/OJZAQPlmJgBak69gI3tp3naKYdCGlZe2xsD5qByhF2Hcbex0e3QO
tHCsP2rs3tVdcljuWfVsNlrx9iqNgy3RwiuOZG3YGI3bKBde2AzYZzkFxlfIbVnzirl27EWhY3Vm
QhR7VkXXv+37mQhD6cuAYEB1cFW1aF+GP1bbZAvljD1WgdeTZt6jtsFA8/2M42aY+025jGMlhULG
dRahkXEL2b9/bA4c/lE0BfR8nwNZU0qZITh9+wDAnjwEqP+JDUOyprFwlaWpxJzqH1n8ICDal0+0
tMSLDe9r45VPJIc8QJjKKhpM9w+RBLOtbgtyAFwTmmbjNMGbULTxYytkYCUdmiJscAuRMBtKQISe
l8pP0CdnAU96MpUpfVIIjdazpvuzs+Gvtn92nhzpR0gAHVfU21Ifn8ZXqGGnEwVr7VoEVhXty4EV
H7hsXhKfBzjvasdklLDDDHh28xR7M9Acbv1rZ9UR1HxaLFym9sISSJWlXkPoAwqNDHUPuC4xH+e1
JtIwLdFyxn0BPK+0bW0FFn6ckRZ+CiXIG7efDh8BESYqgU8ND+9I2c4dp/f5KEBed+tIn0sNSCLQ
u6ZoobGtjthmtKyQj0AZAjgk7bCg8GmseLnGgE3JqqrOWSVPfNzeiX92d0J8shi4lOkv8E4z49KW
gNanFhz2QBw7E2Ix3CGzl2qy5vPMNB7H8p2QK1rnq0TjwD+j4iOGLIEUyEyD/6aJB6O0sPFTet/P
bJ6waxBaqhAk5QBBA51CTSbXvUG5Pdhc8Gtm70rw9J0X8yqFiwI6ZZ6bCs72xWjgozy2aFpDanLF
y0sjxsN7tx6zhPFb6VI6PWkZzjKWvzxILEW8YyiSY/R2Kkkokkgzl/nf0MWtagParhFR7pDPXDZr
wOYfL8LtttGu7W4YcPqQ1yGkYuRD6At9IDbPwZ5JjbCCX2GRhezUDt6l00e62cwPZnI1fRMW/5Oa
2RzGfMpC7GktkH2Psj7XkvHadxaV20l7llXgYbKB/ENvu5rrSQ3FpLOQGPka26i5NHQgKqiATopw
p0OhwJw7CfZiYm0uhWntgnSv1A1WdUhAi1MkTqR5AGvgJH6vkKTfATD3gxBQLZGTEtuBauFy9iWB
8rWpy5EUEHRMaHyHL1lBOsn3hzVM71/ESUZRsyVp+jpnWd16TNGDpcD6NsFnPVZ2y5SGtFjplMOy
hTkzPZYxouemiJdJ2W9KzyX+XJlv3o2Xvj0ykTc1wQLwSGRHXBhB8XGFyDIfm7X2AUG7GoTf1wM2
gAGHougNXnRpKYMY680ResubUyQJfy0Z0ucIvdOIByaHkXB7dmCbM/vAuY+9hY0KAPMHqho9aEfc
dc9ITkslZRG9B2jROqsDwcdEJCl/PEq5oNWyOomuenrvR3/BUZnkBS/eBVvARJe2uSZp3vZABnpG
bpG7Cht/bq5FheBUvbFRJMpKtw1uKGppAfbjDRCVmWfdLoNmIY+pe1V77TNdIEDXFXVvh+EbX5lA
Pt2uwH7S0jPHl97z7eMADy5T96pg7qVF6+5ou4eXX5GgGFmTFmhVdrzWJnez75OgmGugXGMijlWx
n3GZOBCNm6f1nW+SOE6WWfqvqT9BE8iRzHqVycNTkIQWDjrY/OnCRztt0zRpiVas74Wj9V0aEGQq
LfBadE709gRHW4TZmtGxALFGH03ezAHV3fxmSXg/rC+kroVJvxfBX+BeB1bynSQS7xDhNOEFirls
nTqUw1OIwGNP1xJist188eGXzL/QDhIijlypT+oXlxrhnTijT1ITDGtzNmDaIVfQ7RSEWWQMCQaB
VSoG65V/BGlQptBE2z1HLJjCEQunf4ok/OuEhv33kPapTjOVVmdvCVrKdcbdjht2ey7j7jNkjD8A
rCz7qvPYnx9aCH7QrL+r/WfqrUZJ6xTFisceXrc3yj5Fpsg0EAGIOgZEsll5v3+YHR3lMNMO1oG4
GDOoRpRZneMbkOD8RT+1s8Us+QkToiWdcas371xL8GDH2thA300nEvPR4cmcmhr8mZMOUaSaejI7
eKRFUbNo0WxrXUtYV6uLJqvOI65kA5Fiatz5gPBRuU5pC8cj/ngiofCBK5pEb+vuGCo8CGtBFL5z
HSeKu0xJOa2PaA5yZUKV0IPVGBP2Us8m5kJpEdSEsrsGxX7IPzs2tpo2xYkWPOXUbJeyR8TvegGU
1v5bZj1LtKNwiKzrG0NfbxqcXEOPBKpbqSVjR2YJmvgNUD1umkdOBAAzBGOhT4rhZB4zRJDK6CnE
lNLJCDUr8QQkQ28ugrY5gUUK0+AFjQMcK1C2PIWwe5b202m8s+lkEF33kEL9XWVQaSS4IWQn6cCX
2yiFW80dl5zzKKWuJ8PkkKavclcCWpzMd3dCPVm9ZNE8S8jJVqkj+SGEbNynIIEcYf60nfp1/sz+
wCzIdf5EJnEk9iFORRYh9vyHx/XhNYBesBM9p0uPlxCElGU5oo/01atKySqs3fIeaD2cnW8mjoz0
tWC+i8wAZ0cFum98q2Nseo1cymp3IBU/xj1IDjQKja1gDRW7vuaMT9Ak3qMsm1MbHWDTi84PJ11W
HA6xmuPemopk02SRBw656VYLyv3ArkLdMjt+pLjHkjAO5uzl0CCDH12o02OdXKTRFWyl655E/mQd
Przle319RySmaeObBksgnmxuqkNYSd6ebECd7JBvJVppVZXmlr/sj2UlF6idcoN9k3AdR+2N0BeS
y8bsp3crEc0IAlghyCKz0HXO9IdJYXW+waBF11fDBdVkPnQySkcFYhUEsjdoDtQXz3rlSEJ4I+WA
VRUeMG1q7kA1uI501khNei9xXpp9Jquc00m6NAOMod8+0Df2LRHSgAvjy9VRVUYczDPuCDBTWAz3
nD+T/TAQLeA6el2TZXp8MhjkFZIgTsNtP/a6P0crktLdpRvKPsJ3XGbCMVAt/W1jFaV1rzc5/NB/
AGif8mnn4y+IsjD9S2ZyiMaI8AAOLtAU8O1Cy7GHVLdy1Ujhh5RtY+YB8DKSgkxtvFh/dMaRyd80
hNsRSGd6/+sqjuWpGKlqylUIlQdyCJioGjrSzqzoUFvHlhQbcwW5oGZubksBV+cJrmG6EtIlLQt9
z3MsjFhk9F/76W90XtD6iHC3TqYATeDDeWGH0bDCB1qYMznHmzvbSVVkUJQ0dgNWR0S2Cjl/lmCH
5GDyIiNUQrfLBC74fK47LdIvUZ8eWLMXEAe0XN8vj2ywc82a7HoEdYQ705ibialcz2PG21nLpyjg
rjyBz2uKxWTz5tBWgGAaEv3qjgHAgLiBqVEJFVK92/sSRuOIeQN8ib1n8SdmFto4ncNtcW1PuJsT
f3HtBn66okh5E/CBwJfkzb2WwA0bzQviI5lBbFFnzBueRuWBwYA0AvU8M+bRv9RvNyhJPztUPM4j
GyEn3ACH/RkZt3/p43ptUt5UqxEEO29tIErQVSnsjKx1FUmxwPHce4Eyv1SxDmyBmD/e/rjd4gHD
J7K9+reuiBNYLxWn/mb0rQD5kUEU0e3BvbksO+zAIUQROqhyFAulEsubwL0n+Qcfc9yD7sGC3892
PDdp96m187o+VbAaiZNKPaMVG0dOvmZMN1r7zdDgdbQKQj3NSnJHjDBFXY+R1gUHaNRd2iZcPg4O
eNriUoHjzrEzsyYgrVv7Rw1cH56mLIhkwazvOUp4N1bhv6fcXkAcWbVjOU3xf0WI4pFr2vBOT5iL
PVnruhfD+HtY99M2rnJEpkDBKaVi99GhJMqAXL+vMNwmBT7ZrmPRG+47/h7H20kEn2uVASEEsXmg
Sd/cVNvym8zSDVQYgdRy/iNYI+76RgacJ6KJT+qXbM5NduV8sEsVr18g0v4apwz/bEJhpliO85Hk
0EN0p98JpaQD82fbXcSYFhfTIsDr4ZHJEXN0kgTYePAO7bHIc1VgplhEGE5pAL7LRPMLn5EcHobd
Qi5fCliol7G2zQC3rJUdwp9RtzFcoKgc1eeOCSNQ4bLT8M6PSgdku4mZrZ3wPj3u3BnWR8Sjg0LO
w4eKvxiQ1HUZ4wP2nnxk1kD7FbLZk2D9A2/Ae8j9+arad6V5rA2pph/7gJxjx3wcFUq4vo7c7y1M
ytUgUAYvodGo4xp9lpbWyJSa1Kd2dYW6ls7QOQpxl3HOY1dcNCZ3lxfprY+4rgWS4KeQlAf0IaU9
x+7LEVgz6cokjpqBMWpqhG4wLsmfUbSWjxQOlLTjRIIrmv8ehSD4jW9r/WaU1gq9YcQnzrGHNfPt
AjntguiAjJYaLCWqk3h9cNmjCUSnmLAgMDjVn/zY9QM2J5kCNeKzi/LpK2VU4dBbWw4ciD06xyjS
MPQsy0cYznfdXE5bBzDM+4KwFfs+yPLpqg/oF9VnxYX9eES7wk+p3DxhXtsGxBBCOBsBLZGLi0th
Xc87/VRM+i7u82H+RMvE7zMZsnx70G7a45Siqx17O7AJVO9zXkNns23JCtZfVifR6xn9OWwhd5OT
49FCURPJrqRTbMVnfHApN4LA+M6uy4u8JHtTABZl7GsHzfFi42U9pEMz9qmXl/QktjE8FrKGfMuY
4offjVPtT0jCe/WlXUKtRmD8s5TiFir79A78BXYGJaZjMYpc2iGHVyoIGXZ7vKEiEr7OwG9WWb8R
zQIKoCKH/IBJgVVNcgd2Hj41zFKTI/6fceVi5KoQJHzZ05RPBypV0clbNRhNEo8qiiY56VAkD8k+
gYSQzZNcAu2/tSIOPkasHD2CvKDhwpnrVvR/tlL2iNZyf1zg3E2jL++z/mVlKoxMWaoFW3wqbfok
lLMJEtfshmGNccjU4azMO9gwYAx+rK4cxj/J2RdZ3B80yfPJMp8GAo9VqRTl7aPsWod97hmkNDpK
VY8OQC8HTHopVoPqy7pNgX9kmfuoicaHB6BgQogd+6PFmA1lbbdSbt0BVbpE6OMQfUFNH825Zvxz
yjwpONvj19sc0z5GuBXAShe52YwyDIrf0z8oEo7O2M5j2CVsfuvhYg16A06mvS8Z0U0+RMIjVrg8
qGbU6QW8anRXa3O8FwJpOMRMQijsxfuq4kEvgT/cZqaMEOTFAxFjTj1j0UxE+lirkKFftOzJgh2s
j8ZPGwWSH2bJXPQejDhXikdA26rMxM1lgNyc85wpSBtmgkZ+lRjO12eMnwIp8yiOaWl3s2hrM7ts
IOvpGvXgRcZ5ImI3IiR3lFQOEsVakzEvMQpzNfNhcE2N1N9mXYfUTvyoflwtfnwI0X37RthTOgTK
YNK7jfRlhMCe0l+8y1qA4kqpuxwHBqMHO9okj5N2RtFDASPzISDf60VRFdHZ6i5jVyPdMV801lNe
+sBY0x993t0fE/I5MTxAzhrmRLdZnSAyy40z4onw9rgDeNAWFY7smOVnuXmpY4yrrenW4kMF9ROr
MqtsQCUjUeBmYROQg/Uod1oQ/QngovZfpknqpPEW1asMI/iRL5dhuUDjgs+1bAqdHFxv4FhlNbEZ
Q2o/FqLcLRCAVSKZJgggIwfe/kXKcjTg7hvlALCuOwZ9uGGFuJzLnbn9o3rraB8xFYzseqThO4XP
UGQKFdqbdKbdUxnkpSBPLCMgAbyrB3TtL8SslR0Er8g9buAj5JZlc1Xbw+MB7PgqKY6Qfoedwr/s
BoF63exzHQWQHuSjRtLaTrF72IwsRxLAjptZjQNXAq92mfJ7nQ7OFjRxdknHnomgIdhsXeGySuqx
aCvH8bwsT+HJX26aGexQJWg9O0sLNNF/yzP+OGRt/7U1AJfyx6zSU9JEyKsFCu1Ug08/NXM0f9lL
E6c6A/E2jcrU7iuhh6+EekZGXWoxsuc8MHtPthsS8iwmtuoj3Za40oiP/z+cXWtVNK/esCnzwq4F
twnCkhimF0i209s+5jV84cbiIeS8RiuToIpqSaYOT3L/Uh8XE21r8qJ+vQLa+cQL0XYfx+v7B6wZ
0K0BwVN3lHfQI8SILOHksAa9CvBk9flHs6Z1jnU09+UjYNhD3KPXK+b7T/QZBKVGcTGMs8dl0DGM
sbWZrugrw66lismb004OkL6nRfv3hJ3+TSAyKuzClmYc4qa9hayY6xUI3IGe1FPj4/5/eLrLxdDm
EvX9RXbVssmgStr7sUKAi5Z+Y0GduifOlj5NfPtrP2CyDIE3qLZda3+HCF1C6g0nuCepzW3XxTE1
lBYelDo2N7gzB+78uSC09h6PLBLbi35KXbBlYE8ExiI7a7icNT0NMr7zuGN6Sws/wvwapaoqrV/K
v67yNieXBvHdw8HqbZBHk+hzm0JuHwv84XJdOp5NHmAOYkINLzYj0kZGlqTm2emk8GwEzNTMBKJD
NzYzKjeBUwwPRr3tEwqJO3M0pHE30J7qCfYM+2fjTwxZqCVoKzXdsmHWVnyFPZOAX9rMZW1zFiq9
k9XQ7nStiuvlaQbo+/YrRbwXySudHtXyk9+hLLczjCWOnb8NoK+Zd/NPVgMiSuCiAsnWB6sHCC1u
VPFBXnPzMvzRri1uFIwhMF8gcCTk6VGAhnyUhbvhBMNltTtuGY1k5Nsb3ZCEf+ecfT/EV1QieUnk
JtA3tPVsFjxEw+TM5XmXx2ywh0/YcazVmc9Bui/Kbd2+s7/hKKouj6H0ZzMKId5JIxpgbHx4H5Mw
T61vglSWQypjCLe8oGUBKAlbkNiErdBczoJJke4eVA9jm2rK+WOvNEIjEepr3/RILzOw9pjR818J
iYi+w9TfzP0iLwP0JFQ5X7O8/7wTbOsQ2gO6Md9ufptDq+ZufZfTYp5rP/p+xDI62LdWJPYtGRuk
108HPALQnGBt7vm5qoiCSvH63JvH3oXgi+6L72B8BJTmlyEt6sWOLWcxumlvVY7CdPMx3LIA6ZoP
BACER/9v6mgW2HW+pcds/56RfoeBQXV7g9+80hf4fMce3PpbRjR0UeFovK4lZSx2mtNnvyN4sHIk
iF72bEEms/TsFv6p/xozV2B3aW6GsTBd9GslhuQIyUNVeOtQnMYfU8XuKhzopQ0Q/jynG/NvrVfd
SqSkKnHsc5E+qZ7sAfMDQgIf0Ed0+j1elT6X5vI9JpEt8nnV5DFTzGOyNAIKXwM23VSYvwa7vESw
lJEyhAvd4ccYGuhZj12ujNSE0RnrsF+bWoAVdNWeFbjwUfPfFoRMbphpdsLHvBJpsI3nn2HERjPZ
X4WS6VHR2as20fJ0xLNDseba33kf4eXnjzO7iDZYtYfk5XYhNRHmw4Q71gbQw9FfXsd/GrWbE6u0
wTbTVreCvS/onMca6Dq/hFw00i7yddnNq9DRNm4HdsbnmYq+Axi2Iqc9u4XJ20MrtslH2PJVEJHg
D9Frdbh+EAvn+TFExI1J5oRyVa6iPGjuJmsW6pbji6vR8HvasYHy/+sER8nErGQSf0bBzaHObyNC
EcMtGE2YIWF1PbhFggsKaoQaLfxDurJo/5naDZWZOJriwRA4niv2bH4Lbp7ED7KAjhTV16uXRYMX
7AZlzykQvW0ZtxpvdMplUsGBSey5Lsn388Adon2kjWaeUaYXniMmMFShF2gInnlfUfiX5raDCmYa
VNViuOTgf+Kq3sKAPQOGPUIMs2f6SRbSeAw9aobDaV88oXds9XD8unxVpv1wXFE0EFlIIf02EXPd
huoSiChBrmXXj6Ewa7m0e//4Rm+PUCAI6cCupQtz6xfjBDBoGwxr/YMQJfoK9KUf+5ZWObgDLvGt
62yVXEx19wR2pMJpOIRgtkFiX6vydjgyef2wQ27gP4GNKxnRifi5g2SluEV4NTAPypx1P3uJdd3e
etlAoNe8huFoOZ6KEUbQ9MEv+Jpb7eEBNQywRPTjBhKEq2J4oLOrEiYca7iKrn2VO/cJ+KFvbvg1
51+gF0NvkfVBVzcAx68ygQDLNol5Bn/TVrJoFDVhK/CjLa4YHCyC7FT46z5Dy2m2e3egnenlOW2E
DlGKGIo53FwfjOuym4YbtdzMFR0GPCu0CECdxAkaq2lH9UkYKcRoCD/D5aokoqnQorjxoKl9GLBn
G+gueGKhwePFLGGlulT0voVuiz9+M6zUfDjotgRMvne+Y1ecYT/VTjdXmgHlycTbVNkkzKEFXVI6
0z7QNL5lWLPbKaXuTQrsDLdQisH+/CYhZNuRGlaya8xR5QvKNaPN44wvY1xUKDAM9kCZYIik+ZRc
0yeunGoTtafnvSTBPkV8s11PkMLOY2bW/lAzv+AeemJaUMmsUzVJX/AyaE77OLMFFo7343gWFFB1
B3ZWFQdY9qbzJ8+LCLG7uUlPVT66qPjPYrbDHy5pwNAQugdB4jmyVeaUKxbnt92gF4ZRX54yaR3L
73fNk0f3zdR/PAgk783ZZs0FOIHCy1OlVARcS9jS/IR9nbdWQe3jT5z0EcFBUjH0a1nnFLUdP0Yk
zXWaJzXAHMhOb7e1qmDg8ZcMIbkjUy0Vq6YPPdmJ2eV0y4evsLioAFY342zDcM09T0QwVp1hUoal
19o3mErzqzXXStemIECQi7T/PcFE8uAqkSE9JHkv/55WpaK7ptrW5F3LIokUmulJ5plR/WjxrYl6
DBF1uHHptudlg6bmxLbCrMhIzlLREK9bvEff6vcSkDeBseWyQm+azfSLC0pPVWWJDlovVmbogRMJ
3ttQZOhEHVjGneKzatbuS1oMeuD/22ivirYdalTz8bgkSAGvf1WGNMwmnaxft9PB2e4rx+yR8kE0
XZ3efRktkJVL01Jffe/5HtwUgZQEk976+iw61NDLlTDypSujS61pMItWrbZncOKMmLjk2GDjbUp7
WPR95eCXblY6pZx1t3LBpRsro0k5UXfZ4j/TM/OpsKfXXIJ7whK+nLsTSED6ORoDRHWgtfRG7Fs8
sRxqACc0Tv5BFVPiuOSinLES9UYYI55lJwpfSguIeDWCjSvS1yneWiayEb89uPGaYMdYwcfMWT2E
qOOUdQF6h2d1a9w7zHicg/4yzhX3srOWbQT4foO3wtjvMYjp4FPmWkgv6lcTfNvb4xT7sPO4r5Am
RxwWeWx++20tT7wdXul57xabOCu0oTb5iwg3KcnPwbVdfxV78Prldt9LqrsxjMk9YcPEL2N4WoEL
BiK1Cn9dDJOPmenSVPZSTQK5Eji2fYfLJeeYmP7PdRrfTxVszvqejnGu8yRj8VlKNikQ4iBbRG9f
fdSfRWK8fo6Q6htGzkPvzsTf/kFi87JmbEjQ8J68QMBTx+Ss6kHd/wO2u8BJ4F1y87LOnbKAXoAW
5jTm6vPpQXB4EqrJujtrzsUg6dfjSvSKLH23uRKyI1f8iKm5hVWuGZH3feOVuvnQdDsy34ACl4f3
T26vfERxcFaIGt7yQ9bccPIHReGhcllJrDsxkZEuNptbb01sAsi84fPijvW20FnOivOIP1+2RjzB
Iaf+T9Jkf75azBzvqSnH+vu2VFB/uDrsIzuVdQfhoE6n9RttFR4FTNjiXAelmCFtG/CxJHjkNGBA
BxA5hfhSOkjf78UY09RpAYlhCfPCSc7qN6YLiF/74+CLIBu1PMLCUa73tC73o8GidIa/5fq7wJo6
Qv6bfYgaQX70+og5fT5b7YOwo9Kkk6FvgtjBzjtyqPIXKogDBNm542ol47Dhfy38iC4tpbhep8eC
sJ78nMxjvq7a8ZKGdChx9wPvUcM1AcGWNtFCrwv+khJBtqdZCi0BZ2TBk8FHriQww06K8DA+YXFJ
r5RjlRLPO4MmeCOiOysSyL33ZulJNoQmr6Rr0LOfKoXjnvQ67J6MVR/VjsyKecrO1DkuVodmYMwU
5A97c51oMZqvdnFve2LTBmO559oD44oQGF05UWVzzYgKZav/cge4vNp+KteEmKhpjEEMVZVp706X
WgHHwWqBZJ46eUZ2OOL9vSAAuTaWNU1N0Ttj4/fw+W6Sk5w9orRal8IMM8xSSJFdF1LTfstrEsdZ
r6bnW2VBtOFr8OmIiwm5AH/fm1jM1im16H3bp028HPA4dzSpMgoTEbLoDBFexe7gnO1Zm1N6cEjy
190YCpm0yfu5SHCySsE83Tz1NP0g83kcVNfx6CuNlfi60DVqpn4mo76NU2g+OpPOcsBQqtTx4mX5
ihOnz2F2y6rK6cpimb7uOdSOhCx7SHREb9RlIWaaXMfpKuQP+JlJyYvnfjrgRLpcWvskzIX3OXsI
lWm/Ku9XaNTXqUOjfQ/eWWfSlpGqyJIHWur+71uxNyhSN1KkAqsHFjdXL8vUN5BCqezoU4vfZJNc
8tZ6XFyPUJNpp6OIDKAJcCWleQzcM3vKIzUzpvucjroMfBV/kH4VYECfLu0fHIjfrRbMNCuJemeV
MS8CLnV/q/YsYm7hDMumRPBRdsDemfsgfts2iC98B+bq3G+Mkh40FtrT/RBqZGtXuGL2WM0aXMQy
3LZ1dVy4p8+zCRsNLcZNPj6/DWfLPujcL2/21xg7YOZsn2Rclikas5T7aq2JV696WoMnbSX6wZTp
8pBc5Zw4aTbhCGsEQ3hODcdnRpL43BZr91Zac9cNLRcNOUC6UcY+cvbQQtGshqNEzW9QEgB8ITg5
Be11Vyic+7jba4K1GO+BRCxPdtfD7m1i8gT1Zpqruu6nz2nK7izDeHTscWo5euRz8Dwiflj0n2Dy
LpknxZ9bZKLs9MXPa3KSyyJ9vrfOqCbValtbGkZ+DLUdifdpcDta0nzljm1kYRsQVgpEAVgdWAy/
N2Xn8AjGhsWBtfy/yczblKkLBS1xGeSV0XDIHl/A9BlPfomW/BaIlOu0/38SLKDdp0m634lkLs4T
lojBUM0/HJHiw5pCHnN9ij0HBJ19GfBhDxAmSB7n5FGZxfZvTFE4rRL5ZLDiVaCpb/0rH6fnHi5D
w/2czO2ZEYb7TtFX0ot0w77iqRDPFM1/FgqD70f5U9G00heLhdGKt1iEOCn27EdwRG06Oi9HMnXT
8TwLSiCO2GgczkNb01/WK62IfXX0cft8JAeSnX4HNQJMNVE9DevTpErpQuCcgRisscPMqUiflj39
gf8aXv5HNHRuZy2d8UFUuN+GTJ84zHPdyD95PbfSBvl1w//9YBoR/uD7xyeSR0D1BdtGHGkf15mf
XTG06JbmdSN3vd6eFxR0LOrNYB8vyL8qWATuUVw15iE0ZQZZUnMMhA+jUtSDQUjIfN5n+KEa6Bwl
OZst+1DgGwQFePTL1ocALBqriWcnswAx3j7mcYnY1cxCXlBqb8IOi34t9zUUHu+NZOQ5dBd4OnTA
mTbru8BDPBATBQ6uhumTiA2Of6cmKwhZbwYwKDRa9/U6SDzDQEOOcDyUDdV0zIs8i6zJUAsFFyCP
XlxeuXsg9ZkzaVFfT2hff9OkyxBYq2b1yJXr+j/Se116rH8Qa1hxoQJ1kYXblDQpxcVrHTWWWp/d
xQ8ZO9AkDa0slDhk/dz4pDe5pUvB+t+ci1fEixS9eqdNpuea53KyQv+PqzQH9YAdT2hs4VaaFmLU
cT54AT/WBI6cWxdae7ksOVdRnOnNXzvPTUdtFtoLDGnLfqbzlgQqomczBMN/3EG7+kArSpJ6x/pY
zMhEOlbYt+GkrDSQqfBjgPewE6z/QPAsc1qt/2f1QsKXqPphzPTr1Q+WJ+7fHPwVMRAR4+vwevfe
LapNM/TLNP3ruVjXv65dp9wmCblCygLxWOWIIqM2gQKK2AuxLPpcgrn2YhngMy73Lgi45w+EMiuo
s/OWYwuyd0A/WxmBFzLRx7aM0XNehwy97DrUr9PkklyUPyTg1p6Gf0242Vye2FI0PpqcWsKVxJHW
6JZ+a7Zl2DBnZGANOfvgZji4B5vbpEYG5kT15IdNsKzlITDCMvxjf+tmPQBxPGbFLyx/ACc6rRqf
kVlGOg070TiijF7jmTR8QD9MUFrNS5Ccf8H1WNjAG0xAfe4LjSS8Gsn22IVSPlQT2Fygu3pmB450
cRfKBX2dsD3VmNa4Gm7zjIyXN4FdNLk3OrvsFpdEuYmkj/Ju2rKc8fV3SoQE948eKvYvTGcPj7wM
xByfp6yuad140WKLW4iQenSgTfMlhw4vI+HV98Mz0mgyIotkAU2MPBIGWXBj+mN/RyPAohGhQsY8
he0jo1V8GY4TIsA0vuRZeXA++rKEa38+3E2nqhUwUAzLsut1+D1VAWFyuvf2JPKVi6yjHmOvushu
nhO65BchlBXURoz6LDNyb/vjKoORyv4CjdyiFGIQpTvtfDk74R5n48Lo1i3IpkcaEa8AYao71oE5
YsZSo0qjvMJctjQ4jHxEr9z9C4vXJcy/Ih/doN61PP9EyDjqHDfZD01ux+hn2Jq11+wXhuLgoOiI
y3i9yj7iQcz+Q4DcBLuUDnmc2Ngm73gZAIlYAGGo5cHTY99sFKbISebXK6biQ1e9caVt4e8dvdZ2
WwgWa+NftlCGNl0um9PJWGre59aclZqOnYPcUyc7IzROgpGTymQxcJmkidYt1WfDVSQf9vVZ+brA
zokuIdVYCWLBChiJ9TQv7Plu4dM18SrMKhptWfELfIOuTEwF3lgjMo7j9aqB/Csr1JWrYFrDqIq6
ONi8hvDFBb/ADEemwZBz8KLenNASMvafzu3+uHNU5bFkwUJsjxmCMfAgmQLfVzuPprdpr+aO7uDC
EVmCq0cqZEzWciF0nHKPWWf+aPbn4sxNJV+C83cofkR4dPmXd8EHAJ/sMMKPXHlmU1LaODPy6hTX
5wXK/NWtooXCgYv2R11gCyANL++5lptaK1WB43l8JJiQPHHgcf8GwZn6svc11j64fI1NCNS0tY/d
R5K8WanA9qH49dqzh+mKauf557Pvyz51Ryj+Ur3h7yh08h9VDpTvi67XP5o+s3/V3rUHR7n5KFSp
vm/MKw6HJOwYFpee9LgIIjbrmsRawt1qXpZmn2njnPXQHdCKzEDVIwuomH8Y+SgkrtZYMdDxpTD4
16H50U9HFZOF9YGCNjKSLV0sOa2wJ9EbAKXqdt96W8eDXRyBS205hAcXzgL9/wN0psmyJd51f/z3
Tixnva8VrupDyo9MEJHm1XgE7aNq5I+nsWC6x0oVgA6KBg41N6J4SZapemhOcimrn6+dw8VkoWag
CXPhaewLMM04PtKh4/u+LlTqc7PWYFjI7DQRhFrXw57unM3XQ1RFgJtDvqFRn0PWCGpDg5PvO/gD
uxdVgBhcsAYlwG5L47TaCucPd1P41gJMwr17/ZKhoWJ3F+OyciYkfcShHw1iA79tbyhzXKb+nVFX
Ue5F+2WooMceVHoNFmvrnkih60CA8vlk8ikbuFqmoiS1z75UhvZe2XP9m7f4vc7TzkQFh53lB5uF
ALDzAFeDJEDJFgGNkXb2ZTccvV1ViAmNY/vWotYPUOzLUln1SVL+Dg3vQJITna1HmoDn/JOW96li
x/Hn53bTau6jED3CrwJyehWa5fFBDcKlanPZun4r7/uedfygp9/k0VSRZESOETzl5avhHcrH7YwB
ehj0A7BP+MWyr85967fnaKDRfUL83iCzDgYZ0z24jfoJDrwiEfRwoO4iNglLN2neThZotFj+KK0B
zg2991e3b1neWdB002uzv5vKXZrvKH+xUQ8RVabilcZ8KmA5pNGwd5+lHCMVyRcbhyOYBoFLn3ym
R1gd3u3q9GcObopt9iz3t3XMVStGjlpJgd44hDOZk485nH4zfbeaWGBR2P01Jy/TjG37hrqgyUiQ
pSHY6zNEFxsv2NE5SSC3MQVRiJG031nzqD+fClMtQ3uePaOuJtqT3UpV7qCsyNqLNF+k0+gvv/68
QwqzSZvz+uQefyvuVMHccZS3Df084Yjdye4Gx1ORzKa+HurN02huskBdS9DKI192Ofh9Q4h4sIJK
5PlqkL3dG4kXl2ThwNwY8yFiS9leJDbETJuHsKJUhwU1n6CEUf3ELHxqmY0nOcEYQZENfNq9d9SK
rq+yKKQUzWNeWOb4XD+bHhmKlFGmj+T4sQV+33fEl0BKL+RlBBXkH0fIro+1nCD0dEBRBJ/5almA
HW+p4OiVCRbIUk43y+mVqevzNLp2h6J9vgGV49+zJvzXGneHYrNwZFr9DgPYLcmYAkHKsr9pqMAv
c1r3YvYn++0OEe4XJv3qWcVTs60UBM09VRXmcVHvjzS5iEUrleA6OlnIBw9hU+ZHMBSQH2YnWe7Y
RyiCEKDqqmTWkO099F5otWPcSlDFHgy2fbuLNGIFpDq6uLfaqCR/raTOPfFutz20yyNKM/3TUyVs
J+/VJRecvB9xjpe5Qd9lvdcPeu3pV2lD5LLgBkPSSreUICgwsPsEp6vsQ2qnbm0546CRncHAatba
O5MHcX30yGmkFlwgI07pp3jJUWF5i++OJivQpiGyx/mZdD5SulytZBeNVkLw8YgZQcRyZpkHKIIT
Y693DUVOs1JOkLJLUOOLNnzoACmcTK1SDQIVLscMCRknRG378LExPPcp9htX3NyPDEKd6M7/r9+Z
rbBVS6dygIrQEkhH3M0fE37fzC7EJo+HjiC15vnXS7sGptbIpc8yVyq6WUFSJO0JbT8EJNmhDefp
p01LSWSobhAAU01u26v6OWYuYWVmRJRzZKAh8ekWd91HCiJsHvRgIgMp9ykLp1CQ1yyFl+bgrQtB
UzbritXSQM8eAaU25P3Z62h+n4wHlZCPkHv7juAH2OZOW+hVUuFeGYdAFUz+qbKNaKEc28WueGt7
hS3/JZkvXKSqqDm8cqD628z9HoUx6qvc3Sfvp9/ndtzkhKSLL5fQzAanRZNMNcQ1sJTEpVqMdyVD
iW7a/DBDx7BQh/NO1oPSgq7CtKUASza/D3NYIJsuWze65ssYJYbGzjewfVPhSwQFulaoaBjCItKr
OxQftthWvBy2pNaA8tGejvxbZG+MRHuH8062oq4r0Qo8bJ8nU7/TlbTLSmRSDAUOrn6Kms6RuFLd
RD0ZIaKHcm0PP8GL28hOppJkQO2YbIyGdlc/Ddm8h4wQxkvxEuFjSKMsGDxex1wQw9vt+eR7QpL/
3uncEBbF9jNT/rI2ZXmB5SwjNjDKB0kwS4f3gwIMCG4BT6xtC06LqRNMetiQFVU8WskZDeI5Stni
oXCwUHYjLpFiG0jcHSTwKWXowZqUAZRHMwg99D5BJXWE6PY2FB1AoGNPbtsjy73eikVtPC1+BVoP
H0Bhx/Rex+iJ17OpOGtNSTGHhJyRXIAoykOfdoOtzkAOjUEUKkDTYYYxj+TSbI6dU50msG2OSG/t
bFZn0N7Nh2oK/b6YGW6CdooYijl5j4lTOOnBNFEfJ+BND0qBn2iZ+a7AmVc2D4N23vu8zzLP8EoF
QFNUrv96bIumcYlJcRntgwiH1N/bUv4YLRsWkZ/4tGMGHrOfGTQaSZSASeV0WYsaUVcoS290yh84
b/xZHYRjKwlcyUFvEkOGpiLA2DCsymoA2sJVFCWU3hVO98tdughzyyXiOCtBDwgC/SM8R/7pW1p/
IJKQS4Zy24eBxTT+pwLT5BiQGqbtuUaznIH6aJz0chatKi1b+wo1oKyz8FwTY8vFukcB4zaWY+wL
OkSPd9GW6Y9I9P2Iajlbt0n68VlXiPHLCEWDzCqixY7eD/5D+l0M43KQoJaAG/7jTl1aELtqEWS/
83FHZ2GfVXaWbd5HrhsgyBNgjAuaLhEKxXcyZq9yzJyIrp0896jvkLbU2yraGObzJ1HguelWKjU5
nDM8o035cx2CC6HME2ajm7DZt87xhCgWR7K5zZlfOEd+Y3eZ0RQUhy+bx3TE8mdYVaE7ofp7X0oz
Ra6b50J6x+0JUdzbTDziRIQo1UaAkTc2RmxXfkjKQrttVce4xIabjrMH/OYByHTDkx0BJitbKtIg
U5Y+j+wZPCT7PG3X4G+crRY8MD2LeONIItaN9B7NVbw+hk6TGt/BPRxSeVWELncHyQQ9mMzDXo76
yr+e/msp8ot0zkOQ/d3B9AGMQh/rAESMs1BcohR6F7U5s//MnKsKFy0Xy/ZR2p80XZ+MO5SrHB7S
kUjArgPaOr/36B/Jr9Su9PzsXPlSVXt2W99Y29+q2UxRSEmXdz2t+mR+c28vPl3vTWH3KI3seUIi
Gyvnv0pPSWLIqsikzyaZnU4RT5HN6PBkkGOe1uTUGsoQQNo0CZO5gG1it6pXO5VZNZZaBYPliGNk
S6uZDvdnkH8Rw7prnfDit8UdfZ/rMDA3aI37U45eypV3jji1soMw1ONVMfqqlYW+JpKdYjVkARX3
Z6wUgI4IynM8bZnoX+jFnax6YlAo5DCrn08aW4w3jEZnS7gvoukES5im2LwC29FySuJRD1ev+PxO
+SzLOMnAgXNigz0PmakT0lpYWndqM+ynqoKCij48NEjqeQJBK293QoNL1Te8jJTj9GfZJAfrd8pW
+vKucgoGn0ddlN0IKdGJ5TxJdExLFQPiHzrBpcVkBS3iNb/bOWOAsgpQtjZUs1uiacOMZKgHeL3G
3AWO8AslcYwUNB7FPja9Vm8OVmRTocRSd+SmBneRCTi7odcBkenJSSCgVFYXG5AaCoEmD8vZmCXL
tXECfVYiXkwlLVEzC1VLnorcI1TULtJrQdcV9YCv8fZjA2TSKBpWYnAnEJq3x14wOU/VWuSle+PG
IKjArU/0IPQ5UMV6Orv0QUu8sGR1ckgZ0qR8CLFvs5/IKW/iDP2IYHqji3wnV2De75ZxSn+JUWyu
v0hlW7eaHG/aseP8pSRIHajGHZ3tJEIU9calY7Rrw1AE+PRsIL97/HMwSg4824lWqZEcMHzLBi37
z29UJzGVwYdvZlilOV/5UIxuOt9AoPc2I0E7N/Wrb1ew5p/oa24w8BbPHCV2sqH1RGyKjH6lXwtf
YTWF2wG2hQksYjrSiaP8UREPmLxj3/99AOyVZHBMWbSPCuVWwJjmrYqBHsHmqdtcacMMzK3yWPPO
RA3Em7j6MSwt/afrEa/+IGrh3hccujzLdgS6X/2YAzyxzT9oSb1yYcVAdxLR9rJr5W1TN/hqHWjQ
IakhAKbb/NYpr+43nH54tO3Qa20INhy6PwQ6C+CUGxTrt3eVI+8HqPeA9Bhw0hP/KVB6aggeUdNQ
GzCPSlAsehGuH2zkQ3r3baWLUZIcaNuFjI90xcvMJGw4RyQOwm9QDHxgybi4GnWesiCEKq//Van2
/WU2RI6Bi4my2HMQ5N7oHPP4LYrd6GFKCfuaaNGbKEDHrMkSyWgJcSMQ4bRkyQwvCuMWMb2USMrv
WiXOU+8jdz3mWDmwBSufG1nLVefPMhZrnTWWmC87w7p86cR4hLongm4CHFns5GDxzy4Naz++Cvuw
aHySW+boWWgidSkBQFP0ivknJx46Am22GqP86756Di+vWRSw6CEuGv39n0GkOfxdhBSkn+pe1DT8
tKY8QKSzgVzWWP146U8KHfvcilZUXTMTKsHvbVWywwwVF/5zvAV1zhUjmD9nJhk3ehYasz2vG6tg
9joyrw2zdKITdpV4ASSme/sSiJWawRGah37TiuZBdS5SnXfTYxzMASJfknURPEY3cZgJaxPJgYNr
oLsuHWgHCdh/K1W+HiDEIjnkdU+O9f/OImBLOrMKeF7c+MVuoWeawFiKVaP+erUUgGNgTxugkOhJ
1kx0/PJvWseNqIbGYrICjCQdHbRorSWEFu+XW5LP01oG8onUv9azcskq87/UWbhk62QFSqqLwWFc
3keKfkst2bwjbn/eiNgt18reH7FXa8Ct8WlygbIc6zT2W7RMdzqbfKJxDH1gYUvW+wMhHJ2N1JUo
TrqJiivyPZUhOfvjwOZuEK88CcxtdgylSE5T8uKNPfF9L7s9hXLVgumN9MkWYpFfzveG3tXUAfO+
N8aIDFYYXD4QqGSK0v6ESA5Kb9dweWY//fTgJ+rpiqmVrYAGEYopUO7FLRxBJYEsxAkL9XqeqNi/
GsxstHjFjnI5AzsMMLmzUx93dmng4vWjrSFa26lVUeyHSKY0SUAqYPgisof4sdzNEmRTZPVnZhYH
HZCvxqpO0RpNoV/vX+k+wI+CIb64A5wG17RtyiwtIvepKn2awPTIfEcpG/WDMDuvysCChMfTcUzF
LvdtTtJqSMlEsllB02tsuhNnlhhuL+KCU0QFVprD3SQhhedwd38fZHrDHwZOtnzMs6DMdev50TPY
J87RIFzv2AEus6Cx4Th0jGGb//hWhMBKUwha52UowjAQNyxge7Ulk1mtAaZzKzELVLdoaYg8YNlt
vUN2V8H70E6EEM0P4pdh6KYwu3CmpH13nAsA8Jq/tfvigkVj8WWvipGk3xdMpVhF0cg805srbkRh
s3n5Y5Oe79ob6r9hSsMGeDvWhLEWo+Tmy9dMnpgUVyEs+E0TMK8he/xQ64mbQJzffW+P1b8vP+xD
JoMBltzVnD+tCZBAbjL/M49hEntnOn/E8wq/aZAsIXMOJAPMhWBf9SFLWSOROw/9WMygGmWtN/lf
4rW3GAwt/qYAJbZWCfLX1p9m69j2cIPRgEz3nz3PRy+P3aoXa8cz2L/biR/YLLmC/i2bBjsFXY2I
M2I6b7+RpPH2mWxwApYvrjsDQz+l6cFIm8tXWB4lqteEaCHeu4zs47u2QS34b5ym8foRzceCOaU8
1cyqduQD3L5v4ozPXSXHbSYrmm2PhL4HVbas8vX1vfuvuOoLw3Ak/w7JJWybEamA2ajDpGix2Te5
0nCIgXaw+GjGGsFxr5ltvoWCk/0jIViwLJ/RIFTXoh/6jphV+ibFmKaGsJ56k5ehy2rC8+V8Czn4
VpEE9oQtgSrS4Jql+n3WAPqrUoqj0xgBmu2NQi0p/0kegD2WDzgkJ8HWaLe+Ru0dBgVMmquIIlkx
B1YwaRllmSqD21+6UeCdOlRH2yJTwXRsCmhrFz11M098NKwm7/24a1cK8vlzrLVEbzkI11xup7wu
xA5G9NRhQCa2x/EoYBKxtykKe47FOEyj7z0a7M4KI3ZZKb47ciJhEkeXTTV9hWyQ88nfIdq1+z7c
hzVDnOlmZQrhmlwP25pn1zBUrUrBqZZ6wOq+ZrsGyHxK3Wxds9lKTTfOc8weG4WZi2fP5H5H/LMH
g2ftHLrXjpCNTsDJPFGC8B0oiCMHUhX6tw3GOqRRyrVlWxzT0xlIZaYCKis+WayDbEfC81MreXmf
I46Itd71yHzb3rk9/dvyl/JoCii3mI2dF/yT4CdcAeB9mVLPGYc9zAL8VifnAXZYo+M5wmpq6+9F
+ys4qzWcmSX0tC5JrTykbb6U88d4n6PEDjFRYml8rtZNVWifEooO/UG/pL8x4rNX0XaDHb1P+3Vd
45WHbYuD5DUe/DhXNhTDUyTACI/4yYbT/SXKIC78Flo7TTN+JXXWRmhbwHRJwAShvkrsmihZO496
OvTasykJMe1A492hjS0zUl8+cLGN5gm/pZ3BNNTVaB5AcKVuPtqSjGQVefrGVFtX1o4CHv9qcoT4
RB/UaBGYBVw0Dootshqd9mtouSa88903L6co8LdVsq89Ltq9L1Mtwo1dmBEODMAATKO8JmIi/CtL
3Hm6ru6I2xYcfNruEKA62OETSdFNNIsiYaj/yjYQujlNiGMcQ1+MdUE4uyYoL0ZBO3WzrXVcJ+Un
L3qzptPhUT44YTypg0z+f4YdkN4fOjSJrU7F0jvbcJGo/H0NfopxrJuxUjNgKmz26lg4ZDO+pnNa
L5hQIxXRq1oXFBi5Xo24rrFZJzE7lvEctE8xv+IWPa9ST8CJFlNCMEPeyGH/OkQN9YqZiL0IJm/K
9QD0kAjmyJSQSyxxskCcHx9W59OBFIbX472SkLe/oFO1saQtbAIzagZTuit/5T54Fkb9PZ++VOu/
XBHtwuGUcOPnIEwDvgaKs4mnuZUXVaGqsX3Mcr8a/wHbGacTXIgHlMbCXTXsxwd2HgfkcGf17Hqe
wf3t646D6ayDnvreQmdD9yaui5Pse3dN2UjCTvPsqvFZt8L8sbx5C4jR4uJO8dYtqvIAwp4fGQK/
i4iLIizA4iH8qNIlIi1wivOL1ONPoNoV/Xl4fwruglV/DRqC6paK14mbwqri0kXLLySAaHcg6dmo
A2KRo99f3bGC4ouavGPwwvJDwvbRyaTr+A1A5kWHWbR3OKRU65JgHKNcqEMGrX7c20ag3Km3Oyfw
s3WiYbiLPxcPJ6kWXtz4GDdUxCEB0leOiVZDTENTWLO96arn7FskQyGUbspzXJ/j3R4EHRK+tIjT
VnJis8rHWtAvmeh/1vOYhUClQY/55S50s88pm4i95cFYs+DW34s+0b2h90QBrcHKifzI2z3ptyzM
6X9kTcH6A7z1Wiga2KkX9h71HDcjKhDbY+GWlv2Y98bdL0lt5U6eLbo2kzB4VEj3EN59me8G5S8x
OfsGgT6cwu4gK/hd/CocWDMbGUpQWoJNCOj9sRreDf45ykDhI+Fhq1wJQaFzqNb22Gh+61wCe20A
mlpimRliM4FUgyH0Wuo7iEwQeN+dyoJ/yUSn11MvJhs9sYTrMHsnF9Ji4/kr1SFXDENn+hK1k0X1
HUHZQz6uKIABYjkPw1OMLvAMuFmaD38KAl6AfTFEZoP5YV72cgNg2QLHmbRL7tATVln5TDYelHzd
xCf6pm40DB8uX/YbTqCzfQkQJHVtw+oLF1mn1lYhinc7OUyz2/gQzPKJX/QUaGo5TMmdHaTfPaOC
hKwRjHeihhZv2UGOOL+j077RSfHP54cjBCNoyw4+7k4ZO4/Yp8lckYfjokjF0S54BSJWrURM8q/q
4WU+yoKgKlFM5KFinKwjZ31BgCCDK0hEQJUa4q3Ia+DHlMX/OQYzbD/C/XS8g7ygZneg8YhepqXr
PPgaCfGBpXJoj91umxey6MPLPQmCCNpvG388KQoivayYB/t8fpmf5KR9h5s33fFKGShFPM9V8Ysq
wyWldNb5E+4D+opBt+9TfGf97+jrseEtsr/Pora9kl7370+XdeJ2j60VO2UB+xfGP1cpzDn5W5+s
whwAn+qTFwPncCa4RiAPeRdGxWjARVDzoo14Nh+NWvy1qQBovbfYHXInlB8PIiaSz9bScTlLCA/e
ntWcfyWAVr9t90dOyMFqOWv8ndYGhBJtt+LdUCiNbAo2xVQ9kTSVmsMuscASQFlDvq/AS1fc2SI6
3rZQuIgsIk7vzuIG74K+eYeVa7vICxKj7mdT+onzJ/4z1Zhjv6j/+ED2z8weLIkYQs3l+qI8n44N
7N9cSaHD7XZkPlRTewBEfy9K/Lp/j+3uSjlaVAKqKa0F72PVqi/puikOiRi5NBBJodGKkBiirGeW
DPvSQmhP9fFDLsuiL6ld5hRDGeNCOCdvJV5JkgQSi8yLRed3ubayUI3Hp/UPTn9TBQ/n7hSmYzGp
o97jOK+hJ+HyPxXmHVWcvqSAFLhL92RD4kLEOIYwO5hyq0zDL10GRhmCDkQJZYp3YIsNz98mshpm
ruluK1pHXeVPVZSt2z2SKYrVnt9P6fhqLdGWaQRryrBWUR3+sf3YIoxH3EvrGa1bEhb0TrAjS2d1
7IxHwa1Y07/jDExXzaLzVb7ngpkepRXOxBoxRLLF68b9r+YtjYoYB4BuZyNMcoW+2OTh1Qhouif1
PlN5G7Nf4dz6wjDuj1Ia8vGl1JiqmDFMJIYlKSisSaN6JmlLy1InCUi4Jlure1XDTLTNH+emK3Fb
C6gpfUgJcrCip3qVdFnhM8Oiaelhpm8TtyxB1NznL0ANyW7CEPKsaxr2Jqze37j3irJ5HVeAOnYI
k4jtK40zsZlWkEBr3CxQnNWI7+DVUqP2TzRh5djMZr1ioGLo91l0g80rVjw1er3UaO7GpO6vt9A5
C2pOp2unF8zqQ7+Y0WIgb16efMROZ1TdRI/EiTVVzNxo8bt5asVyzePy2DhxdGJZ8OchA2Z8JyrD
+u5UHg2etytxzdwQp46EW6ZgZI2WS4Bs10/MmpynGfo9GBszHzqR+x/92E1S3fW5bAU1aEcIIUKG
vkdNa4Xf+fa44rsScVW+5gZsq/N/BZG3nDH/QGLiqZrxBp8sslz8J51QnEjL2Ke6F6UIG8vIiagm
qgSnBbjLmYCY2oPpeUoI7nSW4/iiF2wwD2rnFsGcgPnD9zBt1hmqEdR44sxqnaASCngEBsG+lwIH
dp2AqOaKntYh9ynAwJVS/KDcK1aISh4a/hZ8eGSNahlsbBCoPjA1oUgz4ord7BZpyjCtyQprYPE+
brA/QqGv7h1IkFbA/PcvWIkoZPZczobFBX5QoJ4vCHRrz2HibiGOzteRjcu+kuRfDmOL3TlJaC/w
cZHLlvTWCI4vGpe9bkNYUyV/w6uziv+6E0+FQk9DAA3kiPVz5CvYl7MIuoPFPYs62gb4I2xeh1Qs
JpQeaxXQopp6m/WIaT84IX95LmBMhdxLvDcgyD0D0CKT08ZP/7esR5cDkZbKg0VYG7FSIdDHn1c2
U0PEDDJ/3SaBJEDkrTbgYDSLrzbfPcMuws0/e+IGyRJ5FmxrnUMRnSEwpre+p0R6Bq+MUgvz9vHP
pRgdyI46p2+o0mkxqUF0cQz4KxpnHVLLOnMMSDL6JVLoOp4GGU/SByz7J3ck3tiHqpIe1nkdFCqm
WLHfwmBIM8AZUl3pwH76FzyzUzUE1cb8pGaH/y7hYk/06AtI9s3pXMhlHZF1usutbJLLR5D2Bfhn
q+pG2w2972p+Q4q7CjG19wEe7WrjQKMtU+kj0jRM4HXRrC8jzcunzQt9oNhOzvKWlAzfEWETjOmP
bygOfkuJS4BYDc/mobyyslnMjqY/1yMT6X7X60WztZavLYhL/afoYOHURPXU4zrtG4hf78grx1Vz
zCfQBjRFnHFbTs3RmgkyaLRmslpzQrzxAIBSz5jreO7XzjXqmYugFS10k/BV7xpYi1hJurh5Plq+
b7McGhQJFKHx9D/Bd00dOTEqy4c0R5TgfsjA+Nksk8pQjkoyvDfeTeHBdQhsInBXLCWBXbSp+vUw
JIcOLeyr5fkwUEK1rjiI0jEf9rTjUBHD5aLzR/nMQ7aM4vUU1ccnox2SmtxCONB1ZNQD9LjOLKUk
gIzgXwMNn8EG0o09bypUyedXuLEucy7/BdS98frs6Pu5fRa/slAYEcfBqAKwGAacdfgYZrtGHWS7
BWXYITaMy4+q4r3Vz1Pk3Kx/yLmli9Slk2pxtCXCZmtPZIQIoIpLL4SD6x4RO9Y+j/nNKtrcYrxH
sCqTqwNrUgAn1ikL6X2IaxUn7RYhOtTxjby2PBxoA4xmvw/p32LqpZe11Uh+bRZGRxpgFpBr1XXI
M1YgSw/TSdUIOnl1T2Mw0G+40Vhal7U4JDh5VThexrrWss/dElvAnzlPdvfWlF3buI07X8NsJRAu
zChsSFDicClzKnyFN0lHgG3poyYGD0TExkJbAUnVwlxV6A9IAs0uaVQmUhDKi/ztohdLODhLoTJq
EUcXbwt2QBP4mlDxuB0BUxbFnn0N5Ce53dXYkLVf0FClcvUB8wcrMSVLnI1FUk6HYyMU4+cIbXu0
p2Lk5DrpVbcyf9jzG1GBY6byoFjeBQWHuV9vmDH+RxEF0MmWVtpryqYqAS7l1hB5y8H3cRaqCZMg
zlbZPosKpWVOk/tD/6PR8UPm1Q9cLGIUjeGdNR5/vjd5vlp4PC8Frm98FPoryukVGW09V/ALs5oz
mT6jirXZCn4DZ4qXAqS9ZdOLt+xvfL35RaAsyVg1Ej4otmVXmBhhOwHKhgeRHDu5ULeKp0KGqAge
gtWQNLRmdt/IYzDbT81kr4aVWP17XuTN/UBJmpnCSOROTRPhifJE2KhC9vcwiJXQYxiQ4VY4k3+t
SwM8peXQxogACjysbFY45ALPXvMNS8pTzutPt4h5vbw6DoYdhu1cUYqrFjNpCMGztx7UHr3IoPWG
d8jvGx/L7d6e3Tg2MiMdwJDdTGLMd3Ykvyor54gybHlbITDRPH9VvkoDcKKreewe51ptVuvUaxtW
22rBoYsLLMet0m2V6nCj5sg9Cd6ExZFjBY20X0tVDQGAMgkR8lqpKFvfrTZQkcTsvhHQcGQctGDi
NueP9DE2tXhkfHXFTt2sqvHFzZudmaDD5p0VqH5dbe9lbAd3XE3b9bFSeTm9EU39ISA0R9i0vC4B
wfj2IL+sWbSFCfw1nOrP8qwEsDfBCTLPCJpDBvWYDvgKo+PrMjWYRlJMgyvSRiQg8wdIMunFDeS3
+4Rs1hUMzW74ash8qI4pWuMCPCpn4905igdDnC9CvkxwwMGzAN7nTurQ2EHwX7W0yclX5RNFgQbM
BKGFh49FWdkWsqOwcT4KL3lUcsv9ffpuGEcK9QffQNrupTmfJxMSJYt6VIajep3kzaO9ANB0St+f
+n4A5MBZRnEqVp2TQZI/GP8diPIRTAdYgs9CIj/1xBB+PLNap3Q0RTfYIxMWVFrnAXRLJ8Fw/WMj
jdR0BqLVPMVa73OSyrTYX+5ctUu5YP5MPJLScV8jNc04rpcM2XOS+ojzus5DkwfW4Dlhx7VfvyGH
oiQjs1aa0EPnKpdCQ2oQAtWJjSrF7slj/m9sqeEbNe+DG+h+Tun1woI0IVxTbAA/IwQYTmUIibub
t+jbehjJdR8noKljSSdngBKJ1vdif/nkor6uF22bwU167xcyZ9RmhWwx6jKHUfBMDvzK2ghX5/ii
5p1h7IlV9qGtuiFDwI9crW7CEFiTgYvAbrIMXTVHz+7WcyAOZOxjWUVBDgZJRDeh4eLx6grCgkZK
JJrRuW+0Eap5NRKnTsg6C1a5HLPTRTHzxQV6C/J0T5fxiFQIN4fAEhLiSRfsktF8TZ1R+CretR2n
AmHYyq/XGyr+13QbXgD1kChvl8JRCEOPAlE7Ms65D+zsfo04lhTJ6Na6jGkxT37IhU+6TqU7FRTA
ntBJibGy7PK/Axwj7NGWOgCRGOv8CGBxW+pRPYMfY6W1e67iJefld9mec6M0WM5aFGe+4pqvy9f6
YBvI3HQSGcETucQbAu7obpEiWeS9c4DaYBnKzp0WeAzgl35Xvt4dd5FIxwTNR3cNETG/1E9PqLQM
FQs5d1di2f5bTMzHaIGkBaSgQgrenoUc5wSZzKpx5lejAVQtXhbUH1K/CTJMj9CLU9RVC0RoDDBV
iXBHIYR6cBK6W+wQ9nWvvf2zZORNgt+L/VYECZ3fslItE07rONDfsVrdSf3GeNzoXTtkM25BLH8l
sOJaGmzx/F6bDh8mBNcFYLGi5NJBjAGt7yO98aLDBnSYHxN21otSt3n8TpAORd2170yZjeuhaki5
1bZWE2mEzP34qobTyDXRgv/94PIBpyakjdDxjA5ha/7a1xa2sCHdiI8e16sYzB/TjAEY8L7yzCZ+
N7GaAF7UoA5M9oQY+25eftH+5DhXMb8nOT72/A2/RSBY3SIViJhLM3tQzURcx/QjYwhZ/RrZuuLW
jGoaMRukQJKUJkxgNvEzjECJgWNouBM3EObAcfbT/FpvHRcr8VCPM/03//Tds9VLJM1PmbNIWYFe
jATIrjuwTx5QgSPqDnFeroPa5MtmDn4u3iFS4nKLz/N6dF8xPdD66OVYDNI1rgTppffjdt2/D4er
CveSXEvRj0OA0JaGJqt0cwtoQHWDznypZVvNp4pH7Oo8mOZtOYV1S5nttG4cPiBPZMtZu6VhkR6y
GxqdKGbUSWhJbXVmWEP6uftNW26XcTA0822+0TYijYab8hzADqcpDSStKuj+aUz1xUFyA+ELhCEm
dLNeW7w/z1A4ULg7Lq5trnUDHmkB3CLnWP7USddEtlTeE6xzYtRG+pElY/8zP1vQwsV9jmmKhoi1
cjPkpxf+t6lIeJJaT+P4ZBRmtbI4Fn5JgEd1E9GvLnArodiMUaIGz2nTfWi2WqDHd3j5OKGRUWJA
8D1h11EjQJxoe428/w83y2r0nPxvQfICt5D93Fs72CPPM5AloaNFkkvP6gI2Bfm5cATl8+Kw5rhc
3MNfcsMjRDuil5mSS2TpOHEhfYXYLtw3s2T9D9nuk5r392pSLfd4hH50+MJRbCcffEAssfGH1OYh
ENtsXjPUbiMrCcyNyDiBKC+FkbKxWri6AcKGcmSBygRTKzqm+TLliSrp9agZ/fKdYBrZGByNAPpP
cUebowRZtjzNC7s9N/xKlfblGd95BpkEmI08teVSwK8mziYvAtvQnTGLqrgGNXdQZAlqNeMDnHB3
WgD3ZR7Rb28uk9kPQ/jKg1DEB8pUb06nbvpcrJtyv34nzceOfyN0gb0Pd0Gk4c72FJgnksd+jPHZ
4wIq/Sd949pVCx7nMTwQDz7/3gge/y46PvtlKbr6WQ5IQmA8XlH1H7BIgrLefbYJOcrrt5+z4zCE
MLskAa9H7jNc/32fd5HLD2TB9swDVcmrT+M5STXVLHY7F/HLBHveRrhi8/nKY/i+5Z4lc03Y+lJf
JuUH4bQhvLXA27FhaIMMfihwyrCYXXRQQIzBLm3niKCS05V0bQtsEFUYu76HvzowqKNN8X6vHST7
JOjTC2/JhNiBp+e0/xekC6LBVrNIMMGeonBioukmUGiQuRIRk/xBcG5iYCwBbfaqD61mXvCI+NtI
GL4MNUzUsUnBLJ8ci3SYMYpeK6EKMsQJkdGnEW16aKpnBu7gvr0cMUPkaLTw3ZUuPBRSRnSJEwhQ
gO0mGirvkTqTgyqgRD9s6f3+GuvazqMhmf1/ompG0z06o0whT2iDSW9ilg8ls3D437ru5PXUcQ3x
FWrDGY0sG5UURQyy5y6vI+qMAQSxX1tkWEry2uTj3sDy9mKDOSC1kOM/Hzif3b0wNqTE0KO9Ch6d
X7xPOCx7431CGXVsFYDrUZV9pL+D+iJgxZyvb4uA75O/T6qQgxg9cBJvbABwdiw/YJMd+KcJu7FL
VvgmA/hwwwQs5nvDx1UpU+OXeEBqW2o27MZt/raleX2dJa9gCRuim2lMS37pO66hqKjNXgw8eAWw
zoAG5moAgHfb3XY9xF92M4q0XR6RKwS2ki8uZ51U0qU8uRwO4XvrexhzVQP7qH+omqF6iGByrVwR
FMxUlGO2+VKJLqIJ24THcRe/4YC5C98b18A4t3eUebMDDT74C46Uo2+axiSLvG+hIYuBHVNS6Scq
tYd7sLzvXSa1j1xtwmOGLW46p/G9F/uRvxaSpdun4ormRRrty1OQDp1Y0MsVn3AdiZe8hr6m1TU3
2x9g88j5Z1FcyBsT77FT/HJtQSsXX+taZWUjl9dZcVLCMAMXgDIAZw3k0VHdbVRKJfxB04+odpWe
bzaMYKd2Q4fRRMsm/lanF1UswLg0rnWOzyxxKMwe6FUv9Y+UlPjQ0YCnaJbZB608mWy9+pG6cfgc
mfh8Jt876tsIvtTIHKG1N+HgBZg/2ofid4De3so3Q1oyPEQKhlmt7IjWqlWL2Pa0r1Sy+YZry6z6
4mPFnpfWco6p6U509Xn3BG0mRdGtUeJUJVCGEZUONwqYOtiDmjSCduXf0zpH+/OowQgMXCGAM9Wq
47U5qgn1zoZIltyzcO7ngVW9P8m3VGF1BuBA444ARHNhhHwlSpK9Pp8f+VWrOI3udohR2TDXSNyB
PkXVKpyX0yd4HMVQQeX5NR9nAJjSWLQWra/a8fFdYk5VzZiyE5qTSpy6fhYVCXTIov/XXVUbNNuH
QinFxX5Vg5t/0qRO6L5v3AuvRAydUYXLD/EfNMjzD2ytyw5I0VMKj+brKhpxiO+MDlsHOc5vvLnE
rop0kv+CDD/bjuXnI2Zw7u7h+36S5nb6b27yPgxbZHNedgGn5zQ2Y6zyVSsLORxGCZayqOVEF7Ny
AuEhR4YYFgMJwMeCZ8urRhrSZfenjAUHi+jtbjCR9EGOOgIehpJubViJzIXAswhK9YAWYqmdNB99
nSq5PmTcdy9yG9d4R9Y5agb4k4MfYqdzU12xLUastiUpVXY/HvBG6aQvyJ2kHiVIjpzqwSwVdutH
D+RlF2lvtDPSci6gOQWcLwfJjnooitT8rRhV5D8wBiF4INTBb4R6qSt0ZJy4DGLDDz/A1/YNzlTF
9r3poFMvd737JdEEr3VUgT9jdP8iGB3uQHJV7cPQJPE9UNiZFlxM6zvWzNzEFV26VR2F8grBz5Ch
8mQeb1Tu6xd4OEfTlAi0FtQUsSt4W30PVflY3Hy6Hr6tS1s2cZ4DpeLr/1S6ZYaInAZlKb5qmgaM
Cv9B6luact1PRet+jwpObfbFEP8LL28c24ZoOgyQCBmPeM7zrjOG9Ah4wRo1uS0hdD6yV3E9w7lB
V3ew6LF03KRp22nXV+B/r66mUgd5AVSReshu5xvwt4C9QlKn1MKRAMiDoiTP+zBpYTWH5f3jwIsE
Fa6fJ8kmhEEdA9RiN5I41LonLYmocNKKaQpl83rXP3YIbKVsrk1ZhhX2czAZE2DS8spQQMukgBxS
BoKmiQtsoaenSsvTRmw1a0FUItBu/kIjYd3rJ1HCy/awBy1Zy0uEIVjRTtXHIFk40pSCe9PXqin6
NnAjVKSL3Vjbs21n4GSkzwVAQXNtsbdnqnbHf8l9USletA1f0MZciAufRdRxigVWD39dykIuqlAq
EBZBr4MCGAAEAXDIOzikTRz3Y485AYrZeVzfxnkMprWdXO4zqL74gGGQX+0yErFFlBDdP85NqwlU
2bcZU4UdxKEETvlsiSD3sCnxs9QgyUiaHhxV33DBszG+GD4iZ8aGNYb+uGKRaCgMqhMsA1Q3+d24
JJ9C7DdHDxJrEnNGgFyqale2/TBgTTWUmffpnLMcojy4Olw4iCkRnDizjgwGlHmMNq6Reo2P1mFO
53ifQ+BiPk3f67hRULpTwtqwRnONNXIrhpBhgftRf1LjXmT0hCjR6hd4Bv/DRv0vIosdXykkbUUc
nLiMS/XH5z2PsVyEGMu7jQ1YBnBSQZxPpIJbw9m6/OELSsSRJ/8m2rg9mhcW/Ap9dffkzS3EMmOw
CFeWj9wABTE9OOheNzcYKH2tSHx6FTCCGd0/FrUDibtDX5vbAlDxtVO5azdQCIHDv1L9mWKyJUgi
C+s4g5JzSNo1/yrGZkRwFRkVpoliaSiiiloyIC3DvfkBbUy8hrW/qm2jcItdb3yRxYWo7hsxkCu7
NQHKMNIzNs4WHfFLDwXwFN6WGDCu8xisxvexGp9tHTji/ouhplmP3RWywSPLxBkMVzpkdAWyCyHE
WlWuy7Jpv3YM0PXeb6zlIXWq+OENjFQ687wFJgz0PqMl8KhB+fRQZ8PG/zwFM4jYO8wxO3OV7npw
91U/WBXx5UT3jMBUP66WCgr/4yDXbfKIUVzdMz51v6cxcXbYOZmeBr8WUT2PIW9o8FmURCJFJ7gH
CNqNLS5rmuy3Hl8PlKvCUzj/qPvf8SmkgCYK8S6qxeMUa7n9fjp9KuE47Qf6lpF4nr3OAoizz79c
tTJiApUwBDSpamefw49Ox56MPVxaTNBpYiehkVAwZSDQb12FjfgajRpHIeEwIPyBECRO1JztCr+v
1yE9elPhAjSkRnduvH0XM4pCUePuqBWsX6xl6sVr3KPAmoWRZite88hWf+Yc29ylzJnRoAYddQs4
DO+6mcFSQIU2rHZK5dl9rYgWTzbF2mZuFhKPNwVUqhcObGX8Q7DLTYMviohenfmmnX5jA/iCdUH3
9FE+DndOoH1gxQ9RommpVkl800bUR0ah6D04UOZRXOUgTqIUZwIKENW2JAu+TUYimE/0o8//YZAk
yrXz8eg1aoC0IEyQb4nW23MdV6f8HkE9t4byGnujkhLvlVU5TWMsuMn5vcU4kFgjAHxp51BI2oZD
dHvvtxVL8ypHqoBHa6mLtWNLUHR5OFfkKgi6qAHi+3LeShYybbxZB+ffWvTimyGYdbI3VetNWRZH
upmytZeVQyomzW7QI9NbgF2N/YhRMyoDi1FtuzY65dRn3pPJtF8wtmnOnCK9IYFIdnk0fu/vBSUn
biak0iDw1J77yc5rUiV2JNRZ1Rq4+Xdg8EPQ+tq00x/kVuKpawd/wZ/vNMqZAQzKLPFgI3uPtQhw
/gopfA+9NEZDGPX8jzbnIRSsiP6vYQyiM+s4kGuaOMb0Rdi/ok8lhn9/8advod0sQ3vPynvZAlQS
8aVmuAjy+0Mx8gPpCmMYSTswmeYUWTB1IuWO35Z1tXW2VQNwguYvLSqafvtf8EoJxYblWDWeQNGi
xJwYe/G95HHKlD6DSIvC4lYnKwirmyNHBKwzubRUYvxH1d9iHpBw7NXFMX1sLrN5TW8RVjFiHkq/
1gLlrVfdvbFv/2+YypzvNOP7Dybq5Yb37GJGV3Ix51G8GXtc1OjIoi/gVJAyLxQMCXLBreX8o32H
B+MNPguY6lRcOGv4LbEF6LN9ui/xUqIEAxR+lDMLeKILVgvVIpwEUQMFJsBeo8nOHx9yOp1o2+1E
SBqhDYaimyzOvPE1quxWzFe310H8B+kGpN4vPwhO/OfkF0hIHnfX4FeYhXuY2bofhkple00d4ALG
jzc7gEhwjrrfjzCOKmOIipn+Z8Fp+p9LERmZz/UUtTtPWfDCy0U0GZIEyoGTWihmesurB+hqhmF4
SbbXRw2hkLKDktZGE+/CWKyEHj6ZRhIRpSu2fNBgk2L2oAhcM0QF4bDMYs6oTBt4qnvWURe/2opx
JOR78ZkZXuHlHT2T1Z3Og279C/xl+xJEMNp/Tn7sk26dzu1OwIusTQYxb7RP9XxnwjtKsIRbWep0
hs2zLZ4XZphXfU8eKfhI4g72ryjJXStX0IgQ6dtoVE+pIFFO7S+tcBJxGXRhm5INKbs06mF1fi2J
28Apnj4PQV3CTmKQu2VNl+F6IBjLocyVUBFTpSGU4nGstEgmHFAi0rolcEbhcpWVi4r/52wbewmE
sx81F+lUUQVBw5DZcFVhhwQTAMnk5c9lqi6QjqyeQK0+hjGPGH3qAouPt5NynoLNNxHggTi3MSF+
fAmLRkJD07Aa3BpANmwXgf+91fdV3JYw1ihcBzTrzHxY7ixn9/rwS7GIK8tDxLVx4YbSlEAzdw3H
SMXRrL6Y924DfzqaD1efueUznuZ+lg3K+bmX7yvNvy3Aul26AdVjBi53x8OkC9pgGmwnrHqRjuTb
n2B8UA5xCt5NfrX37YWjf7nCwbNnYAzGqisDW8PO4+vjJjRTrvkAAq5zwJR+I56r+nANDRg5Rdsq
inZRbGRZhdN8j3vbqdBpLn1iYXpxozWn7soEx7rDitDIokULXKR0+E/1kx97VtBmZf0WbUVDIApD
cGkun71mA+BJkV2RIKc048EMLYfzprpYSHYZvd3mGrp7FiWXZ9kqKLz+9xoHEudJMT8yB/egAu+B
Av4YRj07rj69q4f/CwKuvixxGBL5C8T0/CPnuB8I1ejXGgtWm685uecUzfJXUYjdh3ToS2OSOXVR
rEfKKSUJSl0cOHj0aExHzJYtRPsoKecbhjLvyliusWhFdIRfgHQNDFrnuhTEj5XwxeRuyyvoUeGS
RO/LAWgjaFXa2Wb5dzHAo+qpE7Nc7+4QxmT1FLEdTEqGuZsER8iUvQC2VrGj84aHRvP1YmzyPYRE
TeH5PpY/R80TOWExE6n+fBOoaYJ8zj9H14ekuBH+Pkb581zyDNIpQmXEOOvoY4p419uTJcxBKYVV
HyKL+QurC9PM/6nDrBjL+w3Bq+lr3vfhSp4Y76LmrIno7No8a3LXfNE5qAf9wZ/l4rex+Uotwj8O
/3/tPr6IPBi+tFmRQKwz2Dk5XDqO6EREMlvMNJ+QW4MpfWJL0B1dwKqhShjCpImKX6n0vE2qDh+P
JF5WhlcOBOejUwfZW7lpcgh/32d9Cs5vXKpLPb9i5c9gVb8288n5ntVk7zvd3XpO0b/OZR/dCMJc
95e+JMdn+Vrf5kY35AD64BNpV9PL/Xdseeff7yd7ws8qAREiL67mA17Y2RsOLwJj6p4r192wmunM
FesRJ8i21UEjBEkUma7WXTNZEbSytptlKElwunkdtfcXh+b0zMCwxPVeFujpqUmtHyrWBdDFSD77
Kps2XnprgazbqqwbM0DdNp5MldzFh/cnX5gjwZlXg/zLTeILEdEx8fkvhXnpox5hDI254q7USR7R
/+YeXAt3zCKlzLbJUW0koJony0ZOYmoLqTm97r2fRj+35J1Ir1sn57lSEuFdlt3q6kc9aBSSyl8+
p1d++kbTOfShl0Z8EHudp5pDRvvr/H2MonTPzPqiqW9JSg3SkSDh39ypufTzWDuXZfWwMNKHEhAi
cjiSPvd/DWnUCKjYBy2lbKW42q18wKtWAD5uMNRqeVdO+L81dAeFaCwWPSHMkG8yv0IcOhllEAsW
ykRo8wJWvbl0ldohUHy+PwsDlAmNVXrMezTd7QVhyUHECq8I7QT22nKSruXC95mczAc8qxd6a/2q
gAiDhLVg1TZ3TIJe/edSjeRR/dsG6E+lyHJ3X981AVFi9iyISB1SoaLYgf05tCLFt+I8yE4a6TrD
QjrKBY1oWM1br4FwnE4Z69Gld/2U6I72bC2e6vToyyiLzm+Rj9Q9ljA3RHUlFFJEatcXra4dX4li
/O38YqTmz558Wa7PuSjfsijiusWkvtinNA+J987vFzVjKto1aRLZGPZ8wRMbgmQ3Hu36v6Gqqrzo
E+BaMdZskWr6SMsVNbJAI9hfjYpgC1j5pTxfW0/BiIskg5xVIlcrkqxGAKnHB/lwr3zbQ6j0lE74
Dwny9PGh5gajBYja5PnWDW5B5YGT4XCBoyjsbSsnDgeSE8FtJL8u4MJ+ENPaX+pYtqwHm8Stl44n
d1WEiiqx7bxUKBXUuXcpCF98FFlWUsTv5ZE5rm9UNcqpvk9txFZn8RdBrknJ1XA1PW/oMSwHg/0U
TbE57RQXKsJCWPNT0Vk2TSzFX2tpvtxY+Ek7sjJlF3phsj9x9EBxaKEOuOd5iee5EM1YREcRcZEv
Yvf5dQngeSzIL+qBCqqU4F0Y6JCx6xNeGn0n/k4aLzDs+6KgSDslvmmeVouTcYMtZSzy7of89UUO
cqxivt1HFwpiLKpRbkk2lYMiaQ3IsIE4VRalgwhmiWcUZnUBXfvzmKWLqIHbtCvey3wMa1Ixvzki
Qz+LzJiihgGzPx9C/f4Cz6u9pYQA7/BQrFPxVRrx0ykpnfG+GdqX5KWYyW66JwEShlsH1KMWD+K3
QaBja7Qgaee3ivLeKU1NyLBy9y2Bs3vsFErc28ppQbODvgnTRTzXGqfnjHjAKc8RVUV9D7OIZPFG
RwoLwiw9xg9xILsnDoIuWE7+NlWvV0EE7j6xh4BWFBnAAZP85CCItwGCURjES1YkURQLh4+f6N/k
LUNxELYuOI/VRXGC67b8KMsalSFCKZ1sSGPAehjYEBUgp+bWD2y64KzdEakGJPRm+QRdvJvMgmTL
2lasLi+lbbPROnPKp7BswfciA5/AyAcvceh8scwcKlAKV0MeBQHgzlFfvRHn4Ksssb0KaKKL4rwM
uzCDqAg74ikBPPthCGfX2EzObnOTVbLLzeJqnzT8fjHea7SSM7Wp9zIognL7+kjIfveoZhYtnHLh
+NR7ip2NklHKdAnOPrfLApijSZ6STmEkG0RLnZ6EOWCpniaeChXlDlcUKnP2mbJJW/Q83PYwoL4P
sGE+eNs3CntJfd+KaguWoU/NLphEdeWPm5glY2SC4nmoaWQH0nt/PulPCQ8M6qmj4gDl55aGVCjh
p4ue4vy0ugPtb01zfdV5aDX48GF2ezpj3m53Gtm9MIoYnxv3rSBiHPYsOIWu3VTf0OUICGRhYwgF
UOTdrLVFE72pvtsaca8fMZELVK+bFoXujOBkbvVQ6GkFhzn83psJGrjX2bAq6WvWiXxKF4xfN2Mx
wRT/h3wP7hMeYR0eVTlahdTMzlQdJZjLpN+EiQDaRWKAEhjyOry2SqZaIYaRzBNUiXSiE2wjfPnD
dfUG+ycFpiCTXntk07zYu6SbW9/TRjyKef3ac6B6X8NLtg3j5aCnSg9UmWeGqs05y55LlMzTod/Y
rrdViI/UwKmpjtul+pEriPlF8m45zy9M5iKOLf/RawL+lxdThoPH0FNnTEvv388s10d/i9HQiZac
IiwSfp2tL/wqqmhbx4DQbINH7gIZDikBCI6KX+/Ul/Dg25emkcFRhdZxbFCwgrk8j6SpX5JDIOxv
RgQW/Rs3g4y74+0+FNkQ7FfAL5IFIKYLhaWzs9HN0jLblwOsdcruYfyVt47bjMJ/pnHwfSi2suD6
tJz4gU5wOR1M5GkhmHLw7d+wMIqA88eFgaT3KHyzHk/L74+nt3XXjVfy2UxwQXo/rEAkjeeFcp/w
nsJQiBkr4J7dWzEuTzhTpH7pfCQDv7B2rs5dJh89FsBhTgdBL6WJaNi7zYL1TAK4wvOd861c9yuZ
rNvilpnge/+Bfed03YL7L64ZUZ5EDiBBKIxhKFUo3hDZiC8bIAMOFixAFY11DY4PT716np1S4sGs
41HXPsqj255tpQHOPHofyhLV1S2jGpgreuvvaqQAh7rTXYB9Sc4cV3VV5fXHbZOM+dSGLA0jHmnZ
xKuJcskRHfdzvDfeeXZZbsNihVC0+qnz0fMBO6b8eEMQXRaXjlBeVCF4k3KOdKa1trBkc5DX59XZ
gk7gDL2PisnForgzAzR+job2pAqDqM1ivHD9uQfxZz+V9hb8gNcD0bCnlugS+IYk1iixdNbYLUWL
vAxFi1Xyb6QboqNSEkvw1gw3vjttloLaVOwOXlAI5JXf/VP0+si+BWx0YlB3YCMSx33grCro1FRf
XNS+cMs+zVkqB4yEcFKeyzw1YgJUUOymt+YzRj3jlmkFk44pURvf1bT/jtAwJEAt3EATWDWeEv4v
GoeGg/FXwQK6I9zhXLGTYB5xI3ruiNTbm3rimG2XmvpEIXdaMxg6MrFD+lJ3FrcP/saLpKM7mPzs
br1ewRtxglrNQNZcF+W/OW1OiQtxFlsnFS/q29jL6wZU839yii/ju+xpTbvhTFIWmD1Uu0lUj3Qj
XjzqkulGulznlvM85tCljHDI7zifX2UjO/6aa5UwlQANHn6S1LMhzaKXvNExYotyLPj/3C6EOd3g
r11tK5vXVFTR/Uo+uvGk4ZEBkQA6dlfkf5SW810PvcBqXLwrZqHIhTDmAFsHd/6ZYIRmPZ9vbavW
KE+N7NTtqRvnJ1S/O3cXupI5oL+qFaxCzXKenl6AJ2IoYfITKemuE1CA5ql7yR9XEMrc8OqYXWsV
mocSU3fcAg/2hkirPwQah0HlsieUMpXJDhPnfqsHoeJO1VZBoR7DMPiscCbHL2uZQgCawdDA3K+k
xQ8viwrtdF7Rio3bhKnGLBQCmG4Og6jQ5k9xGEKCC7lOjYudKqHyFOzOtTKv8lWqpm+eIi5bpYB3
myWW8d7AKRvTd+Ndrl1vocOQs5q6OU8apKbz5S0BLa2dpeTXB35iHywEf/VQErnXgMuNO5NvY4l1
XxIXf+KkP67sGgpkAiFMMRGTAu6GFDG4GNypZL5wg0v+qwYcE4YOQxb8raDgDhzxQKFke+COcsnB
GeV3cky5IiFNrpbfzhl93y6agp7ufkTDSQ4G6uwR66B7eJEBDvSyt1Y9/+MWBXRFWOyu8JsN5p3N
vp9TIdyJVBAQL7vKVqZjyw+i4xXyRB239kUqnO+UB3CWQLhGrt/SpygQZlPkZSU5r2A2Mfyu/DGD
Ib2z3kyD9Rr7VZplh+NzSb24nzbSUQLNs/NHz7YZtayxm4jSVtvA/9JXUIFWzJV/qv8vwJDyBKrs
e+MkmxqXCAjR5lneGP6qpjWmYMH1iVR35cryNwER9kP94f2Rd/WXmwAXEBB4ob3seMhY/pIIaQaQ
Us1LoFwMJgMdXfjOhZzHjFz8JkFrXWqSrQ+tzKKZVHW9DFNpaZaKstwBm4zpcwMRU3K/0Zqjs5/f
JlxCXYusIizPZyVLzpvUvbT4ZYqNmRNI59hBNoT8KsqfEsYDBAEVSgfBGeKCR5Ot8Cb84NfvV/Um
XDNsK+YP/RHVpBT6wdwfNRIl6Slmkvb1kWxCzSgaS8pQH7a6PO1ZBIoVUs+oy182sNRoPRSuSUYo
AEzQUCkFpc00YHDD869lXsHrku/OV6mcu7jGqZ/9gir7oF2lz38VPSei4aNjHjq3I7xxmssSSwgH
iK/ZMGo01b9SC4Y+OwRZBNHtWTquxU05Kvlf6N/QXZUfk3tEbSJxQpiOSrvoeVnLfbi9I6xgjxdP
PWckcwhG6X+t57rK9ollYDchWXyuAQJnLN0W+eV4C5S6BBv5xTdcwSGBN3i5n7j9FM1dmebO0kP8
M1kico0Gr62KgPB7d/rlBfYBIv2twkXV7+qjjlve9EtoV4uXFdl5trtokDvaydk9pU+oCVY7l6Ua
PLuXcyy/ZfgDVpov40H8U3ADzI25PVPsGuaJ3ABWe/7DAsPPPXJd1YjS3cnvE/2wXaMJpAmUine/
Q76mHb04JZ5N0XP+Cp8650mRvKK+XOA6ifuv7tnV0n+gSyT+PBsjBuu+J4tLVBOTo0A15iIDmhR8
aHFQD23j8CCsSDJjbon0uIDQcg2CF8lYCVlW1lbeFTKYjfmLraZzu9dAlQUBc2Q8NN/txVoQMXEU
324FVKQJecq8hFMBtWELHvJRZ5nra/tv7fZotnM0TFgp7eAfLRXA0Qk8cLw7ZfMEL9aIKDBgax3p
vjFC8KrfGPH86KYVkoRn2whdLLapXBQRT6hDAihFiABlbk/NG7CnENLJ/c5nDmr8aj0RDeOgxMEr
zXfjXR3zIxojS3DzRH5SZhMDHiofHVdLeeMKv8++ff0YBzmm0js8tpFXZUEO6hsRhDElY5YbhZk3
P9zW4pzelVDx4CK2UXcXX69M0SUwB66yUJj4/uvvL9NU4Wj5IakPoNhqHXc8Zz+zPLDag8DUIr3h
MpP9G7SXJsvmJpiazC0cJ0D7WphTF1XEPqwNU2mmQS/p1S9SWptQO+NyxBlHOwHQ5erTCCDXP4zB
vRphqKFw9AM5QXaeSiwqREOYxivXfmfyZG42Z3ynGT8kAm2QAdFjbOqhfAo2TGkdP+vfllrIek2Q
IikbWCe+qAdilWJR1koucZr3lX9ls65HBpK7VhfQEQ6xidP9J51MHbfVFRuY6PCMp9FYOEvFmbZF
5P5JRvUj+Ivg8Bpk5uDEhnpml5QTczgBC5oPsBAtgfOSBU1xvL2NnqESmqybRqhZsA1U1iI9EujR
ANPRQmBe9jgI1l9VMaa0pOeNsHldLVhqbA3kWtJKtNZt/2HCkE/WaRaGb0ztEHjvOLNiyeeYPO1h
PV+ce4t3lsQhHyh82diHJ3KbGFkwM+ooMfx+BRmsoxykaTr+eztDqWBKMt29W+kV0ayLCT6cU26N
L+GcGLhjKVW3gS2GcidB4sn6POz76qLWVNVF5K+VkMlcPO+7bqW5yITfNUFJ0ODgqd2OG9XD3+vh
4YDngPLRYHnO/XIZZPUV47xP5fDpsMNWpsEYfuzUFPZbMZWjxDrx1BEYl5fCm/ywQFjD1aaRwY1l
cHoE9cnD93GeaQgq7vpU7NvPcWRU41jmIU4m/YD0u8+7f+Af7RY+iNZpPkgC7B02VKrB4URPZ9cK
IyPwGgA9NxI7usBF6he7KWbKrBGaYCqfrU5ZwIOlIS/G3kWzoufMQCV26AzTbP9SyJKWIUsFEbM8
85KkjzGg+ucaaSC1nCj3507Ro0SquzkUHjTpHq3G69PQpgnitMRoWGhDf2JGjD9icW1Ot/XRC1hg
x0Al60bkGcVRekyNPz/a8xnP89LzLyF/3CgLcfcQmk3ODiKGYQwSCOf1Z46beuL4S1rLQU3797Qr
tSG2FQkF5L7g8KmnYmHaTxs4CYVX+iBsYDDVARozTxvTY43pmpVS94B3blz6xVRUCxaUAp0dNdVy
6HvGrSBTD7dwEW1ETegoJ1HKXOz6Sb9pWy5ENg8V70awRvnOuU0SEq5ZBQqc2B3aGoJYgA0u/Kuf
CrV5x7b3z05VGI8zSs+7brjf63E/YFhRfdXQLmoWjvt7U0mFev16fIlmmx2Z+GAQrEgZYfOR1ksP
igoZzB90bTnltjyvEedN/afAv5iJLUPEVc8LHabiGAau+g88C7Ko6rTwwFkL2uuvU2oqYPzw55h7
zVrHANur60oKmAvWQvC3EQ0rqkuVqzfAdcPsAItDdHhExVVoovk4OlQmZxIbVhJjOndOH1nYoGuv
2xibKKFFQLNXeFRDPUoalZm8n8tKUrEbEYJTzDFk70YvRhwrg/esooAZpy8iaOkdqadgk6/SCvUH
F1f8Ts0XhibOw7jm+AtWDq2lV5z3rw7VLDtnweRuYKaEhzACGfXOH8rzYmdUIo6mx6dA3yvHLMzx
lEEOl6dkRhzUyQpYhNwGLfO+4v57en3XBiahKl6iaSOjcV0ZgXoY5A5CNwrzmC6rvlHRu7pXhlxK
ytLpBDWlF0/+jhLAYsC4nldamOy8oGKr6NUBCNwKkVLTIymtsQkzTp4HzyQjTgD0MAnfgqwXezxE
lKvoqD21niGXlkLQb0PzSwu+/ML7FC1hHYclcC9v/hLhJQGKVd5bOecNJGgRdCwJ5o/g6hLTEmLk
Sf2LqYdJIicbqZ8Nfjl33Guds2Ns10SJVk3Vt1JiKEAtqhSh9LuGl9ggvwhT1ZSyD1bb5cYRQn05
RWR0oA5WnlCAQ7j0TWHY+SHVVaqrss0zlE2Z09UuFlNI6f9/wZVeWC6C/xrc8Rx7V5fya87vR44r
HObAVonjkfBhiIvfrZFahXs3C22aARTwiFoXwCAoPHpD2Xy2Ry+ri9+jY9+In0UsVB6kBp0l8Yvo
uzpVgsPEI2T8JPrwm2WII8dQfjlrQtV3/L2ax1vnfpaCyobjQKXIUzZ5sOxy1QB3kX1//hnL0cCZ
qc9AVjvNM08waFn+OmeR9ZXikE0zE0S0oz7bxVSicH4JX3D3aPnYDSXpAzzn9eD/1gLS7EPf3JG8
v24PYfhdPBAcFaI7LSnuzeppiEfSghptkFOBGGlTVmJYdygztDOSmES9lSTp2mbxhRCX3jIilpBf
USnk2COWGgr+Ojf1CtKDapVgomgrhZIgCbrNRKuSt92dQUtDlpn0wPmS1xJ7RrnGbSnlEQMB2l0l
Re8LA6Nd1bxxu5iWjs5j9Ee3UkGSJeg/hLFsRqWzKn3cyxMLJJmpKBQsk4aTs/8lMtxiTzrG/AFa
yVQwRJrUeGtpZI/XPksUbLFJ+JFqkpml4XR4UKDxL+rj/xiGj7Svxc7blc3+VuxmnUBmmMltTDyn
PyZHWT0GG9u13QOdTlX3swSUTvesULG0EVmKEtOq65tl+L3S9a4qV6l73nSwlmzKjAQvf2pA+1/S
NMbZy4mpUEUKnsI0e8vqsozPGFU5DLU0LHUTzlqLBaCTw3n8lfr6HPtdYfOaIotD/2bbkFfAk1h3
u7A7JDrvvPT7fMu2avHIfZ5zvp8n3uq+DkYmnJV4nd1+hZz/X9s6EH6TxGb92Tec6EQV/Nm2XOlZ
uraKcO5WWrXJTHr9LP8acp1Y7Q+ycp6Rh9wB2yaSnLCEoKU9d0BGRQDg05alobBonyppjhDyYZty
XDHFNMOGLd4sqgT0laUC6jrR4FT6uRuMdEPOcg7sy6RGBgZDhcytEFnZM5POO+bGKXS6RLTvVEC5
oN1B5aAMd87wEyApKFKXaT+DQbX3tHtjz+ykquFoDiIVd4DIp+a1dZwLlyxm8ImtyQ5r/ktZ9o8Q
2DfqhIUGeMCyUhQDRwf16KwmnkDYMS6P9IxvCsKiAxymdJcs4fc7KKYDxPwaEjbAIXA7IUrbTOue
Zxji1vks1/vJ2qTX+kzMWAUbV5eOL+l2ZjyM9C3/PJ6U21j6e2HGE2TUelGRZVZ2thHSPWDMrjbB
HX0Nmep2c5ECWzwslUdlYTCVkb5jMkTLh2XhQFr2e5kTxcDpPSuB530OpWcYnvR22sn3mB7U0Neo
64j5Dwil0liTbgCUUZUh3kafI2xRRwDVYqABuTnYe5WZD4EIyL7QJ/x0Lgmyb8flerTNRl90SRF5
gxoraijdGTazmzV0zxJh6SPrOfzPdt7Q9LZx6D5MvjSIhfO8tLktiEx4PxBsQb/oGQFqyI7n+c8l
pDl4mSioXXQvJmEcMKF2GNofjznwPpw1H36zJ6BYSgqbGU9gVodT9yGOUVloebKQKyfQoLZ4ef7C
RiO+pEceg7KES9A6cypG+ZSgySoOjRUsjZeXFUT5WdkKoN4DGImOTkKtLmIsoiH/bix2W0GgPWhj
jHK6kgbru0nXEwKbluXlTisHDdc6TMRuqbA+pvmAwiWmaBrqOFDx6JqQpcVuJXY/8b0lV1qGZvBb
r0JrxCnS6rvTQ/Q//VUU1KkmgM5SzWs8HDbx1+458a7bm4v8sbHnJs5QgDPE3vNVh6Terdiv2Dw2
9N3bXYVcZKzTqm9s7P3agyXM3gLRD18SBIy2O7Qsm2dNY8vz1Eg/G03vU4z/P2wuHFcAAPFT6VIJ
NQx9HJz7WZG+Y6RSh+UD7qzRg9su93D+YABIbVW9T73uUAiMHrfsJ+alc2335hSBarq9HDRE+GSG
/g8KaUCYIz6qOxf7rhIx4zSh1CRlM/aAO3loLGf0zF3lquvE1H16l88ze7E/sxOl1WLN5UgingjP
bAFpweTwjH9kvAGoT0eZ4mF4m0oMxLvdhHMIEPo0c3JqNs2GXjK8uaJMrxhPdD1Ja61b9oYoxNr+
mJ8DrNqcRGEJP97JM+c5JUcVnzLrCUaRrtzrugLxxaitFIjZ1eTj6kryBL/jGEKxz4LlwJc5vGyx
gP2QLiYhzUPqYKapoWnl9p046KsNb+un4xsvyoNaKSMUAFlg7X6j09+iLv14SyZyH1y3hBUh+Lls
FWSol0ncNslLpsdclRL7pt6bZ7A9BgnPk9F/j3CC9yccivl5HsFXGXe9WlWSsrCAv/bjm1hXP+Ut
qxEcMYj+wgespEO4UqmNN1AD16WyDYZBXfhFS+Udwa38AB+8TO02rARNxjcJ2SuSiy2kopspxh1B
ZkW2Ao8HytOZ9r4ZhpO3iNtvz+faTZnG9HuCOhB2MV9JGuFraHEx+UiCYsdFUgxPItrVJFIARwMs
+GhDageUPajYLJQ54b4JXGOTpHMfdNnN2wSPqwe7gfyH/zsE9dbgAh0iR2jf2hczrl+vcVuQlzzL
5s1Clh5YqJt3pNeArJELRa/kb3cBMfuzauhQpgNYnEeDvZjdiFaoym54DhtggWwsAqT7+OFgdgPa
E6tkXZw6Hr4PqcoRljOOGXl3ERpdokKd2TEB6XdHxXi57wxXLax4Xk2jnMTgWJk/s9O4s/SXB+8p
VRhzW2Ve/nZYTP7deGgx4npkdSkmTCDUOdj7nzsHzMKTSmqM6HtCxhw1FeavJQjDWTqK3hUUYkhE
f1bzrlUEMcQYOoBNgp/JCbHpJrtyXe6703mhiFL4whiezE4IAXZZZE9bUwDKYMKhJ1tk2oTSQ/mk
kAMawWyDhtO4s+U85WrVv0hBeT6uXqzeIlnukZIYABOBqYor2pOx7Lnd3j83ybtIlGI7P8kPK8kn
wIDuHhNchUc6oq4BWBEyP0kjH0zPQZEJG1rQwRaX2IdtQ4epTB+4Cy1AQ5pHmdhFj3NjbknsiDIR
hPwFHJw/7IsyqUNqaSdl12/6HrKeX5m0sgxMFkDT28aGmnaH8lfqssYIFlrWJ9NvzNwC+I6jQdzs
M4ZJ3pOqDRL+XAMnUwidxw09mfpfUGanLgp188ypqaTTOD0Ombc/5njj1DXo3rYUYmz/k7E8j1/K
4cngtwoLUXS6NdA7NIfIygKGzG4hg4VVXO9sm1mEO0igHgC5SMspK+h9N0IY0z6KufpsInmA11J+
1PWm4yIGMZMBIVS2dquUBOR//SOjcANCsZlU2srd7YMqq6mtzZFVQIh6eAgJ75lfisKWfx3JoUX3
iZM5W12eMaGw3/ceIWE4LqlVJjcBaXkgraJo1HcbRmHbUsegmdi1sOorJAh97A1U6vugfCEDbX7G
bZIj7I+8kl6vlxCqtDQl6lgTdXr0caWcTXOqa6eyo6WVAGTm2WEBSnHhHXJGR7Ewske5X8knSAJx
iVpuWYwELH2ufMdjyyNspsq+ijrAe9RVq8EKbhUmWFf/CgxRzqGj+bJl7U782D1SZphrrZdzUhLi
EkeMPNzAYEtanm6iM40EdR/D9gO3ES3bUunbDKJG3GsVEnO9oIQdAC2+kMnuSNygTjbEzdmip3Ts
qa8LNOkKaPjTVwcn5hNXRe6gCe8pT6ZNW8xpRgNTpy/KwNSoJ7ccm6O+gqCqRDf679LVxeXXAVA0
ISkJh2vMwb+0rZN9pWGOJLSqGtPl2nv/DXAqciJNbj4OpYgGjs8yp9nQ3wuP87ReE8wvdBa/GV4K
RtgcEOH/Yn8jbQQoPWoEbAr8pQErvBHQP6gKHjnjze5Ggs5H99t0Xg3h/HOrjafAegReGulBEPyB
0Y7YTJ3nIXCJ6Ex3uBFe9cRvbpu09jRY7Fa+pwGnQ7p8Jvppz/0G4gOiwpOt+6Alr45vP58mqI7r
Zml81kHlSoCr1eB+c3rqhc1LI0+znkSnfvJFhQrPjnVMnJS+rGh4JYCOQvMvW0Sr8XuJyIdajZHa
Mb/hELhChoqvHaGPIAbM/61cnjs1ii+EuIvDjlRXPR1jOOLAF8y9WeTPHjRw9IsYIrvsIFIc7YfQ
9KEccem35a0y85ZpxxCt8R7XNwjfxXZu6C04bTpzgZDpjc8iPVLKWJH610AiuoXnK/3MEXA1OBrk
Nh/yGm89xQL5l6Wcc/PR7EQiep7b5/Zkz+jfnKKxPl93ctA2m0QBwOvkcV67LoNWtj29YAd4kjdD
1JxUb2z+zpD9xz6CcVFB/aE1pT0gpg9Oe5ALRniuEqPveHQQsSlZjUjkAhAizITQp7TYpYVd/JIC
KKcB9TwBisOkFSj7rWKSTSxeDg/dutXSm9rdxrqQOR8dXzxudWTqJ7EU6sPNGOMqPDWpcRs+P4Ga
JWq46DBuqwPtjqGZaWqVcGHbp7DSbtnXnfRNVF29XJKZ5CzXgckyIvtlUaswIjtj3DB5yQwBfrRL
P4nXOVhVb6gcZvJ4TWXrHOIJCiOsTtMfyWP1tleukFpEY15Iq3ho0ywc4Qfpk9THiKTnHgeoaNzV
JBZ1XhRmKm7A7n3xrsGoNk3rYIx2HajBl2u8CZCFUIPFpd1xhHOsZewTsRzX9bcV+PuO/eG3hz5G
CBY3bgQenU1jWWRTHfWOPf1+s2i3j+WBbsknSPumkQ9hb3QkoTeAaNgBemWf8Nl5cWANenaAF3St
Sl4pKnme1zTRV+G9mQQGMdZpiINGc9wxmclyNqzcC7/0a0NIWLqUzR7qfCtBcT/VNtwOyncKHbmz
UJiGA+HleR4sgon/6AOTzi0x4p/lYmWHgaIE4KflhZ0k+ubijyrfIylHEQuQqAH9DF8o92bFP5zd
KY6mvfJtgHynmeK8hw7Rjq+48d9YuxTlPIOmSDuFsH4WOPl9vuPPSO1fEhIRSqAdQLKaUlQEENYK
JbemggTFMvxZI8MdiGlKs9SexF9tXQKG1uvEpZh5bdy6bDHUQuOf6L4JxHM5INtQReEHvwKbGYGs
XnUjMgbV/telve3LWSCyy9Bod4VJ9jrpE64waQ57yZl/ENzh5NDGSYWFD7W6gz0CoJQqgCYvCigK
y7Lmf+4qxRSnXMD5kDRWlUw9lVKR2qq1cH70mm8pK/7YnbOkSsKnhAxNh5kLg2BV018b05318liv
LzW5q7cctIaKeT3wCJg7fxsCm56hzPnZijFSWlp9RkZUhANdUWIclvZCS5X697wmEI1sb25h/Ku6
/A9B5NNxS/zjMw8uYe5Q88FDEz9fhElSjaIlWNNDzoi7AfQwHM0UrgkYH5wGqcTPtL4640qEsftk
6jv2va9XRCQbXLr0WH3VYPrpFUqZKZTWpRYiQ6JlUi9FppRmQtWIZ91kNuXHvEgP1AY+3RP2TUWC
3STBi+M+MlPjR0OzGqGZCzUiCaH8VTEZKbS2SiXuHVzG+rkRkN71bUDdYZ+83kOQiHAKqx4uU3T9
6pD/4/2UIwURiWyFuT4jYzNnFQ8NR4cndbX3Pa7BZAvgQcR4xMbwPnM1nxRQxMzygouw6LElG2sE
S5uM53+eAxKtKCg9jOoXmDwZGjlUBxDb2KuXBZ5Km35cEm9zfE5lZMY7TKfvykh4kCUMFBCKOGa8
ZFCqqDou3H6cicrh07CtYJipmDT46fHWxIU6+zBCHB4sGX4DisGutzEURTzsau/dZ/8wA8yN1Hny
ZcITmeaJaYjBHNmmF9s/+TzPAn4grHdahwiePwbpfw0hTWX9IHFYTE7gPltZ8WmjEzEOqTz08+eh
9YhM1GFGvWAryM3Z2jbawCw5TLYf8f+npkYe/TkL7es26kX3fQhdW4awpaS4R89zQJDGaea1GQx0
GaS6CdRjhMAnRclJvkYnh/umO+gQa+6r1dMwS+NJ5d9euBvMGX44k5DPHwDBxfv8RQodaoYheHHh
cPqjh2FUCwVsA1T8/tiLGc0pyIouRIkhgOdJcU5/RRpQg3TmaYuVkoae7FbJikjjWTjDIElMnNMr
43uRzrvSlk6Y5pxoH0uNZCn4ZZ8zZXoP6f/uWKvQpBuW27IKhrzAvGmYH6l23Ul5s5DuCPzzPnMk
8V5tycsj9UCCpuz2RbhFkG4iY0bSO/XFXJlPwQyqIpSp4tgY+eF8AsBqsXZ1jCbQPibJnQ0hmd5o
mVsAbkJbr4O2hRj51xeGJYwufQfyCCHoniQepZtHNRsfajw2uHAmcGfm9algOTzGXPtyNP8iWc1Z
Lr5xuo73vfcnO+hhhXvc+6Fj1PpZRfSSSOM1QmbVi8KaQ3pSwWju54snoXq+Xd1+/JiECgddCaO7
UEPLCVs+QF1pJ5EEJgsuBhOyOpaWOsfxPsN2Gj8DQzY5inPBqps3/RMTrn6ozNxUR2I458R3Ix83
BU1nipzH9UrsA9F55Ij85cpkqBAwr7gR1T8ApFTpI1V088IAJwJyc1Dhf8AdEjegfcZ7HA6QH0Js
Z45vaS9TDN01g8yhIx2KZ8K877MmSYir02bi4dK7KUoxzmRWDHiPu2NfRBVYWY4rlsnokofsy2Vk
uTVx21geAy8co3UgJqcx6lYUOqbVoXhADkaAhMzF2zChcsBWatnbSOhLFASTaSwvBNQi5Dds1rtN
AaZz4O95uQmAz5Nf+ZapdeJFIrB3/9wen3NWus/aRbwpAm1NWdmGnczesjEdU7d3lVRA5GVg2hfs
EjADJQnWYebEVqe80ZJYBRsLd7z7XR6nezO8yGztsTIDZVdj9t2M4e6w0r5W+rzwiWjgsUATTenI
83Qrr8mVZbEa2snP7KQ8axZt9Sm8YeWO0biOfLxRFvcVWwKVPnoLL7fvZcSL8zcIjqyIlEtJrHjs
cBKNFBhzys4Xh15BphVF55J4tpBIC3tN1bQsO4cPV8mTpY5BNs3e1+UecEkDCt7iHx6/xGgLUzxo
FVieWXvEIElKO1KmBW61MW6UsIvbHV9+eGAHy5I16/CKPQkuEEtqgiq9ywY5XPBiA1UpUPaKJfTF
y7Nt6sIAGnOgxExQLtiTgj1xYOqhw3xGBlZqiPY4F+x2RlmGggwSE9MorpsXZfZd2ASf/5RJZ9XS
KMjJuwK5xNRx8bpURWK3iL4KA/hvszzAIt6I+iFKbI//xplusfVwMFU90igF0SZ9dh+krSaaex97
LVRgXA8QafC7kQQAKpAHnnCHDB4ayE2x6eOMF71IPV361ikc4GVUfVcmwSpvNaGt8DdTYB0+uug0
w+gpfWuEJC8+oSpPBQorg1m22n5/LGwJMzzqfdNDSLp+1S41RICKt/xarjQjcd/Ptix6N2cVy1nV
XetgIzT6+s35jKdXA3C5OL0c2CQP0oXfP4n27BMI9yrTVUtDFmPT1Ol3idY53NiCFYJg2oSd8gOa
zRYDwI3o3lhq1095b597YIdsEExk9YgUHlx4KEigBwoPdKiS+xjzDx5j1FeEUiTtarfa79ewHrM/
3s7hLXR5nyFUuSxAE8eD6aKhAOlpmlv6QItLZczDiqit8eFJSOIxNPrhujslOTfba7aPhbzKwtKu
x3RwuS70N4cmkK1RNXPakz0/wUSyDyvDNAaW/jZ7ocbi3dsWzd0d8QNzEk9CJgfgdffssgGfAi07
Q2zMtVqrmL7f58m4oSI3d3dRs3nHw3FhM360X7CiFvhjoUbizyTLi3T69rzY4DljD4tumCVQGRJI
C8GQGNY9OtaFHGfKwgoVxIeDq+PdivkoCy+33iHnIsK/bxw0tYhnFJFgHbEUlZYziWpVmM1iMwuG
Ra/87WyH8QyOxiaBQ7Qc8ssy0ekwTtydOI6uLsbSWjqa13yA/isAMTizaMJN+/2lkO9ptxHZixRW
6yitct8FGPTT0mHUSuyTlvgKEYsP/yoeYelqED46otdSqIbwHaCYmDKK9E1nsp7MhGoZsLRoZiV7
TgO3SwVueVn2gGSzp11+EvCdQUBjcoMRC3CMQevR/qVzsvbtbo9tu+sdVwZk/WRk0qB6R2cNJLAi
3JTmEJregKg7BR1A+9RO/90FMota3WMfrpe9VOq2Pp8MDBh9eK86ZIdE1RVcen54kP+kvoyKrHRc
FSbnK3jQO4MQklElmoE3SIrncrRbp1+jDsXRIFwaynDsdUbXWpIawsWRFyI4zeZ5XPoaqN9/56fC
kcFZkOyc2YB39KY3t2gRaG83+f/suusuVdswCc9gNAlh9zG1SnQnBnhojSiwTuo3ogGed/8wH8ZQ
G5YBt7i9xKxOqO9SyNMtH+dvRIIzueO8tLPt8UkX9GVnhSRUIAVIgs5Ae6tg+rxDqUF9lgIHRgCG
C+Z8l1ydVKews4Tc2/GyA07TtsPify09DQF3tTJKTvFX+2OJExv7CG6KlBaY/37dDD0m29l9w97G
lrw2cSbi1VEm4Rzunt//fPodw5x+7KFIYCRa4u1Hw0xZajYW9LnMlqK4/OecvdflKBM0SCS4PFgz
kCCKU/xIKdQwFRCRug7+FdnJqyUs9x/72kZNI9eIqsxD4vvNMIhhLsqwa6AJ6yfGQWlAGacJQcah
5ja5qB8j9BqOf1D5Vt4hxsNrdCkTePTTfhQYdKj/DPXU5lL55HYm3uVWjtVUWiNrL/dQAb6lWF5r
DuywS+EBxY/qdS9iOY+uv/LXi4Rq9EsvJp9U9nfEO38IWXNgfAFYUd2qPy+N9fzqIcw61QUBCv0Y
ZneIFQY84rK36Xn796D/dTimYC0aYw1uohGKl1tJKKahmew9JNX6UZkPcaZXAV3zjn0fl/JR+r2k
ySGNwlNzZ4w0th8fbC44MTNh3e59+qjAeOEkpvlTbEmB261EtlI2Iqpa3k7rQ67ZNstUKNhJtzws
AoBQB9n/uV1PlENOnarPzeP7H7P9I9SX5qpcxjJX35Eq3RRBJIMRlwJrCo5TIfuv+c0YdkbfcAs2
NEo3jdfuRzHOp/OPNVgVkIeiEh8vAAT6XzyXYgKtvTKmuPbupSphZBrfEzP/nWvoXTnsZDMLdL7e
SYlLIFNGU0/hnCQOaYUf85DE3LtA5K30Xf8ruhwTAj5EaXLWpuUmYHm72UHXFe2YykWOEXt/G3S/
p82TasaGcDXEkaS5SwUlWAPK4XSFYjb2jgWxiyDf/32VpJnMznx0tOFb3OScT2AlFcDh+1u39HBI
hRIyRp3xkefkIKZM9iHzzFGn7xrfMiEWdGMYZJPcPVV5bFk3G6rUtxFmR2z24gZQ0o8uvSPVMumn
GQeAGN30SzaXPoT6ZWYoF/wbh37/Z6qOCmBN32qyJlZ3E4x+6D0M9F5rn2Xlhr5WB22KNGJk+3Sk
HovZAKYkt/4ZrBGQ1AJxn7BRTWh62PkEIC/YCs59VsKCSwJcG13DXsSgzrygGLeKj/f1UZF3Ggy4
GoOO7M7uXIhqLyJ+tHEXkRsrhZzaf8fknqMKM/vnHWpQ7M01oDz4vAiDGaJhaIo9Qxvtncu5ZY0H
YDLAO5Hf7TRM9lKXc5KO4G8DgB8v5dxWdJnOvWEr3CD8oUSDfl5Lb/iDAOWZcJUafHH4fWmBsSmf
jvi+ATh4REXdWjp58euY8YyXtxNVr4c7OWUEYglFlLJomuV7gGhQ9TjveNtWjbVk/j/FCoJjlwvG
HHsp7J6nVviZTHrxpKhkpypsKPCpIOYaDhmDq8GRvviPvyqCLQkUweUg4dZ2NZRFLh1E9Se3TCys
KWttbzw/rU/nWYs1Dh5stUdZB77CrN6h2ijcW5x53TnpvuJJijYUSHEgIIyYitIGY4Tksw2clWdl
3XevbKyOBU41PA/o8I3gisbdCvL5loUBJG7c4u0k36CO4xQxRiOquODod4YDouicOKsJmFp8cYNK
Z+B47GaT7cE9aG1ZHbRaUydic5wmBliVBN1tczVgfHzTJQ4bgfjEvLU9XarSuvr5Bo02BNK+B7e9
eajeKdgcRhQkT7A/f7k6vKpvl7gMThLdSPASJvUorPWoFUau8vQxSSIffGXdff9cO4Wxb5ye8Tqh
RlmO1gqYa34qSEo/b48w/WPAdAhQCyr89OZNQx+Ou2vyLBMxuj5R4T9nVejn3Sp16SBr6bbqkZgG
WrGjgblFCRUWQ+k+u8/HSeiT2OM8olf0ArLVxSiLPuAgOwOrV/+xvdmWllw1CjvVbLpvp6VwAzk5
4tzcQfAh1zhc24oe+kTFUr0CWTOyrwWFTQzGZwwcIgwNZHLs33FbLIPfk0b+9/hjEl9jCeYRfwJ1
b4JunayFPoU6nFpPO+ZfeKTPkiPA7JFd7XnmQHsxL0yPKnJTHYxUXXhWiOzWO9Mdx5odeUQ56rbS
lLKV+DRvhWjfs09KkdZ8xi89XXAKj6y53VXyBgBenZ9AlclXSOyT2d/Le7loe1IkKvEGxvutCh7m
lPyjkBzZ7pk7z1/RPSOzlpw1Tsf33VwFMG3Y2R33nzxnSV/KpjV8DsO/VkYepZCS36g2dgNlQtEf
GeniZ5BV0Mi4pN+pBYSAWog2t+P4DTCc9ZA5URw5PMmT8THSyE3gwG7nnxgjR2FxqMgEUWlT2woM
GeXbUsDH9ggKH3XWZjF/lPtTNmJIOeEnh14wS7yHYHbOe5/nBLlrC3pf9uELFkzNV9zEbkia3Odg
ZaEXCWnPsEoLQfrMM4fuCUj68TFsGM+JpQTMPPt0p1uYh1ycKWrlf1KMAExOg8pcbW2uVl8QdzP/
HCQuLEmhuQqOdg/qWbwHZ7rh+60dCjThUocPwUgPRJpWXfrcwy+qVb9y0Ks0VHobaa+tvm2EmbQx
ZpRwmFgswrJsKHRYwAzyAtRiFnvbM9gozvQpfmkK4XzZq33qgGgvQKIpd52+aRYoSgZ8s8brmkUg
SMN+4PjA6UtB8lTXCwHDsSCN4C3nyk6tb7rq6vaDQH+n56ZoVoYNouzCmKKkt5M8D1r1AgxnSP5q
RYGO0ZlISdly5t/My79On2nIUpaeqPcaOT3LP+X57HYtH33Dduj/adQ6c60nL+tnyGAyG58lKUm3
PMQ+yfs74GimlFGTmklUNkr7ao5TcBxh8FZnMS0NPoHiF3hrfVz0GZ33FRwAtJyoyRWcMFh7cjGE
m/eIFrvsWA549QhDGFw4nSXsFDtOKAmsFQC0/0F/wDNUwgUdsKlYHimOCj7zaPgikBfRQ6wmlsTR
3s3A8wHk+XcqThwHrRvnMOkqQJupBh3BlEOOR+hCc7k2r7So7xDdsrglz9sE/FW89PvUcqhIIynD
4vcwd7HuSbnvgX25rpOtX/Fz4Hg9sBTrvXzxo8kj9jRYGwUt/OoGtcm06ofqLlmxx70KcNUWap5y
252lmwXdQAF2pduQFDtCCSuUjllMdzXmTvjyS4l5LwILKEv9B028YmpkX9PNsq0C0FfyigviSifd
HPwm2+edmh006jsfNdQmnP5y8KaDECuZ4Fj5s1UnTNrRkU7M4oXF8cpnZC9b7rbQ3QdI4Cz+Ilhs
F6zLz5KBshmUscWaabukW4Tu4hmNe4d0VmJws6nkDyQfzUMs5BenVy0tUaOCpg+sLGA3HpYdlp6/
cB8uPnQ1vTKz9GGo4PkNcNa3GM8DXTkVVejZk5wrTk2y9KVRGI1CIfPQzv1/xUEPY4o7YuHrRaRp
U20yZlxF+FC49Za+WPH8ar8Jhl45n3/slCIeGDIYHA8cWKzx+ngI9KmecbifDiHsmEwZ7c9FR8JM
G+UqHSI6U2sGqPRJ+jEM7Ob0dLafcN6E/JYGx51V7wq1LMHBaiS0fxJ3vy1frAWkkH2AIAymug/S
tjHjb9ZYJ8xV71hKWNbgxssg1xzEvZxkVOpRaO2y9bwKLN0g0dm12TSw2vUeACMIygwkXPNqFGC+
ADTf6DJloK5PCakWBPICXj79cTqlwNDqe3ng8m0SLPBPLyCSFMalaz3xBZWA6yj3V3XIuB/GDVhd
q2DeOR4VR5EbuDNfHr3fT5vcjxFjTJh/6N00kWI6EBlL6WJVTbBpk+JcnqHyxIKIonKkXdm7BYoC
TBT188a8HgpOAs6/VU6WljYfwImASX3PZOGz39mDhVAvmFUio/EsD0SKFGwGhCGxC1jZgfisRf3y
a+z8bZGUI+sJQkhgakVB/GcF90IMcfkSJc/BsPQhnUAcwEgfkjJG33bP3JX5QZ7PAjcNX8FqZSkf
s/iY163SQF1oz5PJV7TeVFT5PyKE9mAS/iEaUBp5bxCsot9WrKt29fEI4iL/LEQSbfQxMpebIINq
PKBBwEJ1OWrvUWoPtzikrTxAHIJfAMAs2xlW9DHKiQRn+cXlNJi8UMPqE9fklNlkZpJPTZU1ch48
j0wq9sHtoY+ypBLvdgFyMkkb2Dte5wTW69qIu16qtGDr92l66bbjK4RirgYtpa145rqWLZ6nx8/m
0A0bWIfUTA3WsDOI9WMWvmzaf27/6xH2Ecdpg6ta3pdlnui//l7agn277T3BGSVM98f6fIqKosiP
UJnH+KRSnei5BBnr9i9b6k6/6N9mLtdrQ3f3MrHSTgiOpRVta4neo29BnsNJ5s3XoHOa4lbQfkyA
IJBUgW1phg3pDU9L1rRfvrdAcbiGIGEMBKoi1EMNpRmCQN2ZslHFsHlZThghMHhqKS7YLHOZ6jBi
QRSvyAsi0GVF7ZmE5FF1mQo2e1PUXjgZGxZjPXEhrs+kZVzlia+MhGdbmBAHMx9e0PqEqVlTX4MZ
J8aWFuAAAe6kmciDhPZrhWkfLmBIBzw0q648vKqTL68F3TG9mZmJAbvojYdU724Wo8Af+s+HrgAp
j2b0OzeA1p4jtKL30XeNC1S9z1/hi7urGm+2GxeLAtmDlZlz1BY2nk2NpF6r9pLxSRMfD/40ERYF
A1HQs3dK70dfOoissfIlleFQcwh6AG/fMz4Hr1yQXojXSXzlwt+w/T0y38XTKWKqRKWHpxj5/HkA
7FIaXxauLxc/UvkRo33pPNLj3gs4hZQ+pSMKelfhevFtJBt7Um/b9ZMxcNg+nQfE264lnDYeh+LD
U0nt6J2rx0eIeK6qumzlnD8j8+YPH7xd+EKqCRdcpkFPIVULOO3LhuplQeryqfbJU3ocRAxlQTkI
2seuXROfar2ToQED6lG2w9IMrUIP/92cTQOz/M2JpWncl3QOjrxcFkA1xw8+NjQWvr5opAUhiyPa
4SAjK4rsCnwcU46vYVI/yAS1dQXeDv7kqrBV88IDI9pw/OtIjMP1EpPd3w4T08WkYTR/Qq6no55K
356MuwozCApDaqIhJFCx5l4fzkqSCCY7huy29y4YyKc41rgMPAcaQ+7ri2DUbGAAaL7kCC7WGamC
r3/yM7/XiSudKoGk5x6yyWUmbGXiOsshBLrJfCyESoaXm588RIPJHHd7peaa1C0V8fRQRaGQPY0R
LIsgFzRuP7rhMDQUddLiYhvWi/I1OZA+ZrqA4BPUT2NMzuA1enK3F32L7Zvy2ZlU2OUoNp/XjgV5
PfFb+5byb5HsRJpZreaVWjtyYWOzyXD4sNBcs7EDH2vPnEh649b3LtuC+TDjOTiVI3TUpIAcWklJ
COT0SWtL81JGshU+VjsAIDA7yjrkkysR7L0ONKAYSkVhUXQVtpP2zP3Fk8Jq4NKiY32jFhO9unUT
UhqQgUxIhRfTsfNXD4wmtnlooqqIiaPRX1SpacnJzi36iEh5Lj13LbluzrWT1kSnVmpy/Pp6jCzQ
NMGcLncRiO/ypO8phqZrh7VOC/ao8FDEjd49CUVP45lZU1k2q7dsEr6IKV9v0mArsJplgw4Ga7za
1kYLeeof9uTMjr3qxUb0VUWg3R8BREF3rO/WA8kesOKGloUNiG8HTRbE84K1YeJ8dbu+scnR9ApV
XJnxKj6oCk073V6+coKpsAF7JTBw0W7Y7oefCAuS1J6DMzP+FE3gA6d2FaHXnwKVR0ca4EzPa1fl
hg+rUdJeDF6kJ/2BKskU8EVXtHejeZqR/BXQVsvQ1+s1ugmtYdXZFPc6pssKUKJ5ajuwakg37oWr
4yTrYRvL+9vuLykqwVoUh9WV2fOlNX+tQ4hTtylA5BTrsKwwCu0aM9EwFwLVzrisDc0oDnXTW+7c
lpkOrUGcmg6nGuIcT0cekotEG8FawBjgs9xfosUYTdbDLUNnTONsDgQkOV9z85SjAOVHnaqY5Qu8
UCNfQRebDoLR/0LGPDu4r0ld2p6gr0/5kK1CY9aVYLb9e29CeFwjp5dryLXwJLP+q9ELctinJIwJ
RQ0Y3YVBwwTVhToVmLq4pnh4n/nkV9md6SSB3JOr8LahMfQbM5l4/SlQbIUTlD1oqcFrEmipxj2v
mm9pwBPQgtZJT5AuXyiZYvjZnr0Sh6iZ6Bwj82xy7zz3r+rQfDaQ9qS+xbDJHlzACGCkv83vjK8M
KnIm58d6Et4kwsttGT+xcHdKxbuV/rZJ+gKVdznekOHIJoA0QZK+NEhEBAosK0HbSItAdzpySmin
gE/ydccu6WPzNY2REVpuBM0pQfR/NdHDLHvARQiwYybe79KThwAdb8CKij/ytUQrqcoNuYQR1/t9
KwYB3RKKnBMSF6bYARhQus7g0TYq17nEvvTNUOXWdWuEnODV781QkLkFp67vHJV5O38JB3+DVWV/
/GUe9rvV7TivuVhs6/zObBUjBWHHXGRmv9q+STtRA9cyyrFkLYEhCsT9Deb3JHw5lRC+/tXUeGCH
jLYIQR6QbCzwmYlk13Gl+tZZ73h977579pWH4HclL8yDcTnHv50waXkE2B/Y8AhNgoRt8J9VNpNk
4BYo00z+VG3YhWWaRlyLJqhYUTPqEzJEDqmtu+IOrKGACJbV7ugrR60tOwKPaN4hJPqZYwjzAdQu
zqCsSACUoOwS+YKwbnjC0mVEX0ugFBh+oMHIFfPFsxODtadywb591w37L8K4TOZ0d/nwBehmqhzk
PCgPzscCO9ml0iI2pwTMQUu/EtBCr197x855Oh7wu7xodZ9JjBHZLqSdv+s/WMaqNviC4jdLmChs
JxEl15a84YjHWP+q5C6YxOs3UDHfH1sIcalz1tfwHSRs3Zcv2Kd4j4yukFd6dhgNoQ/jfOTc66I2
IHBpRITG+3oPDZNLntHPkVFv9eO9OpqPjeu6jwLwc6QMFRZTJ2WamN7HDXCWAO3UoMnjUGYwnL8L
MOw4HnLBvH+3K6xXhF22y9jGGfCUFlSl8bDjlc53Z78yO53WgXD+s4m2fl1RbcREwBQqrBGq5+wP
h5E7O+gRX0nktafmoKUl0i6hq7FoOltEZ+On/rug4gzy/YWpQyuW9WYoWegSlcFrjB8UreT8qWqM
sdoEObSQTWhpPzozE5q938FnF58VfupLHL2k/rFuXfjCbnlCJbMs7rG1ncwjIZwb9gJ1ErBGKD4S
jABbP5dvDDSJAZeN/0xGXhU0jEQWOcFUzM/IwOBPY9RWZ/vPKtApgO9xEQfOeyZz/yBsuLK2g5mC
7qu02ol2cRPqs85ySiVHodu8x+gwXzGA0EB6s5ScxS7Z3VFXcWabcHBB1EKm/r3WOjGLs03L/1Ct
9EuVopFfBn3A5fF71FOULC3wovyTQ8Zo3bQsoxAwcgX/BPX7FvyvT4I5/QEd17/v/uStv62G8zO9
3VRCPpUVfCUdG4ak55+n6glyNCRMIFjePyXNeWafKN1fNMX5GzFD+izgUjYKMIMnZctW4955J5pH
14pRKmgWse8RaTeTP7fRdezU6bppae6xCS+UtrK4iCOqUXuZOj+cckilyrfLZbUezNQl+DF506QH
Hc9sXr0bg119oFYDwu6nSgB6jxxp8/tRAbx7c8aAnqNQ9BwlbAFmWlD248aqaeS7af56LDlAOUbi
KAk4Q3ktRFajZMNbmN65Fv/FYmhFbvlOmyNHgueNUZnbi2oMxxR/80uUHKySvan4nZUyio6fH09o
uUufvWzbR52ETsWQpGUkxlBI4jUdmxkmRq2wNpvHTRKHUbRlhX+OwQTdWovkr0Xk9eOk7rk5AV8w
dkENiuhextwzlaZnmpQoymJw28luZGB+UdMLe+tFdLT7c8EBwgNeGPVnWaXIMum46iAw877jFcnI
JtWmGEmdQbF9lXIKfsn6zrtTnPGD1dnEDm/7fDqrhTy8YmZZ9AUVbMmNp6Fgp0UrCIdCyV1COW+d
0Gf//3uJvvlZxUb3CvbTTYJLzSHT2U/uksMMTBqLhhkSu42YK+S5ZtV+p0IhSv16vRz17fKqNIcD
p7DfnKeBecOKJoKYPFJg3H/ng5EfuRKT9nl8h+amh4nDxkrZuRZefBwbXznu4CV/VftgxyV+QS+Y
HFrq4XhDISUC4lQlLVohzRtHAl0x6G+091L+GJdV5yx1+LefxEl79okF3x326nfHYlEiBKOqxt+R
BxEFF74sPodOfL2ZI02KyJAeYQAYWW0wbH+BUKZeheJVLSXYJSDGq8Czrmgf9/U/FnGPr/Q19dtx
0dLN5hMkL/5qI/n3Nakyk3KtcpyBreijbvVyz6EJqUuG6+bSZLbbuMQvsFo2va188HvrX8EwBRiF
E4zEFsQI6VjNEWOctlBH7sxtdCK9mO+xX3UuByqWN2mbdhYkpEtqjljKQ8UD3+uu+FZaX2IcktBj
TPgqMYanhMw8HMv0Wq3DRrhhCu3jIJrZcQqHU42siilgzrpq8MiuU1tKUl2xEB5xVmh1PqtTvpkS
bnLbplw2D8CtiLgxXtCs5szASBvurKq0KIaZMmIh2CeJz3ZRwXf/TZ3BOm1h0ZaCakANymJ8pxrc
a7Xl6Kyp+RKLkbY+nL6+lkCrPD62hBZmT/erK1zdyavDun9o/toU5hzB30y6xiRl/PkyJzelsUHk
4UzGqpRkJEAiUw84GtN7UN5c7rAvL3h4tqATYGIq/B4TK6lu0b7yx8gaRG1FYSHknBQfNNz8eT8T
dMjzRhu3zcgwLWAAHhsI+1+uflYoHJL2aewnidyNuKIVf2pojAUNdB+9j9Hnh6c8P3WAio8aO/j8
Fgvi5PlLbl3+Phsqb1r/BbJuvU0cHbUW/mFDypOc9m3xnSRmEqK+8tt+A6nkeIVEDUBVMVh13Xof
JsSxEor7fanLAqLTn1sK86Y/3k7df5X9Vz/zyWSWV2zAzp/LdXv+D7YnsItzVQbsOrVVtY4PGNay
SLaPdlZKT8vpewWinpueQstUSA0QOWTItvcYliXflhgNX7ddjTeYnzhZedO4aXAFhlzARSbuHFCI
Ui+YZBAt06NsN8mlpOcT/+VL6LajsH9LCdb0uwr7sr/BXl9nE6YcVK7GX3El5yGU12wsI9S3s2n+
ycicZeAhoD9se+CYkIk7QthWXZ6AnJnITwzSFFxNc8klu72BV8WQuC+UBBdYHFGLPbhC+ZwuhgnT
kF+mIIxNPd1NH+Q/PpfveVYNx5uziEuMAmoGLFremiFJAyRukVYLLyXwzs6n7tKXdZOnfsmx/zwD
KHgtsOS1c/QqUNJOD8Sr8aPfqCQnp/HiNAMT2xHXsYf/LlTDCby6Xnd0jX9eLozL2GDiW8WvzyJN
fVJNHG0UF0LZ/aaogLBgbsvFsKKzGLZtVfn41M2J/YBKI83rWqnThPcZK9sI5TVgnyfNwSUG3XVZ
6mWNFBpEZ7+pntpStYlrYi80RJHbL15KOav860NHvs9LIHxnC7eTvwJAKSMq2o+tWrNYCIHg6N32
645wbF1eFVSztB05nEr9u7TA80eDgrf0239pgFAWEDCvN2lW8/twKukUTHwHKONTdXscsnFgXFp7
X3tPzCPfl+VCAWKGDIyNoxN8FLdAN3bsqJkKzcN42UqUWIQFHbmbu9WBekSHA9Sh0pit//EJbOoN
VcOzjRa2ivt14zu4iV6qs8cwkQ8bz39dk/embeTgjI6v9MuF/b3nLJZmuOh/gW8wEpsdtXYm2tDQ
w6FUrygJeRHPLgXYtQz9nX8c9eJNSCh6LDu+R27Hg1RhJzFkwDs3P7On1LSOSYzCLAgh/o8DiafY
fE5hdhnUV0OmG4Q1klMgSN9ucKhzO2slq1wEOF/ZOl+5U0Dm1sjbL+22C3zryfrXQP9jG5wbPfO6
HGTkTeoQ9nJQQSsfb7qScjCD5bLkyPL0BG87rSGDjCTet2TTLbQ3tAXx8XDgbWFpjPJGTxjTh+ny
+CiDK/W2k2MKyo2vF4Qc4xgWHoNl/P9aRBkM/5goV9/BLyvL1Otxev//91cSC617zdyGqokEHerr
usBW32NoUn7ZCPpPeXn48UmMVJ09Rp6tsL6zJslUYQEdoXgr9sjKyB5OTx1bztnaZVq1iqkStOWl
pL3E1Bl/7AsvEa2dlzGELi9ymb8p47wRSoACUY7DGxtOQHzIyc8YuLZwkpeCh8Ohr408JhaZ+pM2
fxzOp2Z8CgOYu1y60PoYFSVTwiZhEvLspXKj+WcLev5pgm4cT3vg7lh56ek59yyebQ0K3bE+/sKR
5jGvAqpVfoqaNMGJpbFwPFSRQcfXqnoxyScqbPAYIZyttrI1j6liooVbGik80xIUq98rn2yER7U+
e7ZJp2io5g0nyfiYpLFupDyqfj39UiuXseACSyCzOEBn5H7IzudNgJmHYvcaeDT5UWG7oLbYnp43
wVBgvmH36VjKLXsR7E+28NTKI/spGBzDj1VB0A6OcEuQWAeOt5PjGDK8JNArIeVOblY1E7PTzYNn
u0dAqMcdlWr9ZiQAe84uSJPV5cfkQU7yFMBicNian/CYqx9W0l2aTXhMgdLzJ/lF0lDa7yd/UADL
5gKxN2kUKgum6lz6C600MWV+b3DnmBY7l2Er9iM9deM8c1m70AvTa2mT1AS0SSe5T0kglrR/O0NG
RcIf/CgR1CIBUWCqmN6BxJQDLXAvyzUz5/IFzMrpO2PQmrJ7n48jW8QZUgTqjzXID93tAhnCNmmQ
o4Rb1RoS0DeKb+dl5MYhGtv5APSBvegIMKax2pGs2dzgwNkCv4nloNFxPrbqzQEQPHFFxTRq1uzH
fck2vkSaV/QGP4s1QDg7pZqW6xIwOEnUuJOmnHQaahwXYkOeWY0ulXFE/5RJYzTnBR0iXRSy+kIM
2/EpCnQhnWtIFyqGyxVRjHL8XH3W+APqDChUYUkvdIlC7LWzV6l7bp6DhFEkdPcNo1jMLNwcIbFM
mQRhtHwGY0CxJiymawow2pxa3uIzs2di5mmYoNM3X6V7VYJlJnn3z1PV1owb66bvUBdHFSTEgDFq
MEGHlZt9IihU/MOsperITvJHuVW0hAk+WfqOpyd9KXPNiCDkQhKstHuuutiv5EIfDn7kWzKYWELV
GXERkP4TV0vFAGsytftoTLQKNOJXDeF7/XuyLGQBPWHu6+27gtu/ScposUIbQODH3gLituiJpiUC
88k8rjX4Qx4MYk+qsTcix0EG/fUd0m15ujisJfUTW8i3KBr7Pvzhtxombgcigmlb2xvgFtklDxzY
G0HL4YU7baCSFgVJXt/S01vzMKilXB2srT2i25wOp7dSf8Kk+nXqGyWALZiTloefLZlxYpfERz9D
mKtLpoIFO7KM3kYvstaYY/e9OSP6kJVX4VHZYvayEXjaar3CscxGyXLwfU8cN51GlSj2QghD/HFB
BDYu3GOM0INKlGjy0iPgymrxlcYYFY8DFaYfwxtwMETVNOXNIUf7jH/Qp6dNZlb8GlnV2wKyJPCN
fl3fpcUsP3rzwVHBU8I1LLrptWHB3uXDjva6Heb07VNKYE6i33qn9xicwuwbLPj8Fev5K1/080Ks
V+Ea50Bza+7y07gXPj2HHUI7dOhj1E6OIlUrH+p4yBkZdsx35VT6l1+Sj/6dj+Nza9tbL+vd7a51
KTp2NwKISrli09XPB/NKNcHsU1px6v2Rrtrkja63ZgREIh9ABOsEVJtwhCE/iTR0sG/qFeh3Ef24
HN5/tO6NpsbgQYD4+6c/Cd+YW7h4Uzy5kkq/K+A2ql54wleyK+GivDjEoJ+b6Sref1HGtRSRomql
3Ndk+sQsiwGSsoydWiBtL/DDd5xXUz5NFqYuf1SNA0lq6xKE//IqO+fnoSh5yov3zQQ9ohyjifC+
pMG5N+KCFMsmWJytKIM4uYO6bVx9/DNO9zhWs5eYEM87TtETRGJB2LHoVWHE0WDcsokiVb1DXq+2
MBicPuTJlsgstjGXn+E1mS+uTV77CMuGBa9Q6hBPBTHST8GgUIKMNtJK6ea2krDclt7BYX+8VbwG
7LYWvvUpj09EWT0qjvBKUFBdz1bc+lp7mCRkOEAQU+iJeDEdauNrY7lXwAd4Nb6a6cTizsIh2UyB
k5vvoVGNSHBVkANIXic/4Gn9UiMlj7rhTIIOwgiUVzhybHCRnpS09NipRCfTY0htD/Fje6dnxAU4
7OqGPhMGRKQbJWpcV/fye3Y83Sk0JajZS7lucCeISZJGvWE2iVxmtUY3FlU+pQUEPJWjF9L1TPME
YQCwDpv+g/E3XIUOHQhImbSr62sqMT/2edRoGo1YSUtdS4uh3AzLd4XfLOy59y78ltRyxRenrUFP
J4WoyFleV1Pk4v2CiEfCLUqrEh3LweqISaDThcxDjLdcHSsx4eMwKla8AvJVrwKJHsM35DPv0Wdb
MmHfWN0DrtcxZjUailvn1DFCRrMBdkHmVzmGdRi/7vxxtEpzKOYT3hOHH9IiDnfIXWAI2jfWbwBI
LyVbvcnbXtdKOrJNSJDN61PfBjx/FnwklWmyqmL2fBklwQohXhgB0vaMGHEfvjrdlnkXCNR8PBdd
dT2FX84i/ODn3IV7/MyPw47N/vxGE4z38LLO2wp0T98C/Oyl43MgIxLJ0KfveRd/Npjh3P3oewHO
W+hdOL58RoESi8Zg+ApCYK512OqYTl7KpNslmlqj4YoL1XbFuKDeERYjjVQ9l9+w/F3kouGigHic
KncaRI580t3db+h49rb3CkvAGZsmNEy/yblxSvRBmL2UKi82Au87KnNfdRQiQMgv3wE0BklRESMX
SWYl5/MknOM3SrjIpAdL7RfqQHnBf7s0tfOqoXjCL0u1+wVt9vFOOFsvMMmmAUQv9C/2OrXck+wp
KBzxDLS+mSriacCuR7IKcvvY0f3GOWutwaWUjElszgm+p7BRyX8d5LCGhuORXlY+j3JXlQ+ygZCo
USXi4gtksd0BWM8rxT7YD5Po+sdyC9UqIXgQh0SmoYv2XxsBDtzOiTSUEygerTjCj+HEQ0WYgDFm
KexvV2ufLnjaemyusiBFzolbezodcXues3bs8Ldq4M4ckWIQYuVPgZlns//zYxRY6z9ip8hPFYya
5szRt0llhKiD9JjWYZtVhBTjFmpSfpww+KwySYNTFXUn2X7PKH2z/Riz+1feOn40km4G4CRgA1/S
hdWdOmyQz6uMGhNeOpnjLAiwMprVITZhup4yhSDkT1kKGClacbQ6GYAsFgjovojjpMf+GOTMTphs
26uhmYmHu5yVZCAPgk0vMBVfoqUdYpyiC2UhTJr+0MDsolVCuYSNC3T5+KVnd7YlvGLnPjrcgxZW
FKrs3pC8uGwjxiyPLNjpFQoPOLkYfUF5T8vkIrSI/MBLx60cPh9e8cu89iUzqBEhtxb6Llh8My5y
t6QaC/TEw98DXPnBlQhrTigway1utl8dmomB0Lxl2Cxi4b2ItfATym5NSs1MYnYLW4AHDALt0/1E
1RATqBdJcrL80TxHEBGo7uHMQh7L+W/3nK9u2pS3pTBvc79opUEGWx+F7OZoWhqmX9RdblIDu1i1
0AFApuuF3Dxe4ERJQaoqXK0RPUO9AWMLQekc3piiCMHrzO3OLQQye2ZAzB+NeNAhMOj1NMdwIOhF
+SU0+mWq6gUX4FmKtirUY31jjDzi9Udj4921T1qvrg3q2diockJ/cPFB2gwcUSB//xOJGYgWYfax
Spas/wA0oFHzEBXvxHqe/W5747+rfJusdHGYI5CUMf5AGed1Ro5yGrS1vs8JeXXHIHbpgE6kKxlU
54i51RifYkArvyXhFDsme2rem8dOz61g2E7kKiBmwx/0a5LQomfpKHK9NolJi1jpEkWL3R3IHwRU
f143NV5KlDXXGcZ4lDlwrk4HUkGmaKgj4VeuShqAy1rgQPTapsKvLQhQGPh6iPfA8K3Hb/KSvjJV
1+FefuCqkM6gjoyd+ASikSR3zmJfueuMy7Mxd0KGMHOOw2ZuxF36q4AH18LGzZZ3kxNRBct6o1gH
1lWf4aopVup6eUf9uaqzrbw9f1c2o8buUIv88HguXghjAMRBxFnNicXQ87vQS7579IRRZ1NJhn2q
BvwOS7PCERnYKuhVDpf9gHU4FaKuhO+fvFqSPLR1c/4033c1XKmrP0Ykyxm5RveXXhTZqWxJniVw
MAqnEU/9s4XRc8JNyt4XIByerfVUXgPAh1K6YPqUfESDguGsMMis0K/asYLXoI5yT9ZtWm5nSZeY
XcmWzWM1pE7Actli+XUVY0LTHyJ49/e1VMfjfXvAEHNPb6bgPeQzTKC4gWvh8SCxvYDZZZRQCU7W
OrVY5llcsINxbck0bg6wcWHLW0zq2owT/iafxHFMOPF+orQxML79Ob9h9/Muu600ZhZkz8wuGOPc
dG/cQVRK87gEJ0lToxeJTWf037O5Xs/qOxJMMKXj0wdh+Xxde2OwKdn+256kj8srX+DIie/ZMnnC
9ENxnAt7u62b7ObGlZSROPt9G6zRKb+PPh3c7C9u1TMa/2/vk2zPDV506fz5HrL0RsbDKFxK+aY5
oOuyf+4VhPrrAxpA9D5N87Hd6NRoYiplSb2Qy0+nQramFoZNzAaX2XvP11ZFQqIZZ0ZF0k4ikaBq
yasoefcNJuZEo3hTixSGyoLgJs3K825HuGOA64TNyFp8d1Ff0P7uHHl4GkvqrWbiUOW+8EyjZL95
5QqZ3e0IDXXbzykh8yhi5NDlbDrE4Egg9jPjAAt5FG0w8vqJmwIowRjVAoSflNe97A5F+HVXAhCI
2ix4OoPE+lPravTFIyDNR+oa66S1bTYMD3pmm4Nw02uql7LqkKbAIWmIWIgc3Pk8YzkcXgk3Sg7O
vYEFbHfZ5/36LodX2q474FP1QQoRxdT8UOo4Ew4BqSCoh2xkzLLQQ+QeoIRW8jXAxK6DNJ7JeWQA
RSa2TGmCv49C60wvkpQM6oIPRi8OT7ChGvH0QRoL31cLGGSwIf5gnDE2HRmwJ4V9zq0kBSLnqxuE
hRtUw2R418OPRTqe5C+i/l6U0xO4xTTnms6D+KzIXjAp5eckC1l1PLYV/kFPKcWNr21A9nczuYoU
Y4ReguXKRKm5ExprnsWfyNTF0rGe/52tvPid5bAyzLNggeqD/uXuPjApk59Pjhegp3Xw/iFxSmaf
UhUE0y0JzO1OO817wfbn0EBBIJSrsGsG8o6AagCTBpXHfnccmb1fuGaYxqtRHfxUdVlVqCaITHWv
k35roxWousU/57D7jX6KwKR3Vv7BmwRmrMcqc8r57yMssBBoWv8eVCg7FuaL0Vto6zHkTNszoShn
6k7/FTMJzxqsjrj6E34WrlF3nOnm6UJKgTKtQ7VgkocW2GNog1L5fYsSNJcEnwX6hSKjq6fzqMsg
X9B57dgI89dQTNJxN1s1fChqXJFcq5WePoYBN/vGOTscYXOHpOyQ0twMf16Vs218AdGQwoRtnYvu
rtLenbMY7vkW4mBmGN5mbshkUoMdSAaguuWIa5SRfiFr4uiXArC8s8XAv/peI8oLaTYuI/6cGV53
hPRBmbDQnTG1QgIcF2P+u8PdR4P+ywBGDFawSeERL1bGKOfhjxQZpNiwMW7pI4IFPH3oyvxJomAq
O86U1C4OpSIvJ8RLq74m8s1U0QY35qChgN0nPpq18Q8KMGS9vV+3u0bWI83w7pOU9M47P5QShc0T
cVzYHW/R3ZfCfkQt6eE2wbSgUWfYkdZyAKYM/97fDQpyaR0PlWeTB3h/ZxZHF3kHINU8nZc1m/lV
eMTH3i6osVM2BUaekuxRykdkv9ofQ7MhlG5ccLGy0boBBF0G19Mssmhje2gQzjyrYY4GRnLyXOYl
cgc7FVSVZc5Rb6NFeQ02/kHAgiG1HWZcARklwfz4fa/f0PB45qzTlxKVVrbdXXXICCf6UKR0+hT0
Bmq5XFiIKazqe3vLCCvh5cRQ8XELcxDjmzr8R3ChJLbarTHew8IR9buLShIpz8IIqiYkRFIOSl24
X2uQ+1l5X2rznvBoOgX3l3H/dVUVTJlnPsqbV0+3m3KQpCUujiNN0kJdD+795tkCuIHONGNPoqI1
gdihK410jB4fSyxX85D/UhDMgRB+nGAexFdh2zx53grU+bYTFCnRxobG5Sra6+qydSWn/7r/pYpx
068HJB0Omc13uKXjcHsE4X0CPO0+nQSul2wkj0HNLf3jsMb9w7P7wPkfEh0pZP8elI4ObI3t3Xf8
pbTGp63TwQZV23fQ+QM754fq8SlmFLjwxFEcV6LlxIOOlDkr7+1LDKKZ4ZnVelzbXezCR2NUNcDO
YurXYuc/Lc8reHLQVNVWc+HJzXNuXv1ElqD+P53drZZLxE2iiwc8et1pKqrrnnZ04IPTPTXvina+
bc6ghQY9J6Td/49WUfNLnpPCVODXzbU0McJIHLYbj8PnzkjjOe3k0qIk1M6K/wXXTbnKqKRSh+5H
O+8Y7IEIxut0f6BS67Lxq/x1ZCLisK0suT0/0acavuuo0Jlod/04iID9Ojj+zclso7RbMgqYFpka
uVkwwq3hZfVfukYRg70Kp34m3Qjg3jXgCxSaYc+cuAzNFBLOXS9hU6rgyAxwj0CPpyC7wpLqYkhm
d5IVsUZKXpe6F687DQg7ZOlDpbmijLtdqGLIdM6ASQf+9/Af/sAzxcJqXUkLSYVs1fXUkBex83tM
I6EJ5WAvLMf3x0b1djdxE0KfPyqtXD7l49W8tW7tFDXnA1ofj7a/HMFfdmkUgiKGwv2EJCVwXwlD
+ET1WG3gvP5jIQLSSv4h2YoJ4zyAldNPwcyzKxhQGi62ykZ56VSbvA3q7M4yvqtF5pnV7rRhgLg/
a7T/u4RLBpFVU4/Hiw8PoP8f5sgVOoilJZrX3r0h68EBMOPqh/HgIE7dWhNkxBaeNHOFFn0XdYZ5
PElfgjbBBU7osoLyo3ZCpP0FO6XYgWciN9xyUOSGoqm6HDg7PGTYE5lxIaIwWCiXZZzUtPTeRlVd
wzZCHyOwvNIsjxkwnMxELL4ocNF5f6Hd0Kt8pUshKz7oGt5/R2CnPuzoYDQdRMZL7RTWA8AgPF7I
Zgz7nh7tyTU/o4WbokBEMmcEfrW0HLeQ/3VWcINsfPg5rQqRIOoqvdBgLj/OkN+83JcaoNUJd3fk
5oqkHd0zZbeHXto8kYWnFTPS8RcpWsCwTyYGYzqkY7wADjPCQqbRDNthzx0pP/lfgG0nw8nVreKz
13+H8Sgwu0Rv4ao0TwFCWFJMRSIBikiavBMFw7zlwR8oyz3Jttbpy9++hquev4WNdR+Z/T768WC5
9NyjrN15ekltX6wv4vYJoz2EQ8qaClBBCPS/Gzdzz3D4jkdv8BXOmM4a+sFpwjECTtTcAZDGH1sP
EPzlur7NMYHJsjBkAd3GteCV40Q8cSRhU6cdTiV5IobGzAzf/m0Kge3mNIUiXOhbdIp5PB46x/vt
8Tl8zQ4e0rQSpikcX49t4u6M9m5yBRmlg1sca3tfzCgFLh470uJdgKqcFvmRHay4TAVp4lsvz1rq
HZDe9G6ViuZSPoh94EFa5+C8m8jsk9QeaaznjMqOu4oDxynTjWJJ84qMnKrjbT/y466ludicABCF
3i4RpFdCUo1itx3KLVmryse3cWqfiCMgDiHpB9s3q2ygY2+J2RPkZtwyJ++OLYV8sW0+SNI2yiNu
cGz9qoQzRZHPjeGO4QmSPTvupRQDtnSG4Spusxk4G8Cg5JveDgHsoxwQfsC7SJjpjE4oyUtuQcQf
TqqHJSwKpa7fWSYCLvZuFLT2O2tRqUgGFFe828LPfOVbeadR+XBeTvtAvOXrtekH1dfbVvjKny8M
Zh2SAxGaJX3gYCREd89G2WvhJqo5PZMbd8ws+g/W+wFAFAzPy++A9PcxtT6Xuj2aR3RS4SoNpnhH
Mul7kexBLjgW8FmzV9IDw33jJhjEGOYY07yEnZT8IS4pL+a7mILdphZA0rTEwPeakPS102ouGF2h
QGWEX1hP/v2vaLBuHF5cy7ARUywXY2uiIFM2Lpu/i3y7c0Q+LWjVE14rU6CXu7LmJUizwszaA4sT
oB7+6IxIdmt56kjrgVqDScqp9fpeJAOeBESvA8nuJYS4zD2ylvcXKZX7IixjpCIO7RMbH9HK4hZb
QhnOBWv8EmqQMidTsdRdMV6JPux5OqEIAZqv+tGWZnm97R+6G8neLtFCX98z+zqZoKMoErLAJmCX
t2UOhACRhq8ww7TBg+bbfzzU1QaSp9LVfORpFtsJBTDNjoNOAvOHj6j455AIkVN3KBNcfXVrWORe
eOQe/lioGkwJmF5BITnIfybNihYlFqyrP7oSz6pMIUpFm2vFlhEvT0rf4REBbz556sgh3hHAP2+5
yy1SzeUFcitC3Oh8RmOQqsGyZlmdiPuVWKgXBoug+jAFghWTncfv28wYhmJP4LsTRxCzU2DeiJ3T
36pVpC8ItHvHWF82fq9z+aFNpUOtAleWLD772BuqvU/hJd19EbGGmUbCjr4Dk7Cpl8zLxQA7g9GS
mBmnqUvBPzod/uSI+8zngBPSG4YbTF9vAMfKvfI+XpB6U9qAAC/WkRwGK54gBE6es3g7gI7r/Nr3
zE+d0Ibxh16pI2jCEDs9z4mpjPZx7i0FouzFsrjbobuQczJIOSNpo5MkKBO1lyusem1L6BnZg3hE
V1sEYjjofkB8lCFXNJh4chZnXuYJloHedDIXFAb1KejTeu8dYcr1R+vq39yetegLetinmfTP6J8j
YfUE/XBUJfai/fq3oborBf70scnnZWGI6lsb1FMsHSvacJXvMiOlbK0OkPKi2Sz1dlj4rkGKDRNu
CbHIVrIymTGOf3o7gsA1FOVBLj1BBpbIQkxm1B/OQARIbk2GvDdewLbL0At01k1r/ggq3toUPuWZ
5QD/2W8UAqOdXsef09nS7e84LPrYqOJox019gh3WSwh/RM0y7BNdzhCkLZ01rLeLViSkWCajSUH6
Uyd3RPeSamMqQPESm/c0FH9i9g76H8R0egrVf8L1EjeEwuXPxvIETL6MKImo7rIRsgwR5XqijpFX
kVx9y9mH8y67IF9IeQJ8SR2OiatkcPMYlyNUEZflJcW3fQRmB6WTtQpims8IgV2qmYU84+Xh0wSn
kQ6TfLruCPIPIfAOnomB8TT1PsTiG2/Nycjsky5mB2+8oKqEyNgAgsgBfJTRYCscqIdvO/VOimHU
gf/KDn/V1O+RDO98iVBNFqr1cUq+fhYgW4063XOgcqhDZAH2eZGMGReUCs53JYIzB0kUL5m0MGWD
XXd0t/DEAvsBk3WOIDkEMeC4nYQZuRYKVSasm/xxG+RzRV6EAQ4dY2hhIPv50iV0BHnQVC/bkj8i
wtUDGcVfZvJ/zKMO0inAaizjdBLxXsh7ZnQSiJOPL1usVz+2DmdlxoKZ3dVBV0NdSZmonUO+l1xa
nYdKdc6WAfnjAfwHeDaZ/7oLIvALzJvBH6ynZSUkTPZbNOZM0IhfQFhWwHXEpnQlVDkX+TUcg9Eu
RxZ5oIvwcJXnBQjBmhckGFzkV0bBWD8AhCiIj8k81nFJ7O1Whv7bHGgBhqLZHB0eO1mUdCgCtqDs
VfjJFPEgxE1ow7OpeyX8gJ8MWqW6K/phGcqzbdiB+D+GQBKAQVsgLUl1Y6uN/8V3gBi8OhT3o8yB
x8ykur3AItwxxJKug/7sK66n7xyOLuHIGi2UERiMfVSrqeGnS0Wceqw5RlZbcJdp94PXoIBxXC0V
GQo3nP1JexHzGwD1+SHLXjab5kiW1GeVpbZ+iAYa1Z1zZ4xOY62IjWV47LdVCELBwEO4mYObdMHv
00nEGYQo5b1FCuiRwK8xWuZV748ZAGw/q5Xmi1QLfRzuR0RK4poUEJiFahEbhaoDEj9j4f6NESGE
FfMVEksNjHP9zA8hC5r0HAAlAcvtWwLYwGIjAVBC2xI4RNP11+QvfXNKADxJGBzMeM7BeGVRP0mP
W7cOHBoJ8mFWUmm0RPUKY3HkJP8r5B/Ndz2DqxUazY6nZHjm3rKpt79EAFprsBc7I0UkD5u8h6Ck
aJ1qxCwHS4qFrhre07Ay+AutivTKcQiu33qRKjkl5rbIoxhxsxm0LagO3EgJKqWznpxC+Kuiwe0V
v0L86x7bbNh1mRwNNG17Vz7sxeEsu/6q/lEyHQUgmiUCKVkPzUIZ9jG0lerVuV3RUP1K7yCG059u
zh3SdTg3dkaQEEDs9+uJJ/H6vHZ4viGuUJj7Ql8O0bnDlDp/VsZT+sfQYIMcw/XwXPZfTSREAbyG
Vx8ySfHaqSYRrtue2jKONzH1CIXVvCQkuluVMgWjmV8fgnRGg6xVyEn4npX7ZWRpRgAE0/hIESd7
ztFWsRfLDYbJg9hOFyUJolruDx3D7p7wLetdsKthcHavZqlVMV/TQaIN2NJJ8PAr8dq0RgEKxwbl
DzRjm41Ulhp1gvFbnGr8XjdVihlTsOi1Ykig3pvCtT7ATz0WmJFKNlG0N1lBXyIh2qtOh2Gl2A23
FEiJ6jfTOEylBhmN9fYugWCh4B7NJfuh52bcL0DpKjtuEU3rdbL9qsZm9IbHPfQ19oyQdOYJP1GB
E1q4ZdO7G83LWiIW3rp8rfaBkYCt7wBqIeiqf2fOZ8Mec+WqGJc83F3sgXULKnypDCd26MMUxUcI
Em21hsp9pa00UFGgsVoHSJzwji0SCSn0UhVOuYEQytJ117QDxmr9c5/PKPQQLeaqcneIl6g9LIOL
5zXKk5JCdMi6AGqO5bEXEwRdYXobPoQ19QXpOU9CJ2gLS+VWBu3ngyQ42R/v0lHrAQdsMCVDF7vL
3HNLO0cC/xHCJGOb9MMlnOhCZGhzbQAw+fgE5yiHFItyhA+Z4egBhIOgBaHXTg9t0Dy3co4UcpmZ
/gIQVf7LH/GvNCdOtEgqHGtwGeBhbWzzyjGQ60V+TUnrPBZVTrgRwUEIVwfohiSXqhwVDxYXnGnE
E+mpnXrj4dBZoj+BcxMpbuIOjTM4X7rPhpPZA1QOG2iNaNPQ5cjsQCnR693Ih02w3DyIIPP57wNv
N254+Nx1LdMx65ECGAtYO/5fRKRqWyuIOmvpVsYJTMdcpRogLce38j6Nd6NTdVLvWU4zqzvYA7m7
5dl1L232YkwbJwAUNq+J1L8FxhmDBXkCsH49gpMXFHQc5qObw4jeN1coaoE22+pAk1yGgBF24DkO
BW8mPSlqzOarm7pA/q/T0ph8IB5RL2CSKEEjJxmWnFNw05WWWZel2M6MOqK9Scx907r2iIWUUQ60
nSAvfvSBvoqhIDxblyZRHxn/2e+hd4BcGJmLeiP7Sm2sbwGR9yVahaxMonpiUebl6IlupwWggTpu
V1coJ+HaWmjxIdlKyG+p9NbE++QmLiWTmFHVQpFj1wwmSa6rmHZC0CThVW+38GNSWyQMZV9YofQE
0orzaKexibye2Xaj9CaPWVzktcxluJFWjy6pm0K5ya1Xf1KtPPFTHYVVuyQ5l4HzS97qmQiuhH9g
TIz6rZ3Bfc7LMeq4GfPgLTdpQp1JU0HM/rPvl7IyFBfXMcFH/eP7bvLw2Wwz9LFIqE5pMhjRhaFN
Fc8epEK72TW0PxzKyo5dXDN3NM0xdnnXSYvet4U+3WXbD3Gyr39A1zrTyMqbCy+9LFmCZ9ynopU3
9abEQJgDXrSPlD3jklajN0QcHp88UkyyPjrVMkmFL8R/xvk/oSdLW54JbXuRQHOnDqIy7XdbfA3S
RbNGvWtWj+3Za2gzJSlkWaK/tbKmcIrgV90fEE5CVTCdY7QWqzi/5zEZLbaANqxNWi0wS0c1Eo7v
atJXtBY7n4SJCYLVvE9yvFdxiycZ5EMXTLnySsr8IHtqN0mcwGNRNhLgqedwnz6R+1T19ttboi3O
CVeG2F8eeXu5CbddRTSpuHH0h6t3qfRq0B7h5qt2XqHkuuGvGwFn+tCTJAlvzMvtaY8PZUWGRP9A
lq6Jf0zV94/2/rADo8mv+OEgCgQTPHXp5a+596Z+bB2te+gRaEcsuNQ0iOmdq3jtxa72VdZuhA4y
Ar6gQMq9adJ0N5lCtABzDxyDTG4v7SCJ3lpNxA00PTOIqeJHp5FEilhjNi6Wa3RiXOC/umjewTyz
jL7CR2UVGUZgCo5liqG0FSzKY37Q4Q0J+W69NO9Huqqx3Aiewgfqpia4teKFNVOAHISbW7pFK1wH
eCELD/RX/PHLrm3CkfZ50wtibx3LDqc6KVCYrYkASDCajFR9UPs4IeD0Ce9NneSVd2etK7QsKdtB
YqSfbvpa0vHlfEv9V0U3myGgq40Xsy6+hGUB6cBM5BiBXr7WGicfvTf+drZqagMJS2GRiqPEigyy
zlxLbasJ7vs1uXffWSve3Qu3t7+cm5N6I2FmbLOri/+lqyTRRhuBREloy7atrTb8uL+f7uEgpa59
zHmU3AUbulpfT5/MSqaO9Xp1y6HzJPfrTA5VwyRrl/Skqq8JlIQAq4TpCG3KB3Cz+AsFRvi9rAcu
nr4CE+5Vbvtqy86eGd4Iqdey655CiGCWFL4WJNElvoummhNpEa78LM6g4HpgItYVQ/12vfgxH0ZS
7CwBzUqTIYa7oCsE28215pwzjRH+DbDRRcwRlaDHx86EmHla1gEiXPMktJSiUa/w82n0alKzxiNx
mnrmlNCy0LiWE7dfe/BgKY4V06n7CDvf13Zis/qhqGi4XUDl7fxw1JfwYewyIRuYwf56ztKzxQB6
/7udJc5nugfzOIvKRgIeqbi0biAM9U3Q5iyJC2jlTJzu2rMKwbdaKpZscOEc4p1XaHiQ8lWKEXbv
ZtMl6gYsAe1O7tf5Ed44KzSOCN/KWVY6ng+ye6MokqIMzB1nWLu1oqRri+IE6XJkDiI6XiRXcMtW
pFYlbbCu3VIjL/EWKeIMf1xlMUZmWPvmUCJAoMrJksKXj8sYpynKNE7WmKoKnWiLhU16Ypges5y2
EHIwFbg1r52FeGVFbofy6P9DwPEY/aqdBtOEXfvVEY2eb/Mkzv+uQLqIXNUeZc0o4pkGKUc68Xge
2ghzgd2pOlQ5sTxz1cehbk0nqud07HlJRTHyA7T+EEOr9+MZxHF+/Afs9Pmxo8FC1Lik9wfvYTa6
33vVrGxNSQGr7ABjrNFk7MB439p9sE72j5XMIQA9qqCJoRfJcAxUwQneQSB8iRzaer5h84N5GkGf
EXMDOjLFV05A7b3rwGlJJEX4C8e9bvCxqvxcNw1bkLDePxOcpZa8i5LTtb6qmIa+OjQ1vftCKis3
07Ptt75D9D0XrHxNmPZ2/RhHCaEugIxVTjFWFQ6S+J2P1L0r6CMFiER6vsWSqHwFDizFYfaastLq
jN69luLXRjV82adUrWQV7mJUgf6XfRnGgQvFmN2gOTY6HQQ1iT/bU9/KFot7mK03qm2/Hc/76bxo
YQhMB0vr7kzN9g5jLwRPd/bIOdJ/lNdQehvyfDkBj0o7KV/y/8d38VCUKBDgH0HSoQKuWJckcWlm
Flsr0qvQB+FiHtyLTClxSbc7AwQ17OAdEvxezWY+thTk37AgoSn9Eg9hXr+tKa8TgimW5y6BVMuU
j/86Pcru+wkz9oXNoddw0wjRpLgwoyMo8SHTv8dCp4RAZSX9C63N9qQzmQb7dfus4MxHLZQwDQNW
TVsoB5nmz8WKTsCcaWXjpct+aZj5PKNq70fgvR9TcJ5uXi15KYWKaf1y07yQ1g8eBlA7Yv6rEW7u
pp6qbVHoCCbO4byCoaZGC1C52904c67eE2T1+tluBveoQX+jw2VZN0G9ZYXZXvi6Bp8bSsJOFkP8
InsbPaE3W5RcByHPDXMXqmhow2maIqoNJQTM9kHwRKWJ5KhgH9gEwU0MOSNzWdfP46ZUVHQrTNMc
XuWz8V4wE4IlLwmNTcV1qgQuQKVkMDY+/jAsKufXJTV5LL/FYghRohY6wYNcFO/ZP/Ufp6xRjC/m
rfMDg4YUCQMSjbVul4NgTJlg+8jaI5c42sb7wpEk3kl6Ha2omTU8p3ba9NnDemuhprE8+nDkBkyx
kPimd0oizOAxOLzprCYgJwWtfIs9Iizya8zPeHbDwD1pE3WjlagvPcelW/rPJ37Y3Xf0aQlePV/c
y7DrAAG9P5fhKEMfW3DZvGw8f+ipTB+dDrztcqOITbqHX+pY+rYSZH9NL3EfkzgGYDra7NmmbrZ7
mKwU1PCpj1t6uiPkIX8W2jWZ0oWaYwiMP4NhXl7s7bRMjDp15On2+iEN0UZvDNM2YUl/O9s7CBoJ
JGIGt+wVndCQ6A94Be7OlxwSMHWivrZ0/JoKGoBF0l42qKlzDbv6pBTtdfIcv8vmcYDU9EGmWp4C
mbChZlZVEZI4/E+rlB8ZkMFMtr9JDQPn1K8VrpSvrtVRAU8qqjdH6N+e1mgtaG3SRF4r5XZrYlwF
rFqzDgqerWxmZll8byH4ORCN5Oat7/ghQLKL9LoLrcRKjRGkSu68se/lxMhRoE6K6jZzrTFbME6X
RJ/N88fBhZn/++8eMQgzg0HxBzXMTVwe1seNLBttZI8BrEp1ZZhd0ctptVRUqWUCZOto281Finjn
oUMVVS4tZh+fGSOh8CvAVz+xIz8LivDNTBROYlSE+due4WOI5VpVq3om+YgwL3TVu3dJA0yfyMhH
Hp5WKTwAGb664WyZlCI5xZSAxCTQnMvQvho6T9xgdpaO/WQ0eQParpwVRiaQnwhKusMtChMUbjKN
9nzj5OtofwR8hCrV2J04FFUAxH+DVZhmVa9flQ2PImc7gKZsqYBVWgD2zODsZiuD4KAPGeUYqPO5
gIlvAu38JisSowTvJx5ucY1qXSBuniRaTJi1lpi0rVKhETKUhg3SjCY6n21Cz1TiDhzhR1AjgUgE
B/p6B/wGBhyzVvjxF3Y9wUbB+BNvaY5Oyic6SWxxA3zWSaBRZOb4IiokVyjAYZp/KEgQr1bJVQ4r
1mzbk+O6GUUuzdY8FbjZBrE+hviSf70wyVZrMofqjXfjjHys50uvzNoXoAF8WCbxc70te02V8tZS
Q+y8VbLe/5+H5BXz4soZBiCsKljvW3NIxNGM9MsKIA3mfbsv3FS8Y7BtPgwJT6sboRqovamFb6CD
qNHRWpnxVFyYCwT57fTailhwOR2ARMk6VaiQ2y5i2h0vkFk9YWrv8fLbyRU5KCqIdQUm50cxZluY
pcDJw8mFrxnHCy89Sm0AF7VKfxyizCtfrRMq+0QewxGM2sKoGgHVYMeyCMwQq3aua6QesI0gnGPw
rerSvypyod2erzWK6Us+vuLAAY4LHxKs35kDFnMs8woYUWYg5MuWLIIDAnK4EBYt3SQXugaecX9+
qidaBUHBQ3o3O+FniauJ6mtBWYrpbe+kgmFs/MMgD9bLAEvzQQTpENDAQzW3vNezdAY/DlMVud/w
rvPKs6xJB3VG5hsyX/neregsjrjXJ8hk7lMckS+5Vtsg0gUZjhfQc/bLNSXd/s4QJ+PQ76szsliv
lo+cJxj8hL9BTB09REAhtwlOq9L6PflCmliB0TCucWbWdL+XX/GEOf84nzSUmFlnrCY7CAE0Vkbm
9Umy9h+xmxb3+taLKAjDtQ8GzV7Jj/9N6hXgE4dRV2xH6ziCamy0PhjeK1sAu0rvcnkskjFnMAmj
Z1blb251gtQhGqzb+rqpYebHhr5xf4+D++zNorLViR2EI5vkbDFBjRqEdWkpVlDZR/CgF6meD94B
OkORkX1q/L8MtayxkjEjHIMzfwS4TVKW5Xm09Nu0Ii7bc6RkA6uMlv9DLczcQXuhOJR4gWvwvpdM
hNU+5SDHpEoUnMQLweXnalwvjQnvLgiB+FzPAHuJpH8535fGxo2ium7HS5ZZCw7ygMcZIj53qgs6
ckrfDK62L3N1qxHv5/jyhRRFyQdcNn7UrQmN1I35P+ebOAaAvhbbgm7ZqgHBhODuy1YCdWIetXF8
AuU/uzDsYe9uVBIyEe+gPG4OxwZp6UmSKGQGSe2SYyKbvl2wNNUBCJHPTZlx5xS4atiq5iNeCDtU
FDBpO29QgqBJqXNTdymnHLXJNfQE51vP5wl02fEoT/jH9fPosdiybEheal5OKY6b53JKd3pIo3xH
MkXHnMVaaJZT7MoTwmx0xxTwGy0c1oUEf+4D75TwJT42YFuvZchFQTWrE2+a/TORXRVINeBqAl06
hIgsGeYac1kQ1S7mZBIWEttbDkYwEHSlcUO2sAmCnvsETvcJpBLK/cQz2W8GGluoJ8oIu1nJZ4D9
vS13A0NT0+bx+3Cf6OYW6VGEbvYQ3lzOupN0rk55qmG65aFp/ejk4W+4uU3XBtiJPdSwiLGPAChh
NtPZleMrMIsTQAtAROLcRnO4YT0V4rZO/IJRXFDYddTPctTErUY75+C5npCCpdHAAaKgPxJtEibd
tM4biy4BpR7kMALdXTRvyjIsgKAC01VD3/ZixUBrOh8JYWM6oGLI0WUkLlpv8sl7ruZZicOH6Wvg
Qc/cjiTZ2G8UFMR5gtD/OA8F00mlymKXMCvpWBrB0O+9GfS90yg4PhBwRa04WgQIc6RQNq1vhR0R
ZLa/4HF+ot+2w3Et2KGoUr3i+fWbMo9DiInPxErbuepj5KSlYWg8mH2tpl0uaBFwlU/6Odfrn+T7
70ft1jldD/YtVgJWLQTVSROwLvg0quVsE6/mPn9dNshLWjqcwhFi59b74pcApEpJUrLdbukRGhl/
aZCDDs+f7sn3PnrHINlLnLrciBzwcnZdcSM5OxygI+dg7GlicuWCTAhKKAN3JC3+VEwpUb9MggSf
jpp5fdlmvwpA4dzVd9zpUjd6u4nWPFkO2S8dOXboc/J0iJh6rbzYNJlnePD8mHJCfGafX+OrgtE4
4HVL75j+GESErTrcFIz6rfjiNUs/DMKwXrY9atThGgnxj1ki7QQXg2oOaIFxsNSkfmZBf2h7y/Ap
yi5u64AmN6cHDsftXa7SnHfboWoBqPn79QIU/rFLvRJcXhJXItAPJMH7KnWSQs0X2j0LsiySvmhi
RHJAgsp4peCMQukkSkPD9rGnJNcBw+PZ3RM1TjWgMacZCfOGWDiT9rS3LWuaqvzRzhaAxlDL98fG
huD7pCF//vjXO6jbXQUv71rD6/QuY7TAZ4XPgRffZckJyOrVZaV0DSGh7C+G3Vi+9qpq3Vsmyq/N
HzBBcB0Ni+4FNFjbb2nxZa7y+SKzOvafWwCKeuc32m9VLBYcp0SyPU7/u1fW16X+osNYu4k2Kq3k
ui/5lVeZg0HnyrgIhOvihEBpAceH7r6c0vr9JL0h67Pwq1zf/bQSlY+u22838m+ASa8yI+7ql1Dv
HtG96oadCabq3VixHE9VwwEW69GRAbrMea/ceHEvnHTzApAgLlAKgsbzn62BMezF9bmBLpjPq8bq
0KKoV5s0A5KhPVfIlTg252ADNq3pAo76Xf70wNrx/1amKS/VNTE7fTZkoNLO9lgl83Sayxsps5CS
TUzjI5AQcA8wpisJ/S/RHAr+Kxstqphn4/h0zQ9ddtvoVTwWeyzpCR2Wsc9dqYFCr0u76oiAjwhm
9UZX2RZYem+1N948fAc2dU7PeoPJd2sWaDXCefKHhiYduQ+Je2QwXt4Qrp6Tsr7Ri0a3GMpS5hUn
9FtOvzx1YOz4zpGbqOviyItcNsuPoJu2FZBrmhFvS5YR7XCcN1siUWtr5zXux+olnYJqIwMqxwnT
L54EGogqSLM8PMewPsdpyqxEdv3iygYJ76w7uI88pcA/S67Y7NgFRLuaVmqrrrwhDwqpZ3mM69AV
raQYoLHk/ZbMuzE12ePsRyq7fqKXrSiJz9PYI4G2vbyD5158o0/eCuFhkirbnWm3XG/DlRRPnq40
QtokkBTGhXBG25N0vX5tRg6UhihZNThlzBrp8e7x9kZPiHuqF4rZW25siaEYceL52g5iYhVbKm2S
kswTLkHBksy0W4uLCKQS1boaUn4OgrH/pqf02vQ2LLI/AxxoyIzvwbiUe4HxYizMlPoCKmYVPrC/
Qunnf2Tv9UYsabOCMTrz7Nq7fJZ/qrnN5rNRwebzIOrBondm7M9ejGRWycC5GZ0jF+u3d1qXp9HK
5AazEvOaB/Py8PsYuEnpxG8ZAnLgEoF4InxqZL8y5A9VryHWGdM5zsg5RRJyuQmZQFLylaDKNeim
No7zNbqn9TS7Ch80cqF7tqArZf6iVdp5xTpV5MXcD/yAHs6Xcu+azV5qEDsd7sUvq8CEgu08Wsz0
SPBI9C3M/jFQqc0fJR1Fg01pwUMOJZdzRfeHFtZZiHmWbmRmcs7m76gtDE+k76Z0z7IJXRO/UH8Q
ZjxGPI5Mdm+jgDmKJFjtwjnWqAsTaWjgbiGjX0Qba/P1qpKFdle8ZMZGx7pA1zF8tHbz+4SV+o2f
NJoj0MUXrVH2+9PsZHNMJh/C3ti/GU6/Tjprl42Fbf/65TuBAKKGFOdFM9WX+s9Q7NKjDe5triJ4
Phg414DhQIVoKOeALNHr9XfzlEyYsY8S+zQ0JzkeYpR94EiJC6iHIFzcuO70uhy2SPTpu0kf0E6s
zUdtXvJyZ6BcAQQP2f7C4XBpzR27DsVZkjIfsJxi2hytrUl3iP5y6kKlj+DLd5lRxikgpR2g38kc
UCGlVgMkBhWzMVYP+chGUCEmX6/FxOr4zI+Sy26TqbBERTkXXLuMW5h5GnpRlpLyQpQBIJeKbdDC
pmtSH6bINEV54q3sxZ7NMsFpiK5VxBG5Fxjq65Q2Yor9TFRjEq1G5rr4Vp+GuAkxbXnKOXW7pL9M
ovLqd4WFtiJoO4ss6YLa+EnuIIP6RsSeY/NXU6Dd6EGqVKEyrBxv2cvkbPbzahBKh50mrhXOKOOJ
52PCdQ24gWoXgTcpyUvMXn+eJ80DYx7KhG5/8J1k7gimUYspHORfF+pPU6ZDNOLyKwbDsLXGhPSA
ntcQicCcUqygSTCYlGuqn1gUVSPY3m8BD1Q1bjtFvrxfOZDBmbwdGK+tnghCrHOxqpuP1yxC0l3i
DWLXtmZfcawhdxW971mM7osQ1po1NFhGeYRkdNYQrbadWq4yEmZQ7UpyHHhExANvBS1J9169R8rz
x6UZLAPR409kIwBDzSZvOqoQXgz8REe1MiH4+9r27WBm7Qd6kknJ/lPPc3rmrCdNr8WHww/CgpdP
JMMXGIS58zwLkYl1++S7iJygq79vzRI1JM/OvjtVR+rrfkbVLGMMkYRt7mw4hAKACpBHpB6dOcty
L80m9AUGIn6NfeWWF7VjMTpQawpTIKKDy+QZQjdEYiCx8PlfWbVbNpo61AJKhGfEoUC0uiLOqMW2
tZJ3KHDXB85hj982F6lN0yoCnfxz3dcrheOb8d5+cCU2SjTAFBsGmfObYShY6yjTGrZoCxi7PUBs
foAtLnCZgw6MA+zNnHK7qLEkh4s7rUoXh/pbUlbWTPsLTLlTtGoxlgH6E28ptYZRcQbm8rJTny8m
7uo1KNtDXeK5kxL2pQpXrnF5tRy6kN9Oux8GgXjtjegD8K/uESrp2vsdB8HEgpAb51S2SWmkMNtr
2sl9CT2k80jlbHyUyeQ9D+KvX18tv/8TXigC/wFo3aBg+nXZE4QUxnp4OhnGbH/z3zf7uYGwhtEX
w2vsAvcDKwIPo1GSfblLjKTZJvVNfels0CTcV6YnC4I8T97skIIGUQi1KlVlNj70Ufo3LGV9bIbb
Gz2nkH0p48GkKKNc8MissaJm3SrGdk5VYgS4Jo6Un0UCvwNspLMW35eXwFdylmnDCAuNMcsWvGbE
+R/vQDAoDY4tiHA+ezO5vLiDxAEcX+tm+ots00HiHUQNNyO0h5jBQrSvcGoFOnQ2wjVSLJ9quvMU
hzw+4UGxtIeIY/v9lw/mmUc4f6S9AYqIVGu7gCW/CWbbD7KeWqIIeISqMczkhgPSCIhaW6i7JvoV
WiqyFm28DkjfyfQH6ovf5fZp7rIuJmBPMWMq3u7xaAiuGOSeAOUT1U/htz1te6npP+IcOb2vquGJ
eEilHXJM8slafARPxgaGSSPfOUIy0r/qSOMyn9WLgXV8//yT42CGFJsVpwayiZB8e9qbPi4eFFp+
KNFWUzc5HJWcO0gsiLxNxVm9tDuEbKFUY3bpXfT05V379/w69MqHOI3zQdidcUNv+zXUFRlKqGPT
eY12xYFMWsbP9sPVK/4kz0yLmHGK9tPXsUp4vkE9wimgF8XUoLjzntAydiYvszpLQjQi3YjGC7R8
dD6zEZoS1pfYfI54OqaeNLgitlU1tCiexq+dFNT3ZXmYIBJ3c97FiSUe/KQEdBgF05hZO09S4KbM
HQGxQGwUHNdPxtD8agwUiImFWtBS0yxZmhw1qoQ2b074fFWPJzcs9ZAwP2Aob5oIkv1lIm3YxxzX
pSt3sJoiDcH0aILjkgwFtakJuDXyovaEmP5hn18wQgh5BVXr9P+7eiurADwkJNLPfbgVXLmXJKp4
0WWL1CjPA1P6DUsKY3677xZs/CKndFDY92F3nLmjTctHfH66HNRR+2cwQMkQQ6bgKenff94hLMdm
FL96w4HusN9ZtCJkC1bxmZLbexAArgfz1nrsmu/kheODh+TvUhyUHsPcxZY9RbilS+pmBjWaQEh3
GMZTEuay8QpD1gC6XA6j9G0ZwbTpZrP7IbN2ewerY/ZZ6cG2YQpsLEPvcmuJD1wPlyFBHbjgUZAX
MBgYU7K0FH1ChzPOnNJ0eHkMehMT515Ne6o6XpKrJDoXSWlSgGgNHvq+GR+AWYbAZCxpLWlFLGaF
I3AxbyGjqpXKFPbT62K80E++Bj8F+i37pHN+J7CpcR2R/1YpK4wfwiy3Pcp+1wa1QqYrrLlTQScG
cV1lP5QUQzl0vEWreMvig92udzoGdpRYGkHs9PSW/4OHlhEE73G6LlIWXHFRNcHXyrZO+kdw49di
/f5EOgQrUeXpSqmquR7/FSioVi+6B3cVTFf/saZjCrXxHOxLQnZeqO8aYQeMQzqp3VL02b+6AKF/
5Sxzn1hC1us4EEdaxqazZJjnawur/hQep9I4IG0SECe0JWq/AdaU8C1M5aXxsCYkUKY1uaWw33Fk
0vUahjU4GOHKwJS5PdnxTzXFskJU5p/aV6RvFdJIr0fpG0pHUHpktZiOp82vggs/4UWR3uPwxPEY
Eb8cDiBv+1K3Fa1uOyQD4BFf/dFpubRJOxBp038vgUdNjsORWo97ofiUu2T3N/JuJ60eTBjDsTUK
JkvMWmuvvyBaF1T/vWyNRxKxCRiu676lWUJFu9hhZaW9+EynIiDhLBMLGqo53XemIT8Z2JjdG2nZ
YWRIomySMFLUXRxOKAZKiCqITe9QvlM1sc0aNmfvJzvhsukmVuxtTF5tEWeGmdctB5C+wYSPPlbW
/j1sHrlriR/mtKoR5Q75Sjqbt6b9K0Z9WbB/9LWzAe5QxhxSvSW7G4vTZVb+EWkF+nKHHGIQS7dv
zJwXEOo0orogZGasnipln6cV5kCFVE2Dnbur3X+z/YEiLAth7hb5iS2Q+7TO8lncTNvCy2FZE7ab
zAmgCj5LYbBG+NpgM2SeRm+cbVvELjJNJRTQAgfhRLU2Nc/TVN8vNwW+WXovVrSOfTfbHnc/3D4k
Hq4Wr+C3jn2lOmddt9yxOm/2t6hs2mMcpniPVtW/3NfAKMGUvqJtOm8WXCjRSun0ktH/KjczY6vO
Od+c7LBmlg6Dmp1psY2L2yyPg7/k5igpT31iylZADTh3GRRemiYsYr892mc0bWgIAhjSbMt6nE9H
lLmAvy0+9eej8kNAonh5kc9S54z5rwBVrpvjLk8MvB6DsUkvxHFTIytnJ/b9a3A/A44GAFF8tqAk
k8NXHOcALjr4b8CVl7Qn1yZmGSKl7onm/GHAQQAkVHNgOsl3TyixgxxV62Px9TAOmdaCzLGfd9kr
1wzvy6ftU8G27tV45Lv6xPIAePz8bWWWG2qdNkORIdjyBVoZos/J7yGHdE6dtKfAyXqYuyFvC8m+
LZdnnBcoqf0OD7zTEJuawUvNPls3Qs0hGKMjRzlTfrf/sM53SWLAUmN/erVbCNDvf2GNHN4imR8U
7JFPw0ezfEoFF9k5wKe43iLBdTduEeO9O/smVkHHIBLfV6E7G24Oro9hLC0nxXphH9cgdooVfLex
+pA8ARUgn8JUvctemlisje0SAjDBjfkG57bvEge49TfuWrRLaqyptJaHR6VO7qoRbZxJdcZE1vEj
pT0ane1dSFWCyngt2rtW7fkzA2+Qt6rL2h02zQ7l+YEf8zNypIFQ5+IVWM5YBVxwrA4IzjZ8LleD
uRv0437Cc7A9OiogrfgRML81uLLDnNJI3i6auSSjNHYgqYSjJh07duOpeu6I97TL05HaoSnGIN8j
i5nFyURQZ6vWKPeQN7YhVqkOPK4AhG6jbdO+hZds1LUt+CJ17+pH9+9w1THGuKO56qksEMlZzyEI
dBsjxd0jWdjC8al5srLxoQNMPP9NSQ9295PxpOksHsBNcnri4ptJKXIbR0esKpbljBxshz5AE2hg
FvZF+tyCIiGo63BefuFUQz8jvWwyjvopJ3L984rTRgOWmKmCJKQZjQgo2OzNoQSgaodE7WMoEnFe
B3SO4dbkOyqTlKSSzq5FDUUABIebrp0IjT6biWC74a97Bl8erQEQqsZ+R+60LZJbdcfQqdms27R3
pqOFDKTL4/XOFVEO8wLCuJl/zztIR/fZE4pHHd7xULbxKtheE3ZP1fIRQERt1Hey3Rw2/eJErLQH
TIJ0vnQNrasyR49PynX48w18NhOw6Lzmt+wuyDwa27byz7bOtX8u3hix17Vgem8RuelxrDmxTFXy
oPZf5eXAtN1K78jr+PQfwkVEYtN/7A1EF9iP1Ah+ylZY3c26X77g7SscMVsXYr/DY0U6pCC6s3Sq
x/1vaOob6HSi4eXpmuRc9UGLWWWKkDmniMn/OUPgHjFz8Wh69Prs1ia2O0gu0Gi3/5gAaclzfPOX
ByvLzCqM2Yn6WAhQe36z/RmTOFLKoiL69P7KZciMr1Z8GvNrvIdN81/+O7gDtZBXfBgnW1MhESNT
JUfpU2mRWnLjVVB4HtROneD607PeosqqRGizvDL6xAzqHZFXSGFfccw8O0DWNa7Dm6m+svFV9N7/
DfJxpHur45i51lUhIi5ztpGmQQFMbWGDU4AfJNo84lLAhH82H0MELIxsbCFvNTXFPSkynz5/V79L
l/hoT0i/C5TZc6F/Pqh/aCn3ZnXeiRIh0vvsf9jCWbNDuYeINATTqkiCn6sO5bqLM7N5nAKSqHkU
vefO2NxzXiX7QRHBpcrGWWpKHRDJCvHuucwMWft/oXXJ7LdP38YbTUaVg+0jz44dPcab0t5wOGr0
ojIo5XLbGzb8Za1A36yt0WBu6YBZQe8dN+P8oS+ID9dvQhNTpI9FN3TL0Mg1kautVQD6thWJ0ajy
CcR7CMx/BicBRDfV3dGKWMR+A2/aOyzHiQeK8OPsgQg5AGxOMCaMb5FfqyARJ4wptuVfvom11V5u
SR/7b6jfuchQtBquwJ1ai59j5ZAXMtZ/vwnCcKOvxVeOfQTZqIMKpU5wz/6ImrwCjGkq9gJCHttb
qFFYRq/JfmgqKaRwx/Ui7xz6rulirnxxqSMOnkn+WGSOjg7XtpxatPKLY/4GsK471P/WHGfe9cMG
1WR8YqbRG1Uo66xa0KHkI38Cg7FuKV2PmwP0iZVG1LRTApIeDd24l73G7UsIJlkIg1PhtK5LavSS
QN7/1lrvgRXP7TWDtGCmRyfMWv0b6AayikYJpK7ALMh6tgKxNpLSyzkrMv8+G1I6BNVKHu0c7ZYI
lX4zAG9C5lU17nVCw63btQXTEAo/mFEj5gXvC7KlAQBeqKe8XzPfT6qauRoz9q0yG4dMG2e8uoCk
IXZqlaHbwC6sfhHSPP1aV3Kra51uTRaR/1Dg3L8nMEazL1YClRFnhGBJ4CFcTxrb4I/GM9/IOQdw
wItQCDji39vB+ymt3ewFG10jK+HeBYaQoqlYVYXqW8fmk54zorFG4OiP5+0dglglQ260nFtNXOZg
Awtr7n6KXmb2E4gFY2X0OcVXGPmPoHDXnFIe+HmAvb0UYbNZkXj62ZPEHAJySu2Qi1MiVXZk2F3P
CwIYErRTZyErV/VYZcYf3HW2Z9tAH0wuk8Mg+TyulinX5G7KkBF4BIM0v9z0gf+ExnGPnMmX0ENF
qQwpqj0c6KYSTTTEfjgzQJMRxlS3e68aCPFgnkq4UYq0iY+PYBHJk23hLBb0D4C0/PLr8pRGIGrp
NPEnqmcIGQMWW/p/VybcjMDdifkySLi1F92giQ8rGmCyO3hvGrf3lDiF8oe0ZJfyjbi9BGTdhXV8
S5WnHK3I8tFL+JBZJYCiUcI0zp7n/2lLmKXBYBUcUADqUNQcAmlbFPD2pB5DKb1WEGrnrycC4A7U
W7Jt860qe4j2OIZMbV7izypcdA8oUTK/R2imgn625GJI8EZLbAczX1FnHcMrr843z6KWURf4wpri
fcNrPeSQUWcDDGrH9epxEzTy85pyervwx7Pd+dpx15dvBnqbDl4mbhYp6sZtwntb9b3jbtgLg3WO
CAzS5Q915Abgm1bWdcWYJjq7pMdEM+6K34jqT2FBwXsQpOkuQbjWhvHnXbYLMzqPoA49zMhUPo8V
u4gtpLm8e/kF27oDaBWJe+1infl9HWTrRtOYz9NE50IS3pMFowLq2ggse2qw1WnqaIqOJf7bbUfV
PzZ9VtuvBEnBseynbmsD6Bx6z+MVE0b/368oQLUhpquoZ1leLxsiHcgo1AmmQ5T8abepxUkIkB7I
fwG0zxSQ/qnPTYpl7Ebvcfr3xIXLFRhL+KkC8J5fjHJyge04bmXniLveM16uPjLrg0kpmhbtgXqW
8KsyULqyPQc5cQYHJ6052jr8VtlvV0k0WCZ+UwrF50lqNMx93tbJbiZv11+iLdrm22b3pCN6Q4+p
XrHsqqGjZXcGPDcaoLRx86nVCwYEgfxrAwem60xUudlP39vum5AVTuOEXsIf5G7O/L5cvHYgX7e6
/ktQ+Fr2ScbUi1tOLOmluhn6EwHFkzl5vdLWMkRDAMF1tPdPmIoCmukbxnDNXjHyBPhFtTs7bEwK
4zGMvdv3chPuqgMkj8+C9zhHsOdaKrnshw6T9Z+BD/xf8Cf6ODcP6MOe8UmvRtIrMuPGO+pvs/8D
OUihoCjTiq02DJ56rz2qiFMRLZLXY9FiaoRyBy1ch2LBL4F4upc1X+er/H7UNnMlJF1ilw0LoPik
qArjlzsgbhr27k6dp3ZWKq8b+Pdt/I8Li+b5G71Xe3wf9havXvrr3S6FM9wg/zF+/gk4es1WMoay
gMfS5z6bWtTTstaGtBR9QzPcsu59G7oygKcr4Fr2hg22TNYuYvEzII4JSt0Hv+9eiOv4T3Jat5HJ
+RQsxx/tSv8Q6fcqnIKF8gxc+tbSmdk0ZYf9TiZjJV66Io7NRJMooWQmemEjap7gD13qXz5jFLr0
6WyzSsFqrXNlt0wuWazfM+4/DSHcZgF91VWElh+dmwPZpldSrYYI+9rx3JbH+2SNK9GdcIwJpMBP
TDQo3jOzd5iRwAwOX0O78fGkTTQaHMKnP768l8yQJB3XNWwQF1QYIac3MTZy8ab0Dv0quNyM8EEz
zQ44mDIY7WFCZBzPfsKbZyxr93/FD9/unqh4RrHWoo1zcCeK3eliXPloqadLTtsxj5K2+qFMIljZ
Lx5mclTGhogAfFkbkluZPpBHcoc1vwtJiXZaKJe0mgEtTOdZ57QnNwccpNzPYbzLRsxqFl/ZGm9C
qerkcaQUeOjHf//bHkshak+EUNy4LzkHnvlkng8ub68xiWeyEk5lsTrN4q6BFmXILf/YqiFSkTNX
OFoScsBqpXfGNcO9wTt4a8dX6wi8EJSldfTlQB8F55/Ez4QzEXrkheNKO35wcUxElc4txLLznCKT
3gb2VFLzCjPXnZHk6FH6SHQThQsCjBrLCOrYWcVnhR4wEjr4F9thBlwyVAnq0m7aZRfCdQKwBKxY
xu/53ha9SG0g9S94whg4ZUK2uJLXQO9ugvhuQY+tM6A7eRxOIUXPhMOsUQQK5ITZytP1qlC0VXDu
jO5sDAY4YFZvs5lWPhhPSPcqxfVACu4UCzQkH6e4iqxxZvlcE1FFq2ORlUz+LjiyXgQ+oAOSWs4o
tE1GaGzY5cMomtOJyf69uPX6833TJnsKPiwbmloFawJPSl4VetMsh54G8UoDzsE22xLtst2fZqWS
tbg1rhpcb5hyHDnd93jFK5cM0fQYR2hO+MB7UUm7KG5RwVYopNv6XBVbsUClEVHzHvY2DzkUg+hA
IIAL7vCvsSHAsS/LAtc3yZBFrqUCVb4m7swGh46rlv6mscKdVe65IwJJPQyvxEbH1ekSyLW0z0Bn
9VaueaDC+A5RmGc/J8exZ10MVYyM/Q5DZRCak1qVtEDeTujPUBM1EGDK/Uq8Or8O5sN0SW3QEi78
/fD3k9B8U8VWPCzHOUmxfhpNAz/hJo2dYjgn61LSU5fFjZscLA3uQwU6EqreJSh5gxitaie37dOK
1MxaG7kAUT+AWwap4k2TZ/hFz/2iQL42KpKRUBhXuFUaKGMI9BR6m8lmlwFD9tJyqIyzMrd9keeZ
3N7EDUntaNbf/H4vUscDxlwOG2iNR/PGsFF/4qKINBMIzEFqVYua3jFS1gw9fXqaJtD7I0kSSzGj
MZz2kfy7U5FCyVWedUcpep1lVn0MQPyNHsxW4eTKYQb2XVghaLIIZ+aOMte54uMSdhbvzC9Sf8Sj
xLxGikSy24NhmrP66D5sdD96GnFcOTri94g24UzdGfwFhTHkF1O1x5ot6g/MzfwNNFU3Ds9edgE6
O0FnoLgtR5sQ1iwy1FSCnDy+OykQUegd8Xrci0TW4Up9TNHQwiCZ+jtN6PHq1EmF4Y6hxUvKkP5n
vMZSa3tLm5oxd6eB9I+vjaMzxwRNCwKDJhmuXvaGPqLJLHlbLFucTtzLaNmIG7/cfXxaTBz2MMjf
9aKPewQYvYWUKzw0h+owfjKE5yXBSHnfzDjMDWKjG0nu4YACiTcaoUzhRWCD7v7S6Nz3hX5LaupW
e2YUrqqIxPGAq42FrwSBkXLBTVU4ukvycM3cy3eU8HsozOlGZsFRlEHvL1gJuaaezcwBKeyilU8R
C5yMN9C2QOBiM1RGUZ8p5UDkRDDS15CDUAK/ya2400D9tZXsA1bAMUXc2Zmt4lLmM+ccEp9HtpN/
tDZ+HsugwQZgO58ONlfq9828NKHZv5Qq8c/xr7RXyvuWhmXtzFbcQKhyA8cIeRjsQ1XDDJNsGiPp
ZSanhip0Tif7354huF4e3sQ8hETwbXKeCA5oqvr/QYnFX8Ch7lxfug3lXTQoXmmYXTe2gyBDKCnf
58wXLMe6SQGMzvFM/+sPwb4fPvBJYB+o7F5Lm1P+q1zzPWjXn6faX0Jq4V+nBG5avVHUHUIQGjhN
r3265OzTjijlZHTSsATHR8SdU1I90CLwUQSB/tHkBP+1byvbkiVGCeSmci8wQKjv4F2+Ya8882Ug
zKEqzRJSV6Hq0OZo6n4vi9nVVKTtlr14ABzoaV8pubLVGXN3KwTA3nJyX85Z+SRq9oIZVoeBVGz1
cJq57XXsHnlPdY11j6MFJXZql2KxJ+f8G8JHWZFLYaX3sE0U5UhKiZvLWzpQiOxSGQElPoEYz8CM
m/fzqsb0NwvmGJmAhdSLLRvO3+Ao/3n9UBO8w0EtFVGMcsqyaCD0VIIsTsZSWzhC824TmS54zD8K
gLhqKtfChzkcm9JiIQkgrFuBnO5x9olm+LaQU2g+xomUrvejdHGAZONgLA3Ee/wjeXWebtj3P4Gc
2QL8ABRYbFbdoFqrmH7cCuAT+BRCDkNvYl5jsDr8hhauo1QcAQ==
`protect end_protected
