`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FPSwcxcmOLJFNKau5DcetstBfEQDoKQLOTxjau5lYgEKTmMgOSCOvQ20FqMLGf8dZP/J5Wt3OW5z
5fMGqF7yaw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tYqhegLt6opNQm61Pvqsd44qn+u1QgkiH8DITWCOWym1nuWJVR78tVGmEAM/27S8uRToN7MO0tBv
gNiOO8hhYjq60OoT2rkjLBpiQIS9awMrgkM/g9AVDIqByrE7/KdbOrRWZYnewdORM2ZjgnFgKD7v
hZeDGdwcHKxWU9ksMRU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K+gYHLvBXWBkT+4rkDvohiS5NTCz3zOA44LmuM5EpjzfyR9llufo2R1RSSoZoxhYPx0Nhnb9IZeI
46Hw4uFilD8k2RQ9m2epoxBUZd8a7Y6VyYjTRXOklLkHHhWgyAFD5zPGB6L0NBF7xVNK3dmv6TLe
gr6lbuKAyUvgXszHbyk0lCWsI+h6xdp9jTrzTQTAFV03xpmJ3EmjKYuHgqjzyaeaLWZuBiQhn0L2
SAnzhfhoX1D7Kb/ipH0ruS+KIlbKo4NMunkuU+BTsJj2Vcot0ebAsl46VYrW1cZRiaY2QEV+ZhaJ
zz16F8ZKL1LgOlKt0Ygu+HaayBZM7waFGCIoCg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ISStRpWhjpuNWr8InQEt8YuXaDvG5lwe7CbQBZXpizKf4bNdEJR82NZxFJvzsM9Q4yd2A5a724JD
sub9BzYKd6GfYGf8wZGbiYXx9IaYrZgVpRCPzo43JvZ4GDPyR6XCQgGLeQT6pNoccJL2FMOaFZN0
dayJvcxH/xwBLvg4gvEd46Uu6A+mcMkKOM6I1sr/WTAR9CHf590SD2/dl5sbVEMsQC7356WJapoN
F4P0aNjkHRtJR2zC8je5G0Y2aAcX9zGcUw8L15glLYrvSqqSq2mBMDxv/1jUoWHT6Y2RPtFYogQa
ufTsC1KKyWLBdiOlof8eBesoJygQBaPzZqvlwA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g+45qipZLNCcJNgGPTHT2CwrWJuY8S902czIUqwfWS0NVR42PSDoXOfZG4yx6Zc1sITk5drO11tq
QOJvcyKRGRJFOh1dsdHThLrjwcxoXzI8B0a5SK3x1o9O5Nv5m3oaCa5oEycuS3hgGfhWPqnqkI/e
9Q+f143/UxQ9k7HBlL+RYZk4OFZJPcZh31J6/p0uvjL454h+CvBuoqDW6Nr9YDdsdrN4KysqXwxJ
c0nvVc3VS/EyzFcydCWVY0zwBdJuR1xbDapTQNTPCkx2Jf4a0sechsW9zaXdVqh6TgQlDKhC0T6l
qTYQ7sPM6FpeLIbP2mEelg6QeMv3MdzQi428vg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oq8hJo4ytcxLOjTf7Ft83G9Ds4H1FkCSGjiygy04a5rE5PpbUxmFmdpbBaNyOSok7VXlLuaa/ctg
PlC7mjfck8MXqOG89JK6oIYsjU3J2ditwlCwcfiVvBACguZKUYo3OJ5POpitRZYUt4foTZrdbpDQ
4VDwl0Q5E+qW8y/mGxg=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfxuWhuH4lzWzeqJCdiPX+JCRAFQPCPmOgm2pDMK31urjoFVyt3cxOgHJRj9lwiq5L6CL0nKB2jU
WacmKzjj+L1pX7wmKhPhmjG/3Dxp2fur/a8gVbTg8BQneyZ3g+J30lauE6XIf1KnXUxCac++kRBr
3qXgCk8rrxbkKTI306HK6CzMcMuygoubtvyiLVD6Rol7QBiUZnOrR4o9z5ZlixBd3iQPjuhqtlJ6
l3xc6dQGX68GPkoeXtX+PjodSpsEkK7JWrGzkFBFz2Q7iX+JAa3Rve24MmqbOM8Fjn3VRpyDf+Bn
UUlhfBpxpr6D8Br/wz+KmoZXN0a2yRXdLg8IrA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214096)
`protect data_block
9C2CJVAeTEQQ2qJrQ7jR0KT4qowM1zSr762DIls1JMZWA1BtrXegfBTFXFCXDJXRWbrzN9Br1kSy
ToB4qI/NArscTAJAfbbue30i4MegWn4oUyzbD3SQZpOSouJI6CA249lk3L9Zy/46KuZeZZkStWgf
wf/AiIc2/RA7Jm3qJanTyG9f1li5z34+w7jrGDhepwO/oRAABNADlwzv0KJmg1mpGPmHA2mrmEJY
0bLwgl156YEFm4VkEqHYMLiFu7U3Twu1VYxtrfEOW/fwTxaDrccQDN6UGG6x1f3s7E2grsCBkyPR
VW7+puk47BDDqf5QB4Q35hO5b9dglIO65zUzh/fJLtpiKoclRapgkQO0b0iEBACOB3AIiZB73Fae
SC9RpaERQN5Y8ZTlQZsju8+35NNPwjcK0r+hbudxDL3v4pDYgc/qRtrwtfCURFFJ4nK8mDDk7Y6r
3jNCSi7maUf8KPWVGBejy1mlIlb8Cq0hScKZnlNjhWP9xURBLnOUOwV3rnhcWJEp5Js17BbbPPul
eKnuM4eTn7JnS7CJ1YiUuBxfguY76d/JW4kIqvHGaUXE1iLA10yNP3lJ9WrjH6tpgq5aNaaNMRtY
xsudEX/dy46g2z7/Dhm0Qwosdv+wB95mi/TE5zew2tNUIaodhSesmucocUatPq4BViBe15wCdcBP
3neJZkO1XI6Iyjs+XaufCdwKh9FSMt9KwG4zkN05+6MTTHs7CkX5WG97Vd5pVA+HON4f1u8bIhSt
+oSwYscHG8Q9sWeK9zyQSQvjIBNl1TDfp41AiUZ2yLDlW/AvVkvhyZJZrEeECpslLCfEo3ccdSEs
EzDOVTOI3lzbAc+hUTQl1NT8DqMMErxtLSG0vDOpUCGwzLJnBsO5S/ApLyMm0adblpSbyLKS8dhX
gH58n5igZSZBbWq6glHm9wj+Qkdw75/StGlayn/Iz9mYFKSMMlfSTJn0WQoptFsJSyeW25kZbqrX
aB0WoTER3QP3U33s8vjUW5htIPB03PLu3HVoYWhEnwgEfRH2IUVAujfwQ1otQuetlD50SPUmCgSC
9jlkzfjL4C/eV8H9t4VRDSFKgA33IC2QOqGmATj794iMoGPlv0lT8E7taCPilzOOFgemtQbIgU7V
BMaI2yWVWzxo6HIohc7ez/kMpph0p/sndbhG8TXJKF9B8bDpP//63E5dkmZb+1bhP+N+Ui36Dq12
mNhzemAOc6RyXbB9ODHoRsD5jVeWPD+5pHuHSxanjJhm5ofA86A2PKRqcbPbFtZVjL6FG6U0aLRL
VIn3AqbDFXm4npKexid8zJ6ZVWSv52IbHULqCk5HANFnZ02n0j9xD/dLm7YJJTYjSQXNMsU1dX4F
+a+xaT+OkDlAaXK7ppvkzpKB7ZF7nmb4qrcwOJd1A74E7ameCenEqWSBkpkCEPJPl39IoLiZ5oPZ
S4pV23T2JQwOyPccDCYLDlkP7ORqwBBN96tEZWSsBuL8YtXEgh9pLb+pfpLyKkQDIt5iSLG149l1
01Uv/tIQ9gd3cKGKYKC1No1kHxo3r/7r1gK041dleRvVqiRVUSzPpz3aS5olB7t0rRTwGFIdGB1K
eb2JZAfl8NEy0lGxZMYelxYbOLys6osf9JoERSafAE8+NPlTaV/HHLCaSssodngvIC4tUp4a7W/7
xtg9S9daaZTqI09ZpfNggdPV/TmSokTkgiRzG2yOrxbywNwydK8Us0QO/B4aaCUeSi951tcYTBo5
1P8oGY7l5Jy8e+Wdq256Uci00pwNCy6cBkcF5Jgzvk5S7PzKzDWom4LLCRzVZuUzVbXKH43I/ZO3
1+UP4VW/xemYdPTAiFc3BNlkVIYttLxsvZee84zIjgZlyI2Z+yP+mxF+yv9MuSEKVm4brKwQSUyb
bZwfNoGcqElxS8KHANTJLbYSfaljq5SF6Q5nLvEtiDC45Dax4HS1cBVj5VKxnExIItbDzHyxbHRe
nHdeDuAMy7NWGBnTycxATIFqTUTnPZ3YxIMgGsqHyMRbXRC+OtjO6hFb6gVnfdq+R5aT5jJT3yQL
AnHDvD/1hUVr8sk7VzNvqY72h7gjFA/uTeGwp9btJbNF+t7fYEVkCddebUswLByzMr6zJleZ6KUV
8XsGQ31VJdKMYHRqCCh1WEk1goJJ9mK0kSoyvMXzXmXsnbgP+CctXszbAHSugS2kpdr8lib7ozTr
14b/kmXDNrzmdnyJCLORB05iXOYWPwf/9EGWXJql5AneAGGQkEXmvxhR13eoiU3DxIKQwmdyvuib
x8v5KjzS9xNvWbe7OPxmXa4q+zNYEajvQGZvqB6TfiSoVSK7dgBkZ0KQSL05kSuu9nmxb/ABPdZX
wvGPuB27q4dJ+ykBQb7881cJCgU/l8RUcy9hKtPF1cd46QFhvqUsZ+2AxH3IWuvVSBXgK2K6S+pr
QscRnM5lnYH43ziFNaUPZbehX3XNLsLDz+32dTA2eU/dArwTxEsnBIct4VrZiV2KYzPQ1oJRglfx
73t0x9R97VDB5EcKzLoQ43m48cWH17GOZ3E/CV7OnCOVyihtYNueX5+SJH7b+RoQJC6Qgn9joTVA
1fFsHjd2D9PF9Ua6RbrhldUrBBy9LslWCOjsqhYAaTVDRrUkS2Rj0A/xkMm9agT26ftdIVHbebdK
A3jePpuJkhs7/9sdXviYPAgBnAiDVfchu9LZSEIxFZHjyokrQubqTlyNKMMdBrSFg9jrroYkW3A7
23EpbR+VzCi/G+gaxt8/bcwm+MVSnZ9Mo8nZOxrl0AXzwPMtJvywe9Z6O2gDkwgvvuUrnqA7nNNU
6s2ii+SzenYkLmKZelK8LV57K+Ewuxr+eb/Z0hjMtOZo0qZFCbKraBhlNaaMbfCZ3DBfWZ//BQLo
OSR3fWxHpEzJ1OT9xoJZC9AC8xT77wTdZlM7HS3awFcoapSoOE1FOY86UKldkURDqejXEn7FFVFU
YfzIjbNhT0cTHjUDo/xvnatggpElYcopGl8/G8/ohO/IaAyOUW9zsX+PlGcN8F+0eEozHQf81JEo
0wgg1QJhycz/fa9/M0jB2HAmHJYI5+W0HEyCDpw6vvPlvKSbTQp0lleV0z2uO4A72E9kgYWQwiR8
ocVwe9FQdCwmcAcsfzBYurlXQLwyudl/dKXR+ApPUmc2IsqYk57fzF1qsa7OXP1S+ywxeJQFr9m4
h7x66h5376IZQE3xSHbr2IIrNP9s0uOo6jKB+Jwf2XvLHR0yeqOHucrKhQeXj/hl2VEPnn1ycUOr
QywUzxRn+DovGXjvezgT0/HuqGIkkNKvDrdBzsQQCpkmGVB3vpi2aHmz6F00BPqEJ1p3lOukXN4E
x6tg84RnM68AXfbkYgNfcol3D+gXtErgwMKgJrZSd072W9jC3/lp1Tzq4swjtdE5aisnZcgVCPSj
drlHNjGnZ15xFAGjNggazwtiX6CE72/aXGxmwykCXM+rtRJca2uBei3U44AwLPZhR5nuzKOOdcgB
bx02wFEMRdRnHrF6AJmhXRm7QsEqCoWH19lBAbds8odSDPcdFkHDzgkzsa82rpbCqfKemzusJPt7
aWcEMqvrwJgISaHsazjneZMf+f5My7Ac8tQbFjSwH1fJ1i/DmM+tHrE4ip6LPQ/sG2N9V+1JWuZv
Z4fmzw46m4wwqlbNBuNiScVk58nWzkSyIbD2kLrJ9tX7y4kTLtuzwWMmPSpbbMKI3oehOOfigV1e
n54nEMcV0Agca9t1lB/BR6fsjHuGUw6W50g4pQaV/xnBiEsKGIO5hYDFqcS5jp3GAIWVKacBW5GI
RxroNcas80PWPMKaTvIFusNmkFiw9l7lW7LlPmiz4g/wP0HyyilenUIEFoCFfWXOhq2utVh8YFuN
Trin2vUfHPYsSm3z5MAw5KgG5yLTf6T6u4qFVonhi73UaPHntQEZYfXfa8lsSdOx/YNCzF1Lr21T
+tWsXtKhyNEkend0kjORg8AcnfI7XuUhnEDTkLXUkjoTqrEW51sjKoVjSGn8rrZCYULCN5gWxp7n
1w/UPLAfCG07pMk7dyodQG5jQ4z9QVbA6clT084ZT0oW6nx8vLPajY5s7h7uYugN+Be1s4aYTy+a
JSsmTu2McUZCtRjLWwzJA3YTNpbaYC7kJH2yaAKhmeGTwRJSvr8viR3WdbWGj2cFvy5bU2rpZOfL
W7vGlYyDahjCZBSuJM2ANptvuirXUTZ3tH/7cUOY8XFstvFo1lTR8gBrJzWWyuWZm87rnqfOCJeo
oBlEdyOV0zHBg083C14T5nzT9+ZFslIrlC7eyM6QGcovByP4a69VptReU0xCTOgPMQ8mNbb6X7kE
EN9brM+Jt6OyWCvrMRwnhq4Ha8GTZs/a20xQPsogv1DsjxQ5PSsvwedgGIRAzTM+kVy67YunPnhT
ckroyzV58o8S56xqoRWaTDhkLR99uXyjkfbeHR+PF5Bt+QIWs5pcjERwLLoWWKgVoPuEzQxdTIFc
tlHrlM4johxr6ylbdURPwMAGGGsfhyM/iXzuTWrHnxpEymNPi7724Eurlp5pexDx1DYZTUuWZwYf
VuW7aTd+GhOZteRA77X4pRml+lLFDsB/AUlXrB5tjtMU2DXCPn8ztxiMRJjWgixoOj/bdRQAuD6a
K0eDxOuAuIkThED2eUJjuxXxjkpTP/ETarTZMFhod4jzCYL13jYHYfQA+U6Yur2DFsD/JXSfAH8r
poWnAX1J9wlE40Td8bzK3L0/Rx0I1zWB3MbEhitEnAAB+BL4jOivChIsSCFNAG0/K36bIzqRgbql
qPe7cyvomrRI8RZf1Tz17WvUOGMGIZUWheUbF3zNYHQ1Yo4EfgkgGxP4DBOIo68YZ6oe3NvvOSwv
aw2B5ymdrmsg47XDqWuobX3Qin/eAjDitNy2b8MzBontnGJJ0WdktxxhyXUk8cQmAp4cU+85TgAG
dyTnTyJKe4hYKk/UUoM8Ps99ojhhLOZRWZ+l2KuAeZD3OJ//ZascYGBb/w0BiUcvJTmSdOPnIXnI
uqYvNqErYkkiwEF7Z+RqlBs2MVL9EWFVklpMQm54gabhz4gdGz+t+c8KHMXuPN0ul7bHESJ5F0EQ
gj1qqwdT2aYSN/xI8Mw1l7ys/xRtAwk0Dz5g2zcDv+G/HBM/mU4NWKFpUq5Vmi1L22bova8SryVI
o5+FxBOzwTpUIKFoz8K9Mn6TDW+11bflfFmE+T2fzRuwrT6sUeZ/aZ/tFT1OlyyQFI0fLlsc77QD
9LYKWuaCVkNja+mGXKM/CS0TUdRhR3lE1M0DSkNblgrJ3IHeFH1elrAcGNKv3GEco4JRpuwf6cPM
Gqh/HsjGzYhp8YIOEbNvQR2NVheVZGtS3kOG/9GpYZeJoZVhLUpGQpVcOtLGcyVcnAYea80QQySJ
WzYFF7BtEyJZICBC2mQ6PR8tXU7w/YKqiVhFbdu1vgnkSiBfsW4Ug0DrJJr0LdQtMsUd4GEMeahp
SenYhvEajt2o4+G8BRdXn1qL6T3gDHvGZiFlnt6W7gNyWCnLhHyjvSevO1EOlfXqjkMNSRyyXSKQ
eU8SQlDB4VCZPppTiTWHLYVxKUzS2De90LLo1ND4o7Z/ADmEYgTjLLtnCRWd0j2zfxZ1h/vFClC9
0NEoycxSmL90F1PqB6eXh4qFgPBwyZBysizsBbrhZovZePcXBOMnVpTNsqM7ZUPuGyWKv7mYsUSU
8Kpp4VQlrCFS1xS1SHMW9z6k+0OQ6UzW2/yk+78VzrLmopMDFd8I3obYiTeLe07qkNIJ1f2b/enC
q7ChS/WnlEKAtss4zsQSdRRhuaJOJAW+xZEbfdxaS+4nw8Ln4gWsw0nlR62KghONYrCZcuMFNYuH
Yg3sHoXCY9bY7uaUnuNJlqV/eoh8mTpUQfYKAmkfneedYBDfw1+N7frj3DYkGyDAqW6u3lOzJJeN
bj9hlkVmM3Hg1Dv1vfc/lO6J4JN/EUflvObhqrf+X5VFOQTGsYojseOVITUvxDy9RqOad83yrxOu
YfH7mpvBI9iD4/mFuIhQXxwqZP8GokFCss28s3JUtoP3+lELyH1GTyX+rYOFNJVcJIPL4PkwoGkQ
tGU79oeuXrTJEZYXpQCff6XsuJqZuy6PA5ZiJMryhlb9R46wpNm6v/nAHOxUiXJaBlXgjHb0Q4Y0
83P10FrR+Se79UkWo/s6JBMXYy42eOEQb8nlvZY+oKDiesyeq6qfr4SjF7YBkLVmF8m3bcz7lrqq
KnTY3dLUfV5LJUyg+GyOqg7RNQ+QN7ni3fKE4ZhnfZtrYmoowEIHJG+v7jXJ3UrLk31vh+5JMU33
j32GLKKXVvH3sInAXddvHqs9oyI75P08ceguuLWhSnKoBpb6tqHhYwIYwxog3VvRgwnLO66KrDj+
wR8hmTAn5wQNjgB1+SRPZmQC8U0sciJGIddoerl7LGxLLd4hHimbNAzKEy+dZZV0HhxYfWS4hAOy
NxJkQYKQOXoO4vla9svofry0p21bBNlQjppsf+FVH4cJmdf3jkwhnBrgrnGzQ8pYp/EAfXDB0PmS
6+z11OjwOXNjlFKVaBU8hh7WyALpjHpL7FK3d5uv0JRfmHla1kqfqwVQI5WYZNaqBqkwJ0c2+8rz
HVtNGYZdruxaj0KJu39XAPLe+YUPCIl9tET2P7KPHtnIN0P6UB0VVKCDDj3xMeEBE2sR7tmj9BDL
5NDjXAVy4/Ab2eAQu4dURERd/3qFVLm/NTBH5MYiUEEs4TiBaUrtEjvf83d+L8oMjoUL5mKPIWox
uTPBHthVmKYyQdEP/SiNl1esC6urpxADtN9VS3oyJkIVR+LIjMZ01wxDE+JsHFsRxLtZSJEOVHkf
12Ld5P+bkBQRJitEV2cA797pfCcxjA61vbw9UxiWhc6+YvIlL9x8aZGYkgDD8Hb1gRRYMcGLAupz
0jgwLCvQfJcpUPzj1cZD19JepsDU9/GTTIraLbmnL98ZMJ3y5YFjNi/INc25VaxjRm9h3niB8NKh
HdqUxtSs269WqA1tZiBL39n0tRBC8JMlEU1hUSAP5sd97W+i1LQ+6Kbs4zUgwKq4sstbrstMDhJN
kPts3PrMRzIGp5QrNWUQqWCdFw2/yOpnCODAXgkklPQ0p1zZ5zRlMqZObkepqGdLiXfRltpgL+8e
PP1Kwc/X8YY5wJmDDhGKv71pRdNGWolxgPh8+98cHeciUiSeonyZb9jspU31LUDTnZDpY410nZ+x
DdXr4boJ1oaOh0xlhPseJZ29qyZ3hMF35R2r+CoyDkMEQVERb5fxyyZ75ssoNkazT4HhtMrL2fGJ
6hEz7ZAtZEFdbFq9rP7EO4uUCfRU9nwNbIDcU7kXK6fB8sXJjIWseMYOfvap/lsZo4hvgEuE923f
FltxXe+rDMXsqqkVzFQhRvUQi1b0rwuuR4yC9kEdsgFS3O0mPuO51egG66CM+Jo//X0Usyd87UqR
JRGgzKy6tZifPh81JKe0AprNlXtXSOzehN41IP4sHwwtkrReZOFXQtW7NFWn4gOhvHl5fdJ02CrJ
Kz/5X++9dmPwEThUBVW3tPlVq6/d5PT7TxiRoM7NaQWDTa7Vvddq8P/tu0V4/Y3DMNv9XdwszGzX
Z1IAcy6aeraAkDdxuMMtRVECEV/yowU3jCL/5V9nvAvt/MWD/sDh2P5fPU/iaCKKKSf/WCknClNf
f5F2uO6IBHYkpJEaWdWjzKzPTq7Qa4iX2CVqvqZkUMIV1wkMQI9+2hqNeRJqnF7ZXKn1ws/vf/q7
6GW0yyoYWlTiPCfk8RpcDtzztvVmmMLheiptmdmAa/l0jmRY3CMaCbogwqPqh3egzgkKozUo4yIJ
ML+ZT8LQX92L8KnUXlZrUWYw55zRk+bCzuNVgZRGZ5r/66JJlY3/JoVsYw00RLczztA5l7Kw4SIt
+BhNU9GoaIJTY9MDGhrjkaT5J4w1ZARgYfbnkwN9dbUuQr3Ana6o+FxIzoH44e9LHtFqcvA/yf+S
DdeLhsoCtwL0gmEC3zIOaFzx0hAmoFXC2qsLmrd/7a+woW14XQQ6oHL4SLtBVVjpuVnLQOh53lRl
+zCAGe/SOigW8K/epVUFHdMmm3GT8KnZyQOAlI6wdmI6eqBh2xDDLYAaQBhA3K0sulkyP6Dzmy7Z
5CeodByT/YB4F+MAwvSC4HfxnCPXlYGe9Ewb2P/iApg1FoQdwUHeRGx6/i7SdbtNP81Od769cDy1
yuAyX8d8NjQZgemsRKrL8aK7Xv9U9z0mXvJZ108eQ9ePcYaOBzuYpbezsddy0LkNN6HGPKra/Hhz
jYEkjo5s/cv3GA8Mrw5QEUFw2tnW0AtQfZPSw0kQlMTCd3ODWaSde8gUgyqPISK3o4q1TfR0nLae
iPGZ/uOg/2WhzLFb0wrxIYK1tlWRt89zvcQrZ8Wwg7eSqgChAeIjYu8SDRCNgkuUcuKm7cHnyiHW
WEBHVInOie4C1mxDdG6RNPMMmkNvZrmc2SBJqiNj0Sj5xzI4qUEhalVCvySE7jWBaY408qu+rs7n
x+d6C4lBVmNacACzu3aZV4zkimYcwKzdD2XXmdTxqqPXFTtWEsgyK8NyExcG9yq59x5mzhSdlv87
v67nTKaaioTaczEPB7EJ6SbsLSP/v+f19GCw7iMr+WR/FZ1U2brL3gJiWTAwpqgYuVnQGO2e4rVO
w74QR0qY0xLlOphfQAirYuJG+b4sX51YfkpATQaM+f3+3hqgLjIKybLwMyg4C18ghyYfKJquFadZ
zQy4WEwsTiaKwdz8zSkcIJRZtMmH7SsTriE0HViBqJdt1/BeS7vV8Rp39dvAtnIJ3lC+imiB1dsv
FiH1nu2/shI4a70kNxXf3jm3rQtITHx3wXFkD1oFobHtDfuo43xNC17sL0O7S8hLmJjpC552wdS6
DWGe3fGpcQNMr3fX3/CEWGJ9CpZkIjoXZWUd0KGz6FHk1ngxYdiYhf9OJgVwG7g2MqC5U+ca0DsF
SH9VB5hutzEd7Ymrs0khm4/l+SUL+179zenq8TdCZmaizvp3b268OSHs6TsYsBJTvWCdtENzG/7k
+6GAxk03OwumYqJ+EkVBNnsDNH81nGENApSqVQ7yn74SqzOvQUhvjw5NM0QNvKwMPjJ8dFrgI6HT
ZWlOUwkoZ0Vw/pLl9WI8ZK8e8xm3PatkW67eUtsPqZKEerbi+fwB+D7oHXrUM43NJ8AWNYH0Hnpy
m4Us/6g/Q+0KHbNDSV93sT4U4ipJxUN/ZXaGte5Q/7xsOAjqm0LIAk4x3vgwbd/Jb4VwVOwLlY7K
uOzJFK9uuBLN1EI7jRQBzNV61s+0KoH1QTGT/GGZM95ZlKO9YF9HVnCkjDv5XofLvxuFOnvP0xOn
dJM2yAX/DQHo3bZcQdH06g6tYzQNdeUvn/k9S2sJeFX0GcaKeQHNQjfX1i4vbSMclKdf0ztPAatx
Y9U/YaB5yymioT7FJrXaK2sMFz+QeFoxRZuIYM1bPv9womTmVmH5knfD2Oe3TpJIYAjiC9fsMId1
SaPM3IKFf7e0ScQsJ2/nC6aO6BiNoFOUw3U8ce8L8O1jG/XGymtjR3PHMlZkYwmLtR4nfVMH+mWG
yaykrlm9LDZWjAukF5L96wBpDPt02wLXKX68e+tsvez8TtIyC/fll+hmzRyEkvA8QXUPVg8ZA7n/
8CXp1D9oGJ3Pg1aeHCPqWix5FurWtrwirMQBQHYe9YtEHR7fvfpHoVrZCE4FFc4njom7DAPcEjvs
tVSqLrgng2cUhRnHfN6SeH3sTgZwVifUfQl5dizBc/6q9qi0/Lsrb/Z+r65jC6Jq9XTCtnaBD99l
9sezFD+ZzzeAhnS1T1t3MH+dQaXnE4LKJtMh3Sco9QniMFiuOZ2UUN+PlllCMI2FX61Lfelj/l4i
0I4pVEbJibg1wLs3ukbaNzMtxREmYL0a8VvNYhBpEUEgA/OHj0UgrlHc6N6EQeqEMmrGxkptCgTZ
MJDTeHdnMuOEEM27mHV8t7hYHXuvq68fBWGtStTb6UJpJzuMHy8yZdeFPG1Zm4OkXQKk+kfdUtvJ
1sKtMnLdJErc/rzjsmlGhlVrN8531UNBtOYjS4b+b2PUmnrURp7nES8YAhgLVxZJbNr0HYXyUGOy
kZYJphzJb1vGoXa1GurWJK1Z4B1ChZJgfedCB7DFXq70hpYzHVjKQ1uRBzAw/hYAayx2LCVv38Vx
Kshu93GaoQC7sOShrnJFOyzgUjfP/OAmzgwh/N8Bb3S8TUxl0JkHKLoPBdNs2bz/tPjAeAzFfDVl
wNteuMZASlPmnUJDH1B7f8CbJ7fTyjcZRd4mf2gtm67F4kBPNc6ooH7EkV2r+yPo/jl/K8vyYHaD
w9km3p/jMulhn4UTchFetZHPAjvcufwJ4819TqpN0XlqEkbTL74J8lkcOrcSR/nAme19+1f4mhm9
viq9D9+RSLaHOFw34jV/6LyAvM7KyOrqbr4jPZqzJ+6EUYRwuL5C/0AANQ//c3jYrF3bm0NN21XN
uJYQ+tRT59fIpoOplD7EbYsi8u6ZVLtULAGq9ItPCoqgqzHrWq8cwT5PcvNu3D853PqZGrAFV3nj
FaYptYa/KGps2DInyruiITJP+sZ1JEZAyMJIySt8hFWuhT8wj7FYdanQBvyltgifvsZXOfuYZxNq
/IrS0QoXZsTUOqMbZBMmfIRpNYFimXZhWiTOwj7woaqzoUuzKMZpb9QaBLjiR+NbICpwjwOwVHWq
3P4be0PEUOJAjXnhYgW03Fxn6epgW8LvH6CUEWNebrB0Ca612fiWCJi9wpJ8uQrb4hE4Ez1yE4ow
33ttlz5NOztI8HWR3GaYqhUe6pkz+3z+e/zVlFgKKx5mAz9IwNfyCCwSYuVH817AheIR01ZVu5wW
BHnMUHaxrogBlh24QuHA+N2bFxMHo4+iqe8IZJfwG/5iHBHZzyCR21DNyUR3EvOL9v+lpBBii+y8
zvec+MSoEqFHvMG/D0Ae4vcEr9V9P8UVFM14B/ZdDE2OA+kDDwUep5DoDlabjUGVfzr+akyggZTT
NIEAgVFgUvYd3Pq7xanm58EgOjW2mEXF+Z5XxbQqOQzal5+uBlfw40MfHaI5akvbDS4vO1JQAgX4
5w8kxEZF/o0sU9ME10amMxczRVgmvFXa7htigzYlrjGBAQ3gWr4QhNe5Wsiy0c5+ExuwyM30DJgf
gtJi2fwepiizu5qWsUQfRTzmTFXscmpMYEVbCuGh7AcWX7el3IY6zTZgrSuJo3QkUbVageQrHB5E
VUc5r8B3NOoVG7eXt0lWIWXRbRfqRWthIp6BT/kGKtr8fyGGzZ9kBHSd9EZTGZWLUYnLn3cgMZMc
oJIQCQGw6wJPZnPxpF/1L7b+JD/hAW9+2TngAERVoF6XNICUGMSjbJpA+96tkLkolVQYjNhH6VUu
e/70aug3vfA3p8CVFAyL1AlIpM0FSCLiGfob+j1KqKvR3HG5UQ+Ex22bacQjVaJ02a79j5puXNLY
JnWJbh/rDg2GmQAXCLSjIWAZALTKPck0PKOpxFhrWlHBw6EUna12LEKT0d0krL9LSHx/JUWR4Yqi
44oEe7F14++47wIhbgS3zqHjpQxD7K1p3VP5iWWIQmLPIJbT2YZgkHR8GiB7GDEgGRixEm8qFtXm
aUDGq6gtV0BTiwA/sbUo6NZUPHKcGd7udB1jvZcoXH/HxsydRq04SZl7EksU6r1011hib2wGYJ80
HuV3faXN6EWuvtRAB2/+GtU5THN7hkFoRIEPANl/qWioPmMDTmH+2x/dkUvzB9vZMpPql50mTvKC
gTVXxwxwr8ooNq6bwy2r+7eC300Qp+NoxWmykOCB3GbY484md7CTQyad42mhMchSRawzx0XAq2Qx
O5v3G/k4P1zSiEUnn/mHemccj48eP9kfWrHI5ySN2EQWmDy1pqlQ6cz23tTmj1FxK5A3vbDw5M6z
uVRFIYLaBsD8CCPyZDFm37F7zrlVl6XEZUf91AHrzRGzQfQt94kiGNGp6An9Bo7szolQLbeTonHa
LVBph2yYV+htG+oEqEVwQL6dghmd9jOqlq6gOsQ4Q+NmHbtVGt8s6a6oGYGX1BoKhxowTx5Bsz6b
jNYRALs28zo0AuiWERIno2aMGwqNRC9prsuka/L19uz7g2lGhs85U/+VgYa+FsUVNSyLhVoFyrLq
cleROujP8OWFtTcUcFbPKMars+MVGEcZY1xSUnKN55v5zACE1EtJYxoyvAPPSBU5ZzARE2qx/2sB
WKw1WG9qysO7T2n4BrCTS4/fxaWIvNGEj6F8Barb2vWpgrkRS6Vd6kXcead3ykxYEE5npCaaKyOA
pteObd2C3WsZzD2+14MqH7S+O/WKP0eR+uwWB9U1QvaBy/QBwLpxry8IkC6M7fhm2539HTfEaIeM
73+5uHCBs0Nrk9GHD644OAisrGLMd3QIeqsq3FmELFj5etSTDeBvEXdNCt6mWDnHn26wIlC1QALN
9uU5nrVS00mk/6fIuUnnpRT4y4sAiemvdwn95DN+ypXd03C0x3BRQMQ4vtw/+m1oVHVLjTq0z3Hz
GXhBMKWeY8Aq+AZLxRe7gk815UT0Gktz7JzB4zeOyyIcnHbG71/lvHq9Yk2Wm7fgWSWRaZZv7lIz
QgLtkKc8S9UlYazoQ2EBSAiJF/+zhaLE5cuw1Ic3XwERRxpNwGKMQvkYpI0FXyGlPWvHi0KuCyQa
nJo4ScxDz8Rs89lw/6rgkzp7TLnfxP51RbH8lGYShFc+TcRVsG8hSrmFBDbX4ogk5GDkFHY+N7Gj
bY+BifeWC4fUDow9kF9x5+/EnKdfFZpxyIc0yaGMyyR4Wzv76dKWv8tsjLuOERqUL0kyIiCYzYxK
hz+nxkWHEThccNTLDfbFFtPurd7U5lTSzGByBT4NCkU2rRVp5LrgajSvIPEW/4Hm6sEeNcdGk14Y
tfit3cIkZvlo371ljKEBaiBOAV8o5PvmikPMpMkc0FjzIpBuUfAlYc/KJhFgr1+fzMjhqruFxaXt
/6i0R3RYu/CDdpBDcsRKFgFbz1r33ijqCx9aiLqPOiqUL/jV48Y8n9YqE3CqJl/iuOGBeowQGyo5
ZxJSQiUqrE6HwLab+2TYZnbRjaFrZnRxl31zn2R6WCwrzB/E1qF5MJY7+/C62V4V4xJe9At7tRd4
vXAHFfDDQ7Jrsjf217oXKtwHTKHGG1uJ1o8cElK06j9+H+q0d2ZC/VKP9wepKOBDEwcZJJMWj99B
oLhMTKLT4ZYCouQ/FAYlhhEVzTLY86NKtAbfuZS8+TzdxJn3rnRHfgQhRgo5Tiyw7yNWew0GlC7Q
YjnN+clXhHOkIZ9Ictg7VYJXbOM8/1uonlrUa2K7bg3BWYtbniyRmRTzgNrWdvW6zuKNTVPdpFvF
nT0mGr1im0NxeyKfQqRR0hnSKbAKYqa8/uy7AgukIuAhpKtCNXqNyI/057CjO0ixCeWmWMWkTztV
O5y6QEOGxevFxbmMmFaSPtNnsuo1Zm70ndh4YcMpyqnq79nVlcVfl50HOUbpnmB0gnQedfG/3otd
TJnbD3s7T77vfhEs/Eem4mEkYSweW7lS9dCWyCjvTI17JUxG5AFR41qXLLq4TqM6YbLnjg3ng62f
DonF7lcpMXTPKQ58Tjxhvq3MewTMHVX0Zd+qarjoAHTeR6or1twK6n/cNww2yhJkrjbkUy0nUvRj
tscVg30quxVgo347CYJQYDPmMpDGPXKTJgGyDXMfk9oJEhbLzIeEhWPYslZjkLflun/4Mf44UOrh
4UgC5BIpb8/08PcPspcK3/oXoXH7/bE9NHN7b96CqtjW4Du4alsqYBsK/70wAH8qmT40Ye4Qd6Cs
kHHgJ1F+vdiamG4eRUjI1NC7/moKWft/6ASR3HfTk2z010/Qpn++jZFqVZca6j9yen3W0/5t9wPq
Xh119oduv3vkY32LzQ6ka/81Lrs7GeGa5QzvJVnhHPz9bBjLbi8VolE7duCQyqrlZp42u3t/Fxgx
Oconm1e8ci00ELWNhGDQ1F4U/G+7XuFOEhfakE160/DjONCnHkagly/Fb2QGiziS7pIdvQ+cspUZ
eA+N+G/bnrowHb2NLc30cfiRsuuSpDu7zNfPdHOQ2etz4hLFd2jsxtKuXXbpfgvpLCjTKQ+qJijS
D5K72Ay8m02GXnvs3CEK3YaezB/b64vTrL5FYImFXybvx08hxg1DU6jRaermskDWhWkPtZrns7kQ
O/EgQXzcB7oNpe0zwSPi4VAdZcwdVMlSAapgG5DgbRyyFeMP5gZyU+mSm1Mi/cSgl6dhqTLTeMAV
JvihGvro8FS+RJdRN/ZgnuSSGWxYAyk7Su2iLSE5hbYGwndJ6sDUzhCO6WA2wLKl22FNEkdclyC+
6YAlE7VHoT8v41Bzwbb9dro//6H+N/wcqydpEHdvqUga3DVKrurtP6Ls8KgTqKh0jObcXqAKmzBT
1j519nwL9WHkQRzcZrK2DkcbPZVSOW9Q5iq5ing8nNiWRZS9wZbUmNwzLEUb/z3rGUaawVSvsOln
e0nMg72GsKWQWp6nmOqU5JwdYyAr7taFtd2vGxLqWqKCbJxuxaeC8b2bPtuY/ccYqeuAUIeHBg2Q
coMcQjxmoRj1/RVFC9NqqKbroKVjWRbgIBhU6D8kKIvweosQPnlB5OxmBP3ZXOF9ickJL9ntLjo2
J4TrW2i8IDpefx2DH8Kn4SsAKt1E6RzqlQp1hYk4bYIfZh5wm7pyv47Q1Riwjryi8xaGoqJEsGIM
4J0t/y3l9+Ji5dq8vhE/uw+faBY0HqiWSb4n8bow3cV4Rbfx6VNFyMk9DzuKSnqVg84S6vupTnAR
ZkbdgxutIHYKzFBmOr1rYVXickwbYlmHQtsLMHCoxvmPT1Di3QSlscFxWdddQrrnoyfK1COjgeRD
UMaRJPRm11vzL7JKElyzbtwEvK0L3LRk3l9ePs/ffqLFqwj2O82uwL51CsHI291iQG3PdYyEQtOV
XGlrv01TBMz6dX5BY+JH2BzxxREJJ5p6oppV0D+85ODJF3Yj9FhQqtBVnVMZXCB/wFXCygsfPhVQ
1FJaMJO9YleucEkCSiHd09kkT56KFBvNpgrZaWQvD+JOt0BeOrgqdjQpk8D3f334DoO+ZjtLGuCK
OnXIzUZ/9TQCx0+hgTDH16WjVO7lQ04rA4uMtS9d6GAG5K7u7RpkpuSgWykuggT4yDF9QcS4HptR
ArCrcLc8fC/rskzJ/1MIw3zSpQXjYo1Nt/EDKg/LnZMg8jweFyln1clUL5XbHJPdApMcs+YaIe1M
OWW1s3x95sR2FQBoSS6vU/E+ZlrjvxCDt7SufJhYcG9uBfyES+wg5vNJj72yu4HyoWcIrEpNRZYH
NE6+40KNYTGl0JRN8eX0dDuyg0QfbOgxdtEhfSB2mz2DmyQkZdxodyA22jbUN2sihZOcDv8KU+9+
3fWhh0HJ+2lOO4eV/TTjMwfDMAOk/0IyDjn0s+gpKH5e7Uqq5DtKTcwBtbs+sgwIu51je7wXTcZp
iIQvXW/Cvlej0hgrP2UmO/p7gcRblsB+SptThsOMaw5XFPom3uR72wjgCbJAPLSiKxWGcAxcJvYw
XGxsJzaUtYptZjjQanbmX9LPMofuAjR/bSMmdWM8vNYYlkP1R723oQOYjhy93t7A0d0LM45PpJKC
JhiRCspFsShcNS6k3gE5DFSexsndvs/R7qvCjf8n75ihw9FDnl66RCNUjLtgzqsGGuhnhBx1v/AC
KiOo5lMDad2kTpR3aEvvZkSIbvj9XrPJ5xY6hjoJ5mCkTtF3OFrqJU4vWMqVZmMw84QizoKczCie
g+b+g356YmV+r8VRyTg7Pb9AZbT5lADGNIDkXqhSU4RYYtKspAA1IvMljEk/t8dSF+kM7V6nw49n
fvx1lQQftMYfu88i8Fy/PimyB2SFFMcrrwZLM4/hZWzfovvjc5OMyP/PbEPJtmXWZx5uYz4mVP7z
/Y3Wjp4RCtMfnfqefjaDJxbgs2GSP3atbO3ImeBCxXD00UV1SKNXz3W2clDerZlSWpVodnl0NyR4
MuLSZmbsvz9xcVmOZhSPG7jIB5HVEHhAQLp4IAm32IzoeVsTaYMIBr2Vp4gBJ54dV26QCnZhjOpX
pYMWmpPpRY5m89T/peRc688rndmD5tSLUoKQAGywB3pFAjwMYLCyuLklUlofIM3ZhnqAtX2H2BLF
QS29vlAwJJfyW9XT7g6hZ3J1GCbmELU794eQYh4tsrW8Uo5b5/EJB36EzVkHcFJiY5J4+1L3Nag2
pMY0WL/Cccjm1mDNVTu9iU7klTOqDXZhOqHsGvsIIhkogav4ccun6nCmezSQw+k5pHI3PRggHDAw
apCHnzEzJAs6VtsqMtlRdndLLS2wu23gxLYcP6j13kTYTskPUcYIsvy+8muoT9zTcBsq2UPXXALO
zczRyMBUM55yFhl6pKwXITaDOJL75qbQ/o1EiqycayxkVjzTB3I6uAN0rLlbNwnPd1CAAOXQU+ct
A/EIuDOJvTfMu7EWRQflUAI8JPr30sCHnaJF34+hYwLU/Ow4WJgO+MFMlckCM8hMhtDE0fqtp78c
m4SoRobktH/z0FrkZKPiKcpIJQ28RHppJaLf5nUlnx13caqu8ZCS9IR8t5jjyKkKH10nTeUWpyvN
EOLej7d42UVOWB2oF8TDjYPJyre2qRXq3NgjTsm71eClWTmAetxXz1Clt5Xcij0KS2HK5ARdNBIb
zgDxPzSkZ9MzljkWwlW18u4Da0bk6tlZ5VFjPAPEIIvqCEJa5x8PN1xgy+CsIBNUccYWkg7bD9kb
0sqLzmmoCeMMddm97jvJpiQ39QP6Te2i0qRzGSo8TUz1ZhSBZpyutVKUaORu27MLZWYMoixw94X8
DeojazgISPfQVaR+4F8VB7h8ZqmM7RxDMwvXbBWfB3Ecs6lZq+qcx2MJEtcbZsYLmhQVHneDRERq
5w4ieVndHgZfmR///78zmNnZ7DOxSYDsp0NMiyH8rtQb+tvfl5ziuTVPX0lSI3det9ACQGUrcIXN
n+4YvR2xRZ8a2TevQi4/dRuxZxjrwBcN++z1mKjw7K2jQOmDhvbFFbNFpgh2wgWuBy9tDxlwypfN
clcPecPtrx+j759ZNXXMTAd+fwHtmtE6HMdsOTJ/BI3u/sCo0DDAR8rJyLqE9lTwouPA0QK3z3iC
GdpErmbM96UzHkErSmxdpD1n+lp+vdL2OU+aUJ7rkncwd+XuUVNPwmoXolqyPmWio/q+tlopDYbb
cEJe6MrMa//wcNU0tq23C44oh5V+DbRC4Z1Ni7mfV2v6b9iPKpKvZgN8AH89lbqgD22jGwLe29qU
tQ35dPAOhULVGPYYNGwSn8r88t266q9y9KggPpk+SlysUrtC6AyKsCKMcuumWETPOSC/hbYxJBKT
jwUzlpl1qYwX9KNTx06H7291Z/MUGC9LDn1w0k+ZmgySn2ZkfBKmmq0lLVXggE+bveYFjIhoi45I
plODnCjqNPQzVaQMO5fUgN3SNo3xbvwdQkBsfx+oO1NzLfP3ucRnbpFe90IC5K3i9cjbVsJizO/H
yLutFp14id+0PQl/E5ZnaBB8sI0IniwdZIPO2XpLQ4x1OcWHQdMQF8fdNI4keP7YNj3dKZco3JEY
VnoVQopM12Gm+DsDlVGtgkl7LyA8tE1v0APq6M6oK5zNeWLqChcu1cFtUvq1qXyJJ72ozZTHjXUm
Bh+TW/HoMhevufIqE1d9pmqbnYFpH3zObjqaboLExMZoDMz/YtoAefkhTG0JEyvA2qtXNUCN34Vo
WwASZroh3+08IIhlp3hRonJEoHZqi0Tl/7cK3d2UhiCdiztj2eg5xYP1Ua0wjLR6tjHGY+HpNqBu
rtJXyASNVZL5BAeFRfYVPsxNINNaKHAioceP7xHMsOU0tm7LYIh3z0OVilc6yza/Jv+07NszVB/Y
/fHOXOwgiuhZ035ldTF15p/pdjUAnWX2aY6bwjHHnB4nIc19whcImB1f4gd6PUgMdRSbDaVGx6xF
W6xSbqkJICueVFraES78DNjeIj+67GRHiVESIujCwFb6Wde2OUljhq67VF9UDsdYg5iedspcvI6C
hHurcdTcKqmY+O5/tsaueteRhtRo21j8GPH9vVBsvkTlY/XFx1JagwXA8R2HLsEj8YP5hmrTr73P
95DWWRF+jvvzNV+SP0twwFaGYAaS0PuXKhMueeKucP7bwCsvQqXMIYEUD4s1R9Fmn86NLKQ3lrM3
ps4cl4cp+gA+7YDgpRBzHLIcqhzzubTItIC13aSQzhGSOqa3O4EYLb7H0+p8/Qji5AGGFULPWPyU
J4AJ7YDNd45NSuSLVYFnRlDgz/bdOZ9KijyUntzEh9LufIJS39baiGMrGnl7HBTAgU1TcR46BN4N
xdcK5g1LXJf2+nWXz4mDyYdfkSBq4cRJlA5jrZhHKn/ZP6IP0uIrch0u7gI9Lk20IwbAeYEgTmUY
xg/iC/ayQxkr6lLtoBDQY8A9HPjw331Ywkkqn5k7Ly7sv57OwdRY3N0b62PvRnMAu19cTaptvSI6
sMtPp/gFPg18tdvPxuiyp68jJ9Q2dagWU5zsoIw41YGYI6KnJFRwXcsupB0FKcszMn7HGmzaExTT
5xiSVmCdwazNnLgEyxowihHA+Plq2qRfrhrHeSW8Ezfv5hH4+tgetgGv+lktSt6mf5FZpsy90XgP
t5VorYESncTmgaOTMfoATTIccsfTo4yg7R839iPSWB2hbTmfKwqTVT7ZxQ2oSe9nYDYkL6Cm409R
gVk/x8Ix8woGiO7eyt1JAoxtQrIntBcnm1KTSaTGUiyyrwUQpkjp1A6yGjPGLbdZBCy8nEye2Wl4
7OLZirJUegoaE8CvLmVuhQQV5KRH7Tz0Z6cY3S+vR0Q6W6CitXtbOFAXHQDu3rbnZkmcTVMDhGM9
OMLI7RpQN01YqJLjEkd60+eujMI0F+DOzW9Qk4wEhA0uZuVe8y0MZoO48ZdP2qO7+iqqYPV/QhzR
0m90cXdV4OtO5etkriaAfmnip1U1nkHMLrLUt7LP0uMNo4OWuYd9s6zY+VoV1V4B5Umm2SOY0Smz
GbW8/D26O1M9UvT3j1UhJ02CKO/x2IUoKy7GxRV5nBT5vz9xAzQkD36nqQu4VZtoS5O8fOEWmyIF
UMNoDN/0zvjsOxFEsnTbiJ4PO6qim4YIFbBRhPPJoOWDuNUmDmRs7GwxMS5s+dcWFYMs3nJCZm3N
3WgdY1VhTb/SlDLFL9nosqXA6KX7HUcx+nscAaWlauIA+ti2KLQ85UKaNSIpEehwIZ/z1tWmcyeE
iHsvNUD4yFbkMgRWLstaobpYs7JaVRWKdhTnNVYinWxZUJScB1c45GVZIL4n6RbtX9J3SBtdkdG0
gPh/XtTUXOvsc51pFXvNACUMdNoSNxjRjPnjr3In9Pn+jCzLijISrKP9kijcaWpKdBgi9pfGnMSM
EhSC6YLRNS6n/HQ/bss0zmx/SpucZGrNH2aLbG4ey9+aDW5h1FXSmk53ABx7JvmaDVfV2ek4DxeG
np38DRTJBLS1/GmA7sgMXqOx8E/4ekJKk6ek1Z3fZ7ifkCBzAbdHGzt8nNSqnqUunRjLL2VcEePh
wW4HxGuIGE9601/io4qW73fzMZWcTMm7ScM/Jho0FmSH0v8sRvy08wmPl829lLB7IF3yRxoLbBgZ
GM0jR5rJIhxiIJZnLMJDvi4Znkqqms4uO/TQWninMpZF3eSdu583sun2VzqxniiBueRda9Y2ad+Q
GHnY2af2lTVGMVSnC7u7atwC+L7Odk8g9PEpjj7wg8qxf6ERD5y4sEFRMYJruHtkNopAQy/CyXbF
q7tPwlnx1lPGNDBEFP72Tt8yzHzqykBUS4h8Tpe/0VLpm9qdvEG8PBDLa21li0RPSD4246mxumoW
8x1wUwvdW/DFeEErq+0Kay3VbvR0ab7lTP+D1qrSDaO92FdyNoUEY9eJmUBHMlzFfOX63o8TdiPD
qNHoITe6atdlelUqmcul/lnCVcGVVn+ULe+u46uVdo8E9rYW6lXytwVK9AsdtcZ1gtiq28zz1LRD
NvZnbZlt5lGgFcFEjXZmq2ndOudGzX/aE6l1WPvr4Mjvv4tHdDcblsMjI7RJTU8nmH2ZyBNY1Zum
ik+OAQLDWs3YG0Cc6YGIWTY2VfzdnN0WNBgesDWv/jct5dxUTY+mfU+uqYQ3Jgajqph6cjxHyPxR
Vx/zQLkRmn6ojPHqkJtWr0UfxuO3o4mb3/3WNqtB/S0FHs+9HiRnpshWUR7mJmRHlj0kYgfrLvNm
SD5xqgQWnnI2KMU6bnUQKjgQMQqG8HLhT52ThTLwwBJi80+JkzwqAwB4ZhPr02Wr/E9AReLTbp3Y
raCT3HZM3lhbz9EoKk83oRIVWLEIEd6EtR0IvxRj04tTwh6+R1Y+oAzxY5heS3sZ2jMkCAm0kAPu
HMee7hJgpJfasmC5E+jymZvNzJ0zBKoT+Wdw1PA6jTS5eWVQM/LcYG5GUJI9a6/mqdCPUGofepUT
ZaEQ9kijkVBPDxLCv9HwkYK66XLi6TWCdPENEOFMIlwZSCrPnnHgdXAJ6dJe4AyuYX/JYnPbZjw8
zJbilcR7/NXGZH2MjHIhWoBcnHTye59333K059H2t6D8Md1iYt87RWAFbGt39rkDa4Yisxxa6lO7
IRT15RJSyC1We8VajJ87YrL+w0K4I13Q2XnEG41QAiw2Gl4lclAnqPJJO92a4HVaM0/NtxbiV7WA
+mZwu5lw18/P7Q30/sy0kFIys3pMtj7Fr5F4IM97spriqxC+x9tPPdtFNNTllOnXESVnExbL2S96
bpuaHWOy64hTVxlbZIuuYQeLY+g13FhqGAzYjT+RX5m1Mbw1uohfrT6aoTJAjpjyW/6lZWznpKM9
/4/15kZrDz5cGzlGwDXJ6FKUCv6XjiiIYb2Svy09PEoGWcEvc3+oikHcFtpSkJq48lOHvimv0OYT
lg6G7WEJG9ZbEWv9bLkT25kjfCuMKK504w6MoYC/Lqi+NoxmJaqOmZ6DzwNKgB03IFk9f9kR5MFV
3enOzTUHl8p/pv4imLkwKKQrConnZxLxDvKoO5abpe4VocpVcuzBiJlWBBRF2injHf/3eceffMjQ
hzygRMXwt+s7Ja4MWcvR6n1Xtvopsqx+6RbPQkUbDzsi4ijvBd+uYfBlpIRvoPn8qeFNVvi4HJMj
okaxpu+U7JDmNKViVWA+nk6YGhiaOk9Sc6bdGc3jDdVHGkXvXbAvewO631cZDpofJl/SSUmYO4AL
jNM6B+RgBLfoGSIHlEruzBtQbtLgTk3qlHS2tMDedEg182flOC1YPYaBFz4OFvdc9H6kdIJ9lfBv
VRF/7qyVhlI3KKEvA9InljN/kRgZybjjm6N2+3pRvhUNL6JG07ROMjK/cL0V+HY+Z66E9qOJq7p8
6XgVs7RdA1x0dX0YOPgOubTegg96xKaOfU+uLSGpUq2DkoIKzn7GgzgWwF3YP5WqCq5H8VqZJpRL
cOC63Sib/eAhQeMeR+e5XrlkRsHPSYKCgdH0bFE/JxFnkdVlSKJEOoIjJw3asUPMHbn+sYMthiR8
Wia2w5kd1DlZcYzzEWuCMqIP3hIN56Up0pvpBnt/AAv7CQA8R5vHj5pEZziSoxg5KOY8gHn+UhFq
2Nw/u/e6kX3lYeQ5mI3a1mn733GVEaVuFL+WCpllzRT2bGogq2RzDY8786CgWdJ8WDKfUtgQyoxC
wGE47h8PEYA94/gypPyzL6T+VKvEUwdPnaInAuvMqBcbs5sqo1r2wcwRyBY/C6WCf2vM0U7vJM6p
hvMuo0ZV/WrRgSEv2wh/NlvkRoZTiyxZ4Zflfe4AH61Ti2/OsPdr9cb4C8x+OEUjvvGl74daIyk1
zXcBizJn4OR8ssij7M26R65nkNSf1v9le+0VUBjSb1iiYLVRclkFaKk7x9y+VOD06HkGxcPuWr5s
lJFEOPEI7KnGNjl6A+P0OUgYDNwO0PJS46jl+6LiXhHKJdU4cRTIH7kzGv+wQ7fqzMc2y+X3AKGq
Ptft4wFAwmZpMZH+jAJ542jgXSNbW2vWxiL3ITEtWKXOhuY6bOs2POw+PgkePapkK85Gplyew5eo
xUPCP7JqlaEPGrzF9NW/Kldas5BfXHNWhnXtu7NSEbBQECbKp4SN2ZlsSzx6lJRiaWi2+loyST/i
AqakienFKbsdMDpnRWJRmOoxePd/KxJeEDaLv2JSvP9AaHRyXRL+YcITu30xHKi5yc8a8lmg1cfa
rPsAD8WbFsxqYzl0pf35Z9QMfExMBCdhvsy8qkRm1ixOQf9BHzYa7NAxKry3eKUgzmYDi16zxsh3
OYyK9548WMEEkKhXVaDxsQ6fFkbvQcxoma0otIypDyUlJXBdLXddT9U6cJwuQZdtGJzJJXA79Zsz
1dU3m3nD38W+6rrrM8maQHAWWe/T2zS/LACd9BBnfqu9/HPzLqgQg2t7R1IZ5iy2ryrOBYjoSKt3
fZq/DZ3fNCt+kUKDQoCMrPSpDT5+jleI1QSYUvwppE/c+JtXbZs1A7Rxg2gd1f7ZDC6rqtUO9z/3
v9iDrCCANFVrO7vdEX+lz/pP8+kyrj61JXrOgmlMACAP6hs+iTbEHZP+fbdqtBHIk6UGKQCr4Pvp
YLjNUbM/vEGcNyvGPKRD2JoVou6FEsTDXv49x0ej5gJf4nCNv89fJf/YaKwhPUlz9cI79bZqADgz
JxLa74t3jMu354lEdd2kqLZyWKT7okmMfV7TOQCmaAhjfFG2zDFmp0Oiva/U4o63yYHMk/w6S1y8
P16Ijnw6tqQIY3Ii+AcsWJnAMpp3LTLtT6bt4DF8UZoCPRCRPWKHRFJLu1sFphdOdyYABmg/XnAT
vWCKyu2BtwWccxYizu0jX818lDme9R8Q8Ur3q9/qhByDke0wtdS17DFsZlNla53egvsGT1WBLLH2
kEt0NWzMivhmVZXuguJyTss2imi2qdEQ9xKh/Qf1hg7Na3a655h0ky5sedRaGB+65oFeY5IFv7ws
FXodMbnXiXS/k/nUDLeZYkgv3RKO+9DcyUSSOl416+RvNQ9qA/RM1P/x3cd1rdKbb92cK4ENg0Q7
d77kE9+rJFcbfH5Hs+hwFpCq09djtlo94Si2H5v1x3h1ckQHv+IfDAjJmIMGgokgq09XZr7EF/Yn
B4PmDxwfTbR4WNC16wCVg5b/5GrYi2HJ+JNdcDI38eKHToXSiNLJg1tT0qgXKzvkssyjQpNH9y2N
bW4Oyro/5kK3uIvGhPQ4PZXx7hUZqDHAORxRdgtqNMyc8YUm6RjCjJNrzxxqMAL04zQiNv7l+8HI
yaF0+6POt148pJZUsdkhqBGjkjGlqz7lLL8OZ9WGGWthDLsyiQTGOGuFPNzfdKZHBns5oz+/Mv09
776tUq6nT+mY0LnuAiM1Atl1319N9SWtBffwgf1QGD9F96FufueRCN7ZgJrwSFGiiR0X0n9AMbL1
ZIeYd8h3O5GDt3il/5Rd3Iu9wLQwm/THBbCjOReh2XSGjJkaPfijsnw/QwBMNBF5NqlmmhwZEtak
NIQvwXXxaXDH8bFsNxBJt6fyes7aoFoIUOVGZL+IBlzl9A2mteO53AVF5eNFfDeG/SZl804i5Ee1
W7MPpWBES/We2eRtj/BzWy7cPa1jXCMITarKabFnGcnytMnmWHdP6r9Tfp+Xhyc1nb9mG0ZKJb1w
5aAa3WDEzl40EUF6U5ng/LpjAX1EANXpxj5s2/0LFYLeZ3keJu9W/LcIuOACG/86tGZ9KuWP51Rm
sGOXFi3MMPpBFRylxL7XIcagVzT9Qjt/dNJz8t1PIVBs2tNbyBMZu9YZAhAwYkrA9L7odgMVTYYs
CiZP0z7EA2kXX8V/LK7ovHlhe+Dvg1rW0v+QzHM5lxAMpoiEdOvi0R7Snxfm8Y+giBYHKUjcefqi
3P3x69cschL+NeGRKs7AOrHyHKTceFFAIkKkWtOuQceSL4CTfm03FrCiUadRpZ6dt+quah6d5nSQ
m1l8pvQtU3eYwwgee/E5JU+9TBW1y/VuYUmKaCBUMOUjvCspkmfYqDmjUiuc/xuMU8NjLrirs2ue
nGyxTihMnose9Ek3kgvPQFKs2HNo2mTDyAjZtakw6KB4Yf1FeNLGrllHtRKANoAq0wq50J/tNVGu
6aBtaSvPe3JO8da3zajh+JrfYl67j57ufHiIOJrtk4AR6RBN8rqZmhvMAnnA7I6kSXRDnSI8Rzyp
KoKZ7SQ7jH2I7ymQcwrbYxzo8MEZ+OTS2e7aQLwQx9rPaORuGssOt0kQaZfya9SCJ5mB+WeXTpCx
/c3oNlx6PUw2CF3c2N/Od/wduldnaWko6l1kZJ96Q9uwy/8x5uJHhdmrt5QHGX/A4gOTjdF6alS8
TN4Is274mJdKCoLWQ818nFdfv+sQ5WdGyCREx3dYpYr6mTraS+csA22y3H7o58ZJ22cqbapJU4+O
+5tG2JcYgyd4nYJWfnFZz0Jx0Bzn/7REVmIe5CDWxeV9BxkyZnGViNigWmjUKoMpicVWRI2mJSBS
/g7s+tmEvAvJ/wafdlHHUDUcGqs/Rm6XoCgV0M3vdos5MfJRgRVvkjp8uL5abACdWdJvLH9gI+rU
Md/S7iAmEQPddAUm4PZokZ9g1wBkneYwaKDtUsMjhZiGb/AlmpcrEwDhpKc5xEqVQN88UCnIVI2N
9/L8oyNXssaIRnIKoN3jh4cnxYUpYRq8V6kGs6iTVn0QS5BB14Ivy2Oi9J+BULbt4tnmYE4dcYNq
rT9Qw78nrVxbruDyMIe2tMtuVrZqEjL/jidiBA0Va62p0uJUzSoFPBnsgHwcdOlmvFwh89hTZL3X
BAUwlgtCHMbOVPl14uAzXgPjABSVEqO0+WejO9jt+ldb8hDiUyTNAqVWVlRVgmmDqjsS0WQgFyvj
a5XzRnxAw+92K7yhbw9DFbVdnfU6MsbKVFWztaTR1rVzPjdGvaSNUxhGBx2TvugyuoGUJvlzYD9i
tiZ3Y4yqYYoe7tqrzVdojh0/RSYtYTHwqSA6pwsxsx1yZCakBy70QPpythz5cQvjcMeXxM6ByZNH
mC9/BC5Taz0nmenZ6nD8AsDpDBgFi3sF686TBJ+Zc87uniWOVrepC4KJ0h876SIw1OMdWxo+H68g
Xlj/bJMbax/Y0DDPVF4l9DA2pYTo0vONeRwfXKDb+XGdktBlfUb1KgMn7rSFKipm4oXfJrfszC4T
Cp2HUrXuAVW8BCX2OyBkB0+wROVOLueGIcJ1V7y3CaWe3S4WUR54FwExzzFWFJ1Q5uKlSIc38oDZ
Ei61ulzKLsVWb7+eClH0Jo/wLj+ZxJfBEo+d20tJFJ683IYUVuoXH+XF3WO1HRI+gLFruHDvTCJX
RmOVWpeQDu9eLmRiWC4oMXG2S+3tZHnhwAm3erxmsa+Ttk5OgKMqYDj3hE0mBSh3sxLi7TLbnEBM
Y5SSySXjSVBXWQTELQghlQG2Bg+p2hzLwis7rpkVNQh1ikaDfoxPBFYa6yuIDhHMwR0gKXjPPlpH
SqLnnvufVQQLean89CT+PTKpHk83CA3KJ8RQ5AjZYT8F59+523sc01GIRErj9peM/sOB3HWSpyRi
K52kMSfeHIUvNFR9XOyRVZEGIUXVVb7KPShb0C3T7nS9xIw7B+bAtCcFs2fA0GEjDR0V1GRtmXcb
NHGvkP2cWtfGYPlhGZs49fRUDrm1bn1xXVMAIFkXdURv9DKVrt03Xa0Fw09KG9DLgiPxiUFTog6E
NTGCJZim8wVTbU8VrM6X9xHNW+UkBPXBS++7YAsxbPak50sWJCBzECwjv4aQPwSzEQjitw1/InIx
O99dS9fGcpYSPAo1EOA/7eAOMxgCJMdo5h6kGdq1fBy5ufzpJ1n+USL11nhngW8sSellGb2zZRfo
ywcXKGuus8dT/wQYIKVT9qeN11MBmYw7CkUBUH9U4wKtvf2Pw8y/AAxnWxuU4WBK3Bh3GmB4aOEF
iSoVZ7cUhCWUgPQxVngIHTv9j00noCrcG4JhVmuWW+ImhQYa7bGGViSHa9M9MZ5cYHCOF7PJtO/9
WiglfgD3xiL5QeYFhzUmIB+nZYNGfjXcfaGS0VAkKURRNGCDCV1MB2Wat4++5PhymKSVR48Dq5Z9
WBUnD5/KPIXHokTfpRzKeo/gVt619mcSVgQdkYbz24djDeYNaECVtqfFfvf4xRGHQoZhwRIogtZ9
HvDBsyYWaxKPhF1gl83UyyMkAqKLMgGQ/XCWxmw1Ui1UJplshLbyUl6jvM66ZATb43Ti3LUG/Qpc
TUxufQ/ZjWSSBv4HFDPfju5ZZvwBFgZJcY7xIdxKxRLwgv59DSkvwvqu/cTyqvS03cl21FR/CXcb
vFURYrQdvV+2W/1EoCZ06sLmUTKzhtklLJnia2gRFxqn1rS0VjiUyn5eULwGSEFgrcrhFd+XjW9/
MFtQCTrk04iw0tWZJIs/6hJ7DG1y6X7MJnFB565BX2C2tIftRD1uVKlpasSIicg23AYmQTbdO6N/
BQCdCjuA29oQzVQZpO3L9sbk8Q63OaARgkcMlY1fERsi3CPkWbdw0N6ufuhKy8JKk8rUJ5cBW+DN
eeRWdNGSl5GIbS+av+SDj6qB4M0kd1/5L8jHJyv/qh6Q7CPH0x357wVWXh1CFE8lfrkTHhEGyMSQ
GAsKHywytIJ9I9TD0LwllhouCPTTAI6xek3DHIdHX4hv8ddNcUh6Tx7zFnsEHZUMAHbZijXRndTi
Cyz/CphKS05qJQIeiA01uPOTbmKXqmIV1wfGQ0smiMKWbF+HO+OGF2ENAdytf2/FMN2kNVz/4W0P
I8wBWYXGbRdwVhHr77SfPaeWqxzVgtiItrV8jbcp0GF7uXX2sMZuFJmlbD8ePH5hDOr7zfYYorKH
H3wKG+/an5eabdBUADt6XQV9cx6jqamgLf+4rbu/k2zrBSuURyxyCpUJ6I+SO+JhK8Oq+XM5zv34
CDRTL1yCGXorQkcGhvF8F52maQMHz9hJqXRfTgwEP16G32Oq1ELvR+6MVDWMW+uhlyRh6MvUWqgP
+5R7KRDZjuEYn+tyGQFdtVhSq1M+nsqNpx/geDEqyONh/vekPM/eTa1DfA5bL1inhK0raOKlQt/g
0/tnmBl7QAd12yyfawfycVdJvJ8Y2Yr1iVYkP8oE1m1COmuwO/PV2sIYE2deud4Y4Vp75UABxzSM
Y7uWT8idHW4rjc1sZ5EgJ06SRwkYYC4iDWr/VPWXJ2YCeJfJUz6qYMPA5IMLtEYvuf/Ec6aPYUVT
OBZ6B58dc8RyHGdVwGlxP1+QdxOBlIly10NPXY9/2Rk8WEbDTPxdI3GuT4lOShTen62WOOwvFQ3B
4v5q5tgK5ByfJIfBHzoVglvgDtj9DYQtB+fkj1f+u8BDPJuEuPr/FXvsTm42twApzaKrFD2xIXwi
VPJVqwOeFfxX/8hifmXMIva95xRDKnB8UJkmrgS6KnyWLSfNXu3/xkJa0j05GhXWYWyaYDHAKf91
sM1Buk8JuVhM9RfMNhy9IIS+z1dNAnntZtklV1RxsB6OBCpUxpvIfi+Tl67V9l2SgCq2d9OmUYkT
hi312Pc9qiTFwvOt7uqI0fRwdI+PAUNpdnjldO1Q9GaLNgkaxUyiaGdUXIaj57tgHSD3yNeRUJBz
YqS90eKBjEMPxd5pIGjcfPUKkQWLWnOldN/N3AWYgtBeFR8RHRxCJnOU4h+Ro8qO9nZmQAsG/XL2
P8AMsoBveRzj5Vv1YtSJjZJdcE90fUSXWYTOkFR2z3YZOQfY2f0Wv3ZGf33K6IzAv7jJPGPAu5B2
v2Bw0OaAZGZxRdiiJg9fQ5KTy9ieKg6z61Q/jh/XRLWiSqX3xY4ysBHYz1U+5zHROGbGqYkwqfrj
ech4lq3fe+nv8L2/UZx5x+s57HW1xijNHT986YcCGUPB0aUFii6o00S6HvMR3NIMVoGNf65W4R04
PI5GzUmOvNql2cZaCcm8CyDODV2gihuIrCnVWXH6pO4X9GmntGHj6+aIgsQtqnR2ZtlbcD7xFq5o
nFbQ79fUOIDHxCvAIJLTGrkRq60yM7jmwv7zMCFswn5mUVb2IcpPzBhAqy1zcleR0xwrfTzL4ynw
VEKFteDB2kbJlBSn5c6dnCZm5qARuZvI44PztORwG4leYZHxZt3aQIdHYg9OWbrGEJh0YPALc0Sb
r7JKYOfHEiRsaosVn2d+arOSpRkiEciAzwbK2bQoWBbg8pG41FKNpoguP0QRo+LVawxhzMZoXr79
sb4ZMUOWXIKrtyJs+TdpU9FgSMJ/K8V1pcLuybVPVBHvavYK4xTV6vxDOfCiLeHbSt2tNncN+Ows
VkxSZC2ttivmhEeBl9gaKW/yVFdYF39WSOBq5ET1kkV32VnMjOriPM3EXxWynfU7nvAF2q5+x6Ad
f+tuF63sfTydiFGR/7LD26od3IwfEsfxsMnvv1an7O4KLgSysKEuM9E/gOCcpY+nhBjJJ3FQk2dp
Jp+3H8/OWeEXVtaQ1jGnKPkwx2zk9N04/JOOo7bA2cK/jouLXh6PVA6JUdDul04nJRmUMa4IK+WX
bJu21TDsCucvvzWf/PBNVAc4UamEQdlgQKNP5MsyIcecqZ55jXZVixiDUwnYO1Js9YNOIRg+ZIrZ
sBWwt5mv+2pYnPY4EXK7XF1r8jt0n/jPv1HYkLZMUklHHn0wABjf0hbiCDFXgMH/wp5U4Ddz9KCb
9H7cFcf0azaXeDkP4j9VpJttOz0P0t+h3qrN0AYeUe2b+6zmt5d0z/2Fy4AMA5Sxh4xbR/6Bsv2A
udYOY7bhoGU1ryAcUtO9oi6Yrv74SjZ3yPlcQji3DmHS6IQDIXoqyrbFUn752DuuAJKB2lc0PcKb
K7luYKB9EOsTfJ9jYr9m/jHLCrHOXfOPiL7m6hleZtyCQ51v2N3h5qfXn2oUyDBfnmo7CefYdv5A
u9LZKXwtApkFJZLr+BfLUr4Em9v4IyaV1uEsM8fLALESKLGD9Ks+wTyQwIYJFoplVTeq/O2LY+Zz
XT3e2hs5aF0iNY0jFN5SVR1WL02pm1MIq1V8BpFut4kzNhsxYqTlIw/gn2XqktLXKTvdIKsZxVMg
IjXgWs8yZsgunV88zTDEvkHzhuijPtprlV/MUTXTVOouqIB6bknEGDqpvROxTYWaaXUKkBrpVEl7
l57g3id4kJ0Wz6tdltMuQK8OOeslIaqz/vgzclD1KLX7/emiZIlEXRZPl2MgasuWxoKSWa8LKB3g
T/47etpJnGAGtlrlGOJVQxRJCx2xsxHSe2nyBDR6woPeLlm/YofjE/wSUMlqfvgSDzaP/N94x4LU
2DkgfR/eI3sPd6wrzEkIYelJio1EIqi59D0b18nMELDOeXrwyWpCT6FDuTPxvZR9eCTv/DlKyDXC
qHpTJnAIcsJ59QpS+1DGnHJeBYrw4uCfxgtb9/J8ZeE1LGRGneZm3HEA7wwV5fk/HlbiL8c5Pvew
pB7/AxH6xlkVAkrUwpWCzu8892Cwj71AQ/xJRxEYW/9p43ghzYM+fltfM2ATKVEKzPyvJSdDa5R2
BUZpGZKzjE9Sg7eo2zOKsGhGcuM1l1bGU+Os91LTLbZqT89ofcWKlB85MzU6HbnBSlSmVMgC6SGR
z174+wnGvOrXYPfAUwONpVwbSdqWaHWfonLhwu9/reNn/1qQLrpqKp2kWws0z4n4cunN9xkU+eHL
4ZUmrpwJS5Ql9xqR4ajjfF2J30uv4Ws2GYVFNqM/H79NQveJDykda3ovDkuD3JetA/12ft0cUq7i
NwYq1Re8ZMzD3Qgqe0UHm0bJoKguLtq5s4lyFxqBEQU6VEaj2VWR/SazRqGc6nTY2AzIIx5OY81B
Zv2P+BDX8p81VZs+qtVaghWZTsUBn+8zilWlFl7mJfsGQEwvLYrdzbKeuKgvFr9gtExJ/jjqUm5e
4J7MsdCnpVTY57fzVjOti8MKriu0CWKP7zfuSfi1btxyCy6MVCGDGLfUq5WiIMILu5I9MBkxWeJ/
njTKTv/eqPLL+s6VhjTB33pjPv1zp32EJ3oLP5pN55uvYzPEfTP09kR2+R0aGHd3yavLLy/v4hfk
jAmdOCAmso202SW0kVeZ2LRl2Ul46Wnx5J8WDM0WcaW0+qtJKph22IH8tmCnodUJ8OJ7ugizjpf4
ZFz8EyDXDBIHPtH9L7cjnQDk9KpclSAynT1Q4XnN+ndERB2xILiIjTjdcK4u0GtTqj5SvhsFtT2J
GBLuDeUOS2G56soYdJa3yknIzzRfGFkV2yYkU9CbNh7HlA9nGHq7NHStarL+QxXKkblX710vO1el
1PU7M1a9eYGXNPXkrJ5tx0BQnXDJ2e/y4tVeY3jhjsVfycq3yk+48vou2aSLe+demRy0Kih9ZWV6
NqBsVHqNa2q5Oq7Cw0BPaLZsdzVW1NGTgtFPv/1HrTohXgFnsULxrRHBLwYuuFwlsDHN2v3ibyaO
bgR5/OcU46A9lkXxQYjSlvdTtlvEVwQhUx1OAuE7z/BJhFzBTcCTangLWxCb8Fax4Y+319U6/MiO
2NNpw3olvEC7sUva7pVQ6vE8vzj+pOQVpg897D4WZBB/PsNUwkdEVAsj64+lrMCZa+ihNYg+yaLG
6V7MX2p2Em0lsxvyJNx7oTNi/sEmsEpPJwR63KHxgw3egCL6rWHiKCu7ay+vd0bEuaee5Qpf9Aub
10yOvkxSGI7OcAUNw8i5zo/yuqz9TL+/Xu5D82ynGchm60p2fLHDP7j1MRQfi8BKtE7WlPIoaCOX
QZVUDS44F6NOXQGOikMlB4yAErtAPCuJM7PjccC9nCvxUXBfIwkOwj3KbNmH9v870Ai9zQn9ZPvw
8BMyphawHbKVXXvbUem79Sdl8FW4DrVV+GqGuttpeRG++eSC8gqusyhSmg1mJe39YV0i5HJBsdfH
EPozax7ftfIS8bS+VV6Dsssdny9lPxAnHxj/FsmCK8qlhygp4unmnlVDqc1pM3Z5G3f76PuwTtAM
Hs8+UPL/pvXfAq37/vxKYN8qcYiXfMRsqJhbROE/V30AK5wlPJj6yTmBgoNxjpPvIgqAUnV6xALg
tWqEo6cRen51JKe4aRx6z/s18MagzcVpb9iXFUUmk2uwimi5jqhNveUly5bfOIVbuktAYb3hmPR4
c7ctBbGXzTdkB+lS/XucP1nqQxQTQgLrq91FYGnF4olsXTqWtGsqZKNIv41haAIN5zeT38Vprs1C
o7XKbnocSrVRcTof+FDyBLgFmutRxlfJS/8O093WBRFe7crR4jS9l1F+LbaiCofn0fMeoGeynQ6D
Z1sE0aUOmohH8ZnRY3+YEDRTihEyfBjpdl77mamjphLEDt58utpbNTy8KKIluva6kIS+Cdwu4f5R
cPJIFdyukzNZXdR2kEpC3OPpVam7E1K55VNEmhv0DvI2+O2r/HpXPVPGQfWuZxvE4H5Ni5F8R+8E
Bp/SnzX/jvELY+1uPsW+nnwnIfURvUg7hYfMDB/4nW3TxcxsuJdxG9cwQ1Q9xZ6/L8WGEHOg8gtu
X0nyERHse9iI93M9lqpww0rh+HEDLmg2PSsvzP5ve7SUjNz19zxFFnXaEpSBzB7hz0fYSlfzn/wp
hn9ycIhh36tHD7d7M2oDJ7LttTXmjYPZAoRddvsy4NkFz+Pg8AIDm2c3FzviZykwEwMX7Mw7bDjZ
VWzYxiru6j5gn8mumusuDeycietL/tLT3wIVfqPBFBA3RTcuSib48k74I3TLEqOp2f69i+1f6/Fd
PFwWoeswusuUb7zsq42D2Vfz3Wo7nfu3l9LN7Ali5YGA5WVEijstYww7x3RMjmvBPQQKZ6hOU6gd
y47UECNi2fR1NEGeC1xZlIxZr5ZBg9NjdC+iny17GqI2+8/oe4lSVAFNbvD7f4nr+WyTDAeYXhlP
S8SlOUFjLgNaicr2BbB19qhj6rFJqbxiqrY5FCMfmo3hqZrmskNih0mIrgzr8m6SR65opujxgk47
TRsQ3MKiKAJ0ReguGKK+HDiTstQI3V7jFh/rnjGkVA6/EpLe3nwBKV7ELMxp8zEWRIE2QKS6N7QZ
QsPkmrzZrE3QwLboGpfZgN4hcSLbEGPHTbfxwA2C7+9vwa0Irxlx404sY2q2YPr9pm2dQHYYFBdL
CSOOsngwoGU1mdxl2r9xfsUVkS+td/H/GTXw3+W4lXs4Q9T2Cq9vP94QrUKMjecgVSDjCgrVg9d/
m1yscrnxEqsEFpCtdEvK9d2//N1bz/+I7CbslTaIpJIHkcq5chDjPSEveY76TQKiFDTjTtzuZvsE
sd1PuslOmkkZeddbTU+4JUKuGCyeu8loCmPaNFadYvyzML1VEzHUFT9LGScE6uhxPqI05y22Vwz8
99hPEDtd5os6O3C5uzcGa1pYkQl0rl6ENW9KroSbEJ686SdHZYKmIeWkxCBRh+9FIjTHgyqPXowj
MAXt/36bpbk9tqnpCTbga7nPkN5LRQXCQUIEvpHQ56IKk6SSxphuANEGzzkZxc2dBqika0KOkelN
ulIarKEwGz0V75ZzW+BkAfbsviM3/5/AT5xlIHTW7gh/Ji1rpAMPqaNfAnh2pXAGZLO+hyVq/5v1
66GWtr0FUerogMK40rTO7fqhMy55qAcxsv9cKyahslltEk2Afx3hGcAeptsNwc8V7LSpIEBZdmvw
WlJIZmHv5K66WzbY6fTGD4leo4OtbX9ZOv07y5k5hSKrfnLhvc3f57rhT4LzMRCf4vDWLa5fPQEO
MaNkhbdtVevnPZcjwiFCRSiSGvzDMjBbl0cUGvlwYcnEu8wKbW9ovdDg0cMrv2t2t4N0cTsRaDdd
6TFvjYkC60QJCz8YsCO3PmKnCBCi97LbtSBtNGf7dnK73uQBOqdZdSzKxXzf0cuetFGG6cTOESSD
iWLUWYrskRVQbUitwBdqDQLVaSascjmwJyATYYlOy3PFgDQQAB38qxMQ2ryR7EMxl2c+m/xCQBGu
p7gyzrvSTxIlBbm+sgKfT0Lq6PBUrc8+nZ3qXU1bwn/VRSS0Qy7FTDM91RGGaOaqB9aqTgdR/1Xn
B7cgq/76PwERJBaAIbC7W+h9PgOXzwP/vCALi0P3cbxx/y9DYGyDGfSa4cWD3xLZCQy60/1QcqFG
7AXTLeOAwqXuX3Mm2qX0tW8Zp79/BKvwrl6E/Kpt9lhbxgkMyyOe+xlOWY6N2bLAbhaATCwu/Ek3
GUhv3K4pfQ+OBsZ7Ksd2/ygViOneZpnIUOJJLT0m7BFzA5UswRNKVXrgnqMEk/cvRA31GqJAgKGZ
ogJDX2dqQyZyKvVCOewRXcaHa6O9brSyX+oxIiEHUBq8PvS5uRhcAnZIwEuMMkhf7LFjbOWm+sRe
xpGNMn86wffXvwrLaQJIwMx/Tyy+s57+2DmjS7MOLrIjS68mw3UQSPwDKQ0IpYTOfanPBZhkQDYw
8zEGmg+WvLojylKP9cy91CfHwSWBOMavFnQArxJ7RySej/Jd7kmu1Vhv4DT0Hinx16kqhXzYlfEt
wFwR2/E9d09omF68AqmkCZPobPwHbk9x/gaqKQU/p4Sk/mhyxPsOfwF2qPR3jIwykZE6TIOBSFcu
xbKjYTo4zNAeST31LA1KA1/x5gUovaz/mtwJUmkA2NSEf+gwSzV73p54q/tP47GtQfjaKgTtYfZh
NilfQw+DUgF1pGzQy5dICR9Z0UKZnqISDjpp0fFH4W3RsPaDEoGCVkKdo/csvvSI5N9w2DuCnX2u
YJ9j99VBdMS0WkTKDxbNXC3qe4hB7g23+KqgQbTt5au1Om+hXe+1cFngjAt8c+blnyIii4Vx4YSB
9upjwEbE3Yd6AOZ6UFZuwClfQu8+0IOnXT0ScXMAxb6r9oYKaqvO2pMdK8utf7lV09AF3kOBehJ1
sHcOAW0hdJoJrjZ/h+m0CazoKWvYdp4lEzisKlhAv21pNbbNmk8Gvh7XbhqN6xhbsJ5DngsVNqqC
Oz1AQ5nG8t7G7WsN/GRAbIyMBPoYtqipw6DnSwGxnfVTqAIAdyABLhdhorciA6Q4nlVJw2v8G8WO
DwH/A9CQSOPb2ucNGkBRFTY/QY0AridkcK3eyJiyHAFWI8hiej4ROpRnyloaI4KWisRS/8m9P41H
r3seJfE56P4MdrRAl8ue0yA9tu/sUkvP4bbagYTck392vf50uJZ48AN3JQ3DTagLuuCVmZxmTWEL
9hgW24t3wMEwtbtecBbTQscPV2WXqu562zlUeito6ns/0GJRffjk8JemKntRCv0ohkGLbz14tDJB
PvkFu0rRWL9tjOWw4eaxuna52BMA1x/RTsI9kajrcWw5a1Fq4AafBzjQAroqfTr4T/sjvmkwrRSD
qSZdLI66I0QzUxiR7iQSLMQvbc+bZTIfBROBR4smdu9g//Pd2FpiJAI5ambrS8g3ytcb8YfQh3mS
03UDYZ4o4x3GwSGBMncOVX5e/ONzxGLkJmMc82VZCUJnxMcGg+L/cTjVpsm9aBEX8XVkycEwhwUF
9HCXPS7p2+G0M9zNuwjOO2vUmUtquJRlLI+/8UeMyXHKEykZffePdCJITmHhm1MZAvisxacP37Qv
oU4c0PMVQsQzG9iX6YDWWwwF7WEd3NMKnv+XEAaJkhz4I0OmJxNqrBnyx1rktyKnvXtgn6kzbli2
OMRWLwOm3GMhKY6AKWhpmfY1IMTAlt+JHQlEXlS0ntInTBtnNGD+R7RoumcARbEfFV7UnSCU4rJt
8+p923/nCdlO01lnPa3DdHuKSnGsWWG8dQlmJhYDas+Ipzi219j97koqqS06fWe2XCk9JDOTNCVN
48T75z2GOPB35dHlVavAyW0b2n2X9vpz2n68uAbow2nR9+aSggWngyUUCgZvYk1w6O89T8DcBckG
HB3aiaVq51OL3Q73lUydmaPyMjNPSjE+/CYRun8tfl3D1XMBdzEqLFtdWY0Zd5Fd2mJ1/f2/HS3d
q5Hq4kz/yoENw7Tqk264NqPg+X/phRF+d/UOjZJLS2bFt9xB3Gd06bNVjpFbMndBYNX3+QJ6hnpw
hWa5Mih6OMJG4q1UAE1peg+QpR+SR/aOWAv1+45CH7ppiZvCVWy7RnAbcxFjABzvqn6N1t5nQdP4
V1wmOd8uj6SqTl0Hr4eveLs/JqMQ4W2nL8NTYXQBXkQpsSD6J1CqLrAYvGaa5oiKiWe0sLgxH98V
H0J7SVn4//M3tb8Uziuut0Fk2aNIqfKXKfLMC9Q8E5Fli6W7wNWXbo9AtYNvya3U4z03u6V+PlpV
6ObJ0MZsmggZJcQx2df7jdeKZOQ23hbjU5x7kaMEe7MFvLB0XIQmB88fSr48NccE8mhUqGsDMuJm
8oBivoBRXlsld3uuRBmO/P4AE7hhL4tsQXzdWzFlJvPw/vJLKtWe2qHo+f8PjzNjklo4TffBmzjE
MbO4PpHxuA2BMJnerwFkHt6GEC+P299vz8+DJ9gOogqs7G1siVoK7Sq6I4nreo3rgOO2Fofnx6JV
SlE5KOOUB8kqu2+qIaJeokEiutAEFjh0+e8yVo2viFL0EPYDay0gVedo+rLW4hWyBV0XzZZDdYWM
CKLAXC3HKfXe8Gl5sFXQX8K1DMZTLxLNPLda84FmRRpNYnsm0rzNIGuYfvNo0HRU+vcwR1dp+Syk
pwReTcNQdnLHpT7N+8JeU5FcbD6PU+eqKMMO6hoiYrhGIQHvVeQty3d8eGw9h4S0ELNzhRrUzTGB
+wxcbuF+X89rq/CYjWuNN3Fm6s0AoA/DGNhChJYGzURtpAYpK+4EGsVT3/F5GFagr+/fna7J6sdZ
OsxhCiIMyOiQR/qyY+KlWvMCoF8FY3MGZUPHzp49ARtrstwHYFVw6lcJmwHcpkDysZLN+O6FXSIy
9V0MEGZXgwlp8RGw6oxpCPCH+EyXlBXpJqGDBC+lViuwEz/yxoxau31/6ZTQBGI0ivfZSNWLeLut
rG0jtk1WOokVmP4Rbu5CxPsMnx+N9rm3TDfR8d71HcoWUMByBM9N9MajQARDobVIVgl2UWHI1j8r
V6vtxYHKr08oYw/3WZ02WI5DiYxprc0Ia9LgUBOnlBDwHuaiWeb66txQ47GMdzJLsoxcYmo9tADP
EH2dQZKblLdHoE0QHUBbX2uSXCpoHyfliaIoqqmk9bpX3F8zmUFaKpWH5NKbRaRDlQFpaXaAfVPO
BaUQ2W0Y7556mLaY5xczbJ6NgWEW3fa4JKEy1uGYFpDXvF8x4urry/gg07/nfG5k/RunF/2jjOgC
9vvEk5y4XKQJWfctiVYYDoVrgpOlbxunmryVN91O+o7f+18o/woeG0fLnMzzuQJ2ynQB3vtMGKsm
Lc5r1hW6S8aAz0om3bTEmvvzYlL+W7JNr+3q9VbenrMBfP1jrnA63j0d7qsGwrpDOq1FvWuYX+4n
5ZCCm3MIH7h4/JSyWK3GZYkzgzx6rjwedBI8/RWl7JvVLMGhpk2EDQ81rlzsqCVR64SU/9hkG9mS
mktFIjS6btMeNEPTNUC25Mvc78sKByRTxlm1e4b6UWIIBldgwZZjgI3e3x4YlOI+QPmly64BQ8OE
UcB+RVmRyMMY/mNbRYRaFpu3uRZZyzYs4hOFMIS90uQrw74ZR1ifd7RqYf2TcGOvCDBOXUC/sICx
xeMk9sKgg3410j5xGJ5ueZ2heqwbuzPZbLPZjeG2Mri+0fUOlK/GVlcjhLukYT7XgwtsrvWfLxyW
Ydc6c7Lu9YdgXP5dIKcx8Vbgbo8X2u4LqY7HpgRy3qBr3nlMaapPaioOs9atGh4FyklLB6SbCvZ6
bqDv5Xl0503DEF/b92pWv6asSSVIZCfzK2BuCs7w//puZhEV3hYJnEgem95Cyf0u8e7hHSQyBTpN
1bg+byM7Dv9G/5mKCr0XOoNW8aV/6wRRHsSqDjX8ZOr1c8UIPPoVzQMH6IE9SwFKEU9sLC9tv2rj
1Ac5bQGnVDdIsTzhPsNUH8PDONMlMztq8EcLW1d5FWtc4vburXBPzgqn4Eg1jiV+Ee3vIxyIyQcP
m8Rx7TlaVbb7UGSnWbaz/ArfQKFX6ZfX4nIWxM3sjDqjRJNaKUWaBs1kZekdznv+sz7bg3Xx2jjo
fNYORISj47JJam00jVLRk7tgx2SFo4rW6WgbOoNPOJDJ+FIwd++icV8yjb6DJ5/8OylpuCeId70n
57uGO1ewrLZoiGqrJTIR335c12AtQQzQFc61we/ZKzPExWN/ufhdwW6xatRDfwvMKO8iIwg3uict
+T6EjtQmH8l1Wdk+VswY8mqGSdE76HcHwh4HJxJzztQOcyKxNo4SX6UnWcVSWbCGI3Z00rtCTkdV
1sRnyUAQZ1BNaUZQi+U/jNJZzyjEzHeijJpzoNpi393y58yxw2EYEeoQvAF+BFzWALZ29J7bCJhf
a4kNzB81FDytGlwET96F0ZBDUTbUK9RcDiHgkuR1/tdYli/8D3n2hCVtHLKonB9RqPsTBa4jY0G3
6rzkZk/ovl1jKgxUx+hK1htdciecyl8M8b5XTUHPZXsKJtFMzyHJrg/l/7VGcmwNFZHiEq+c4mX0
G5pKZGovUQUC1LeVauBQQuxY+HyzY4+IwABrBz5BR1z5LUiKKozzfmjj394eQAyrWNH+MUCEBVSZ
/K8Gei/TBKf1Dow1oWjW3TTDz5VxzArLuC0eWMuKRlXi0H8/NcNPaLuzjTIR7+BKlD80ZuV6s2fv
wlexDJyR8x1qNE3mUNgyb6sRyZ2OIjbzH4Bahsi5CcSBG2yCXfsmkFrLdziOPU5XGpJAv4TZe0BT
bPd0kuQvXEdlIlUVISS6/uWhOsJBavEUyGc//8I4JHD3gFouSkzbGAJ0YAOIWtFW9qOqdJKr3+HY
5CD4te2Q2+IgSpAyH+OKc8+WtNlK/WvtdAUjzawxPEqhyCygD0kGyAAv1Mh5hmrpGpjMGzmMnzbb
dTAqHviozSjpJfpLV6QHXFAHYjH7yipK0DBJykLwZOadQQHaN0EW8mrcjaSyl0Od4T5bLi3TMoAD
+1WAHkPVvG2xOmu+bn+GCu+s2XMjIyIAOGQgQSBhEUzB4iquz469ZaxXM8stRWXhMjD2ORS5RDot
zxzw1Z+e7onmbacIaiwOXu/Kt6ecW3S7mnUlPEfCm8lc726u1Ejb26ZTnDwbAes1+UBao4d/dDaz
toQkCYLKefxVkR8MEyVORY27AonRhJ3qB/ZfPJOeLJPxHQo5X4ldiwVy8w3E/FkGqLNVArlfcdPl
pW0uLSUXsdEDwcI4Egv78+Kuk4ZJyLQ6XYO5mscfef5DmzvLTAfup4h2VJACZNaNmwNVCqAoHUOn
r5am3lHGYDMWht07nc4aGMtXhxLb1zlSeSmN3kaxsu+8aKdpAV9TXW6DxSOvNg+3SHYIL3Ku1RD2
t8+uU1UU/cGtc899xNjYF7e0JoZRFnanwn2QgYEDo0c09WpK60+153l+V3PSDerluSTVnT0f2hwz
0znKEv5GSSRDS5+xlpL6s9kRb6bbOxa12zwYJtrzeOUviZBV4iGlCgMMAZG0pOyRq4zoaOJPs1sO
6A2JM0MwM/HjxwsmdROazJcvNxFpcvVTjREUPce/ACCqKvgyd6obF0RnCh0m9abZPicFzv8WXsh1
Sg34R3JYxD7cLYbjE1AZAodnh0nMnUdGl5FA7sOYS77181/SkgbWzyxGTflxHr3kXnbD8M9ixwVZ
LoC02Ci16Rd6Ytu2OWMim1aZqE1VEu8NfqL1/Snx+lN59Zo0D/rTfQ1GTTdqpV4fesQGlf7ViGfu
m6irbk/neUOyr4cbrZfZUBjsuS2+7SuR1KpCJD2h/bppi6hbLBMFyhZPdvE3JtD7BMlvJGNtxoo5
kBCDUTCjHth5Ws4q6TWgNO231gBCqK+aWCIClsLX+Z0eWcRAojocp8V0fLMG31Temaz+xfvMS2Qd
05Ju8tV0+IYkcM4Xunq5NLa7BeCgRPGpXwAozh0FocKV2iIq29pKADdn7sQeA8DM6CFiDhSisIY7
hcHlWWP6wQZtU4H6Ial0zuX0Wn34txHMUlAnbdIBBgI3EaToDwTuELd8rd0e0WCOR5KWyy/Rw76m
hcwWhK8k6vqP2oEJ1S2zY+q7p5uj1C/BpGOP7TaiQwhZM3p6fgVBjq6xByyP5ZaioGV3udHp0yXm
Sjj/dWHz0EyFEz8y5Bx3biIXxFmjRdYL6x503shhmobbu2FmgOn4CuMEqGNoDnkhYTstF5NQecjU
XR8rjZYZOs10fuhyseqPMyJrul+tyZfp7z/EzLn6jo2p/XuEvaSyYZ1I3Hvm/hjV9j18y+xUSd1N
oGuivM3bbuHvOgwAMDRUA05gerdmn9GVcGL0uZWqhWoZG2ycw51/7GoY+2o6mj6ScclSreNDPayq
O0gxMYIJTRH3+JwO2g915ksB0gbhZ3eXXknbOz1frB2q+OpGhkuieQIRsYnv0iSSsva1ey0UpWug
5kUNwVF2mQ81MC1PbUqxEXADhZ4Tv2XnRKYC+OXhaA/gt4asPdmxksQH6r5HPco4jpOiJ0cvDdgR
rzTRC/36rh/mtXa7mKweAQyVDpYQ1z/pVnIejv2RENDloDC70tby1I1/usIe9ovNNty68ODNG8md
H3FGfif8MwAzx8lqFP1cn5XQVyOHXVVZPenp7XrnLLIrIVaxirOMqfCuL08LsEkQLRmTV55zgYeN
3rRnlFD8x21BIaU1ckcfqVZboRGpknUoZDI2Q0DiSEAx7cBmKVkuWGAcR1/LBatrDhFNQFS2Xh1a
kyH7NFY9S1mPXh7Ndd+oMLXK3d5Bz/Ds9AaztPhw9UtvBW2cEXz3vkhN5QY/Ci5/ZeTKuffWeGlZ
CgCIr75epwznygctCo6IQ8h/ZqMxZqhLiVNWU0ix+aV5tbkmBRcchRn0sePkXjS3tmaFlHF9OXqW
CKbvnX7U9F22mWkJtjyoeNTDZP24xMsn8DPHYFS303CW+OS+qiFZY8ZzHqUNQr4xljrpexTJcppK
07N/kgzcnNqVfAUJX5JbzGC7dX2uHC3E0p6NH0NUKR4gj515lY72uEZT8Z9DWbjcZqxC+LSaFavt
yC8fciRoSrWTv6+08D/F056HvVHlynBZTflrnytVZomht+LyqwXFykKc3Epm5an+d7URo13uhpZq
lmh/JfL092Z5IbwdvWpCe04DAsw21h5MLieDoqG7CZorsyspiuVQz3C9OZjxBiLJPWH2FuO4iC/E
iSWcYfgVmrWu7A8g/C9Rdc7fjzWO+B0tkXRdOmS4gLbbJ9eEWAY7hP+3AXXwl7DtEvw/LvEob2MU
0JjdaElRpzlW8PSZpFuwn0o2OyIvOokFIacthoYRXMiKHcP+zBIZ980lDWCHSmrpiOPE7BCDJTgf
2xtTOHya/59vmH+Yf5TBEg3fbayqV1S6vzK97zemMlH1ILzzhrH4id6hdghNA+ZuSLEZAEsNB70A
EqKL4sjcQkUZYd0bhXBiSNbMrxz7aCbIgxYXKViIbRG9mAv4NQiOx2u1C8Gl+u1xfgVvQjw7SSHg
JdqSTzeHddKh7xwRQ4YTIRiJMaz1X8+NHy1BrLmgdkXMnQDKf5Mjuim2uonQOK6CoZDOYuWxsU1q
v+VG6RLMhXnB9VRyhH/qqbHPBUhshpbuT4i9s/8WvXv7RvEVg+Zwb4J9Todp/OHOOvkandgdwcLv
uoxrE3g8sJx6lcrTBTz5DzY3Q9GjMG81eEkiNEpVe3kvKGLYnkNqfizr3Wi2RCLU6dPpCpQfNhMp
IYwJ5YeESSjBkCzTRSvKMCE70IQIX1EgJLUeqpr/4iBgt3zMEdr7Lam5Tw71gydcNUJ7bIAnFCM6
lJTWOwhjljM7fQIz6lGdRe6pgCGZekDGcUi5V90ywyMPuPhSB5Tn55BPaQ6Ly2ywr6t+QnkPrqWs
Rs+Z2ZrYh0C0Ub/lZHqldu270+9iYaiI2JCAZ21vpBnC9CKGMoLtHV6uwI8YnYnR6IFi46BZyvRs
Oe3dQRzfzriUkN1U+YrLcASvYrWq0wtLhTRyQ/1G0xMDGQC085Q/jrixXs+BtF1wPP3zxXlzcgdT
Qxd6/zQ7fdUFf1vOtCpcD/BuPEYof71Eg6vbp+wI/ApvigiYGeZFzjwlqI1CYkNkpxkOGbtO4c0p
WFIs4eXPUZS86ZBKTw5f0koSdNI0lxhS7qcmp/vn3xR30SeW0LlXx7zP/9waOSI3CHUnxiCkYl9+
nc5ka072D2u6sVYcrcAOH9WGZ6wQv01pq6gO627mjrAagv2dVPWkrMeIklGXR6/34nTRASNx4iNE
gu08HenQHhh+1KRHUMUYDcNR/aa0+1anLJVIJNq723GOtb6ER35828mtvJGJrrxxDUfoP6qjgspH
WtPCNZ3T/bQCCQTb59r3WGiTGptEZTJkXpBZKsfgcintfEdWoE2vUklNkj8ZrEZRU+4FWAfNq2qb
usTm4hF3EVVQK8IZkfHEH/iRu8TnWxE9UkKNvSdj6WlIDAYl4t2EKwURrXKr5nXGy6C6VA2H2MMb
lbg85dTsOzzPi3Ayg8JyUpe0RaKdiA9X/bJuwD3vFn4s4Kxqa/aKQ4HbcHoZwmYywL6nNVSDM2ij
NzuVZrcPEyiYUpXWc9EvMFTH4F1yWOOWdbSx/7Sw6yIcec7vCC72JZwuQCvnwKt8xCgbYf9FrwI3
oqFYUuDSY34NNW6xOY6xjtI7u4wlk8sGPioGkGP1a0zZ09p8BpAkokC3eCa4D5/j6cz+ZMEoFFCR
5c5WIVQsO556BQdmf+v6Qixs+RFQPb14Yukvlt6HI26A4xgzLEG0SPdMHkvitg8pV/LPH8kHZlfJ
SWNj/Pg/T82MUa/pjnHp7D8O80bgrvsS/39Yfkg2KIxM1kcZwvEGyfyZR4Lv2cOcs09wKmxqQffg
1kb4huk+6Y1vR2ZH+8LNM2bc/7JXyOMComYlZXTyTLLGs/1q5ePKbp9m3xDixdQSTXFNKSezWRfX
32aHSz0arD2cNZc2sOQ1JARoh1clIxe3w2wEgECsZS+NMe9jARgHMd0F2e3AN5FbLpXQKOgNbZl2
O8Nf1nbwJ40sBjC6drw/Hw1n23MnjteMqS9Jv0PyGpC8XKNFQTWxd29w7KEoZCWjkk4Y3qadS20M
5YLpvbaPUhV5JnvTdBbFvCi5ojG6yXy2Acy3ZgWug7nrLRS3GGVdR434u1PINDRmPeBHMWaCAEPq
qRGt1UnOcZl99Y1452yhXgGEx6L1zxbPUCjrQa3whx7XFaXNnb6OT6b+LY3Cq+PRILhd/wdFysJH
3+gl7ogNsQetXcXbzb9GvJ9eO/CMliIIfedyOOvhuRWq1UuB8dgQwPeK2S7g4ygjxF9GFse24g55
DNF77hKbSBtb4c8zuFs7qYt8CUZWKrVM5KP+CkphwjXKBy8vFls/0urMH+Kh5MjLP679qYOhW46t
qEQVRcuB1SGXzCpFGUm6ZaMEdQtuDTeq9WZ2UOh0HjCIVwNk9J6ucmvqY1rA74Z8kVynYe1C+I02
m7cpahp4LtnDc8G8bI0jMg0gP1mw6jdA0eQxPppJNrOgzewdYR+GV3pGOEhJZIpv9zvMQEnj9Ho4
dm3A2BMg0qSAz4K96lAwYyJRZdj/gkcn1+qQBFaK0Ykoq92FIEKq3uHisi2y5hN8e3uL+Fd6GGFO
sj5B5C6WZ6be5ucJiqUlVbtXwrfIMpMlxiurIHY553wSuOih3/bx3rXmGunuWJwbhkpUijxhY8XV
eviKwTG8p6bibF51dfkQ37ld+aYueYsTjCfZZ5Dmm0epzkZn2z7POEIr7xdl17U9QWERWxp4Fbwu
oQWf+esG4XW5+SoTHxMl8M2z57zWTS7zDwyAVXlxr2u8Fc+ddLrhYcvkd99hARmCgOLM1oRppIrJ
w3krQNqZ/xa1i3mge6XZJOdx/4dOdQPKs+itjuaMp1jRllwuljPU2qnoBddEC2H8MCVHh+8+ibzl
fhDHgeV8rEvLy/ujGBmk36x8Rp36VaYPvB6l/UhYRLw90x1kvkCz5LkZI9efVfzydZE6wJZOfOHm
YnapjChEyr6jP68eYy2k2JIx8IlwxlTvWyrE1Uz0Ts/qvYD7H36hZEXW5a+U5nqxcJ07jU3KZUXd
YifFLqv1qTDjaJP/k59Qrj0aIl7KERWEdA1iQPcKqaAPkhlAyn/KQp5fMB2cxdVbo/ky+IGIauBm
vNr95VN1XRJmASx8biDJMBuOWlYM3sUjXKD3jBWujpaS1uKOuH/OheEzm7NjVUq/IzgKuf6CddQ+
4PeHTjN/GqX4Cb8uEo3gonrIpsWfMOLsYoSI9iTh/+L0wJje9MNcc+YRgR8nJArmkxE5eZoutNNn
kEvPwf6/IJyYOrgJ9PXw6kPb3jZ7Rwpv0oKpFJ6OiIKMnCyLwBOIeMtHcHfJ4dAjHdAd3hgXRfDV
JzI5CLbbIiuNNu/ZubjNEYrKOeDloD2YtgtzhztSyolGWhMYmEFIEEs/yE5EgcNLebrAz7RJHKsp
TXcpOJ+InTZOsYIiSR/xFAWKN7UIZtDcMKoSw5zXhQyfIBN/2ZQ/cBm7kwY/DopB1Y6uUUhREbg0
N0rHJPiZhLOI7gXM5XI4R6W11Z47Iw0T9QiKKzfo5PD8Ip44Y52eZTz0QCa7aH1T+Nt6l3WXTnXU
PDK1gclq1inYuep9+Rl2pfRnBPFqYPOqVF5NHUBN47j6M/fn1iRzR2gVRhpjs5BKj0vMpr81hZHk
tkQU1Rz4tjS8N141TFb3zlrRHapP9SYabHX4hYBmEQk+EkDcFQxY+7M3xpjzup/pZ6pJoUb6L5DB
/5O+xmCuOvN9uzKHZp1lDqhExYsVSwUb24cTtEokFPCfRIG1CNXTwdmU3M9/W3hqYXWwZV+wc8Nd
OSX+VzitZu6c5/YM3rPuYrKq9siTtUSY/HM5/MBLFB0RbDo49SpR4ZPnXpe4nCpLt+zdulBUK71x
YT0nE1x6nayrDMaTJSsHSuDQT4BypoHZEmHYPmlwV+vL7hJ5n7IKxM8o3Yd6cj1cVJbu5ecf6+1L
nZ3tznjr+xjD5zdBpbyNDrxKJWYtmJNgxX2Pki5tHJjYLBNVdabkyFHlQVHmZS1aYkuXIlljcrtf
iAdhK125Lko8g4dHCgbnbmV+dh5zbWkomAshGtawH1aBJ1wZ1Uj1xMtRcYQJYMe+Lf5Mcu2wL0Av
0KwDDgTOG0ClLQ6YPSOQfecThrBMohLHIoSWDzavfwj1GKi0ad+FOeDEJqTRkf8/6AqRoaqOeYCu
YbkOb7yehyfgA3NBf7YevU2EaDHnVG6D7eMnydphgsXyAqI1sbe+cNCmhAGW+3uWAiscKY9bLl63
rJAZUJ0WdKdueC22MhNbHfpNRPzcsUNUFc6fGl7GCWvz++lG3XD7P5jUL9WV17qZ1DPC3Sj5/2Z8
8Jhknh9O8nlmSFMqfZCX504nzvk+ylx3fpQcSvse4wrO+LfhhplQBjTPCQP1FjyY5XS0N6p9OUVh
flvEtzDNwP/pNK1s03398kj1XEIN3FbkPhHh5Uwi66FU/kDY3KNvdbNVHPljqc2V4ZdFLF1Ti2gT
5wfQXJJQO2kb0QfnkJCP8IgcmK2Dt5/ZOdmq7IkiqANjmukLjvhQgvdJfQsy8AJnnMoFpxfOjEhi
rdq9EiEhz9ik2OOLTrwEFwoAQs3bZ+waNvYp0EK94+78gYSw+vyIgb4FMJeMlZ25/bpAF+1c8Pq0
GKS0YPIDd6MVo4va4gRbapjcbGEuUQfFjTikUHYi+oNRQywK745XQMQ7LKe7fzuznsKbXPlnAV8L
xRQpV/otGwa1Lh0F536XmLrsVyx+7VONuqXyYsHz3IxOn7SDAy53eCe8uo3Cyw2vmnCnGp6XQK7s
t0iccaYY1LTP4AsxKlMuXCCs+w0Rx66gUbo0r2m804dYwJ+TLOty7djESMX0aqy6PW6XoQrABKwZ
6dGP/JNTQ3hTs07sQPo4nkMXsR7x4eriYVHG8N16tkxJXaRG+M1RUUDnARr0eVWbomclznCyChr9
2ndpWQXNqxYKXWPTRXv+fnBI9o4RJrjor19ACcSnCoVG2XUgX4MAiS57+cQR+JNaSSo0fQyCnQai
BvVpOWFLOPPobaDprv+EV3jUevyVxsgEZhE/sL2j3ZxR/XkVGyuIyGkUn9G2MmE4Yo1sdsL6yBc2
DcXRYcVs+W1DpWorRJXzH4thBuuukKE0DH3KqT22gr7CErHHFasRXhUJXLht1Ynm6ODKwSvo98aq
5STHCPBhYqj11vMa3TXR1bsPLSKSbvljIOrZdjtDriP9t1490rQZ+hxXmtt+v0gGy4vvNOqrv0Yq
FxNUW62WW7v7rfWzgnRVD81Ffx6v+q8P7IkOiEJ6zsIGu89HLoVmQglZDJfVv3+mv3W+ej38Z6PH
qPN428D6tTtCPs++kUCWjYGkgO/1GqKUk5DGYaswRjLqxJfubGDy4bbTLxEoSQij+wJfo5On0n6x
1738K+YoXDdJjY2BPKf6E4JBSpjWtx4412bilLCDoz4LfJu7y8HahzEdjIRua8e8Sb7AIx2aUfsN
/kA/TZgGk4CiLeldHNKA3O/k0upLYN9c3oTgC/nTQFaL5BSigiL0Y0UEe/bs7qCjx5UKtuBdSwVb
6rBMnLt89IgYm9lyaZ+ZJVx9Li6EtZMZW2cV9UEBO3xCWJ1TGGHH6cvYB17JNMzgHpCGtyu1eLHI
jEl4YJXxErcW0LlkhMyatDMP8stg7POAqXZ54+p+l1HfLst7f5TC74UgGm4prcr+IzmzbIKLG460
PmgC6HGWYFu2zdS5obXtSfDYKbzTFDi0ur+y2UuaudbEowtw+0hbajkc81OJEc5IpJ87p6hrW0Jl
QYUy25B+GjxobMwzIkk/b7v29f4GGib1B13tnFTvu+5amfG1mfKbzNLtmra99aQMbojaAMY+cTNB
2O7AfZSNNnsSs8HP9R9Ni0JQNIRrmnGZKBlNjU/K3vk0KGNKm7PrBntZ3Yg+yWXfgjz4TlYbM9mi
13nJWVtNtx214uUE4s5+AkUpOJF209dFz4nIMlIUe5wBVLKmN1MzfoqHqlQDKiRQwCpT70exogw4
tbBH8s8uIbHO2aghNiqvgDelVMEVDPfkN4mIvXcUpLyb2ld1n9xToAsI60vvOXP0qYT8M0Eos7HL
TiihtTcmDYmIkBBsQucM90e1KM3mDRp/PQqzL4Pgj8RkF5uYWXGXaZwD6i4sTRz2e/fotOXeAzk5
jABeU6Gvbu7C9LTIRKkkWirepXHHs7r1/dAaHUV1y8r/JZ0Lne7KwA2lKmFwaDW5HWcTdADGDldB
HDpWFJfVzndGP8JxSGmbnzxtELM/2FxiEnWwRkFDzFnx7lCWe7kykSnBWKXMNJ6uSsh6IvIQOKQq
In/iq34/Q0mTEKMNUNnBEL2fWAQ+o3jGctaV/YIndZkYwJFgXhreqniBnLaRjnhUdhZKQNt8TbMk
BDmKVVyTScXczXIRlfGE7+2waRmfTv66FEFoxIW4Oorr/oTOWrID23+yuYPK58ffIOVLAKmwsWZe
4UvdSffn6b6s0HvaJLojnvQOzEalUxPugycHlA/JDgFZ+xTgw+4L7g6XBsX7vA8lX6XKxGzt8IDQ
4OTqoyXdpYrEHrIANeXM/C8dvTlWwGcg1zknSqNpXbJIhNz2bT6s/ady6YC5vUhhI1+CPILyL+Fz
5OF+8gACmkE5vbumObd0QIwdSZVVG8nrDpPYnedg+ETCdBjXYGd4Wc7Qwf1VctrU+jbnXg1y/RuL
96JPO6oFC0/ooT+ORs+S8dkWVuhwERFBkAIKZBz5UMEIulqMekXHO5RXHCXTl0ay5L8WYD32tqch
gfBSqscQDzrhX4+xsm+LUyOdpM7b4OoPhoQfsmKP8odvh1HBMZ7GepHYIV5e9VhbVq1Q199/tl4U
YRk6RPWAByyosup1iB2ei97ZzGkjUBUqkzz4H5AcwvfdGpgF0dGA4UqSHTE2xF+RWCw9VB8w9ljm
lTq61R8lZ7XQtZvBRP5Xh70kDrACmj9TOqauz0imhyZeouOpDpAT6reDB5VJqrtheZnIaAsI09Eq
JrgC/PTEx+53UErBT2cveHwTRFDyeWg6yzwuZDLuY9pXHbg6VGIRhsT9ThiUBdsTvAAuzBd8urrL
7mRNDC4EQAPoLgyXk/ytOeQYjI39g5q2wF+dIvMcHFLAIj6nUIsrgvPvL/I9wZQRBHd4ni3u90lw
r+dvMPyRoCQcrVUtnjIYr1smTbwjmoTqqEfR4hQg9wcjIqYsHm26LTXbzNVdCYuBA72A4iXF/lpL
Af2OhIic3ECoKj95n2bfzAU+1d8W83pn92lou1Bvwl700dmMw40OB13z8qMBlyjZDUY6PpfgVQj2
/PuU1AzW7yZMJH4GxIjw58Jv5QPHMRqWVgWQUqjVj8U9/4hgFxRNZ9fd+DD8fETZysP16QpgRNhG
mpYfs368mhijn9yK69cqTADg3GuITZK35oAWhab1qJGUZKGmO81mNZhuKhiFQ6Rf6dKw9Je2/DnN
8TRG0w94FilmW/PVHHFtMfSkdxfvnLI8i1FdlMHEnCrGOauu5yCDokAt/QFik2a9paEH9vT2Rp8J
Y7y7WlRUM6kR3O0XrWL36jH9MjfcWA9BK4zroWy7THbET/gpdVALDnLFe2dZyt0ghxpzqRDcVOIK
y1zLADqofAVknQpDbWmf2IecjM/Ydl/nFw0sihLp8sgQov0gA/WxxvHhrFnZwvDf/rKhdYjWVeZ7
vL9sgPQUy9uzeVjjgwF9860rrGbvZmUdBz1HxSEfVmuXM3a20DjluuJ6Ax2V1i8AZ38YjOL+kYn4
yVxpF5cpXAzvuAjzjwejpkODUjIQ5WbupgaCBm4lHbT+FX8JK1zbbOcNzGo2Ww2csidwFFwGZJTu
mRu4I0U/g9Ynu8dZn1ZkdiALp65cXIQlWX7Xq1sGGcnXtk3JiHsgAWCpzumTF7q+8sEMUe6MkKra
tXX5E3iwS6HZFJDgNyAKTtJCntLKd/UICrTI2BV1PPPtihhhD8Cyf5oF+2Qj3791L9t9n8pFgHnm
cgdgfUgKnbBoHnoEro9z/9SZDRLKpUSAgQaVnsPSnZBGErpt31GIz1fVoaPZ9acEHnV1HYP2QsaP
3n/eE/4uugCqrrRUkbROJPdCwlqRZUc+d1ZSqrD4ppSGJJf+F5bBd5AbXi+nX1mQGFzTcGTuwaZ9
2rHHavHLzywvsioJSTB8GKWAUJ1byllmfLha/Tc0EuHjfVdmrJzUR2SFryEIrcbzvxYvFYidmCG5
8yjLtYOoGduzv1uibgmb71z5EGn92jqzV8p1xZf5w0M3G/UtXPwCV2s327oFV9XkdYhvUm70VcJP
Rp0gL8qoB5UIEY5LkD7BQmKUqKxaJasUdJJbvp+CGwW+hR7xU49F9TNvuqkRuranYoR1OAUCc4mq
vo8hz9XtukHW4k23NkhorU7gZF0nI+e0xY0xalbpl7N8u/eNeB5XwMlaFFu7w9zcVg9cJW67fzK3
tLm2+FJJAW/KzbadkJcrq6Q4pjMbM5dg+FJp4s/D7G6d6ayJKjHFP5OFLHkUxVgLROL0nx6YRip3
IOZdOzVCSyK3lMXnxqV/t8PFHYC4rCdSfQDEfhPDGdwYfrxQns5HMxAjqfYUmpc1zFN2Mh6cqVmz
QusFKqKXpcYOu+SBi0vVpQvMOIAYmLWGuioap23MkeDw7ghrsRty7UNlR54eJGh06bapDVgo/8z5
vknB240CVSj94dWgN5O8FWUlSiTNa6b8pmIYJ5JSrqbNzowynRWSQf5GRvuRia3O6RXZEYewEh2D
qoG3DuwBr+TsU68YuVnkrht+1Gb80BPtggSOaKjmY6aPFMMnc9bIoPHFac3pFrDr6Fd75YKaC4BZ
ysjbOCkN/cbbFErf2rcVkTkfoKwMQ5Zl0i9juneTB9cAZLpyjHJDnQsJJgUIwB8x7bRAWZTmbdZJ
Cz8UgaEf/4YIj1djuCYem3jhGkgBA6NvH6pyuesvgIGzdz9Zohwfavt0XXCnHosVG3vECuD1pp/i
95h2jXZT0YhXNrLnF8093qaTjr+4mkgV90L5GE16+Ue6yvEYj01HFQY1U1Icy8Dk9tppJw5k1cEl
CQshVnm9yqJnIx+a5T2rj21TnrcYrfB3/Rgm/X+QVQfguqbQJWEBvEr5EfnFIDF0JLvFhTLd9S6B
JtnCxbJBrmOd7KmUgjeAza/Erp/BocwORDyu1jpW92kavkT8LuSbZRJx9rZbtqFUP0kVoVoOcirj
4ai6MWm9pnld28y+IoQZV+3TXeaR1H85aPhBNlMtmBhovE+2Rb4grU6EEBF6uHscF2uo/dRZjLKQ
fssbL9oetMn6Pjaar3xft4fGh7W3Ys5X1BcpgH3+8yb5xeqK3SerlYd8McPV0L4TxjZ66fow/kr4
oJtlPyvz0YE9yZgT9GFxRC/wtZ8EmexxBPuGoUA5SceG/aCGx+fXGLlqaYnm9uigaRqYlmhp90c+
zcOTAPcrQ/k3KPD3H+tYGHCdtDhU/MwahQnAaQj6/pUrFJ9MyHirXPZd/FzcngcZPUq8C0QkUIv2
lTDy+dsPObuV2DASqjbdV+oZL+aRFjrpF9jQeWIdm4klvbxs62fsZfCa1JNIbK8fC20pRBEoNF6U
0pGu9x55543Nj9UcBbivms7TWufxcMK2OzR4ZbR8GI5AZst/sUXduZApyyTjxKsVv2zAen0MY2n4
2gT/z7xLMPcacDSWUPxFW6e48+0o+T3tPTWJWbopWntL73/kFH1TAZt6YqLh5ftKfxPKvVvYCBiz
YCYyggLJeEDobIwPuIMRapKKqUrMIbuRFNMhUjbBXFu4Ir2qS8sgR1AAp9L5uO62gFFNVmhNGyAh
hUmpwnnoswzcSSk7/aBhMcAXB4DT+vEu+vxjOP5afZO1Pziaa19snUAVZvzhHFu/3uCbSibwB34K
kjKnBJInaOMcdUda2v/3qRX8Nhx+O3FkWRbYwn9s6rW6gJREsKBh42KZJ1fSKlRIy/QAY3AEMu/w
kkaEhFNcWXNXMAYQOVx4dbn8kaV5pOySvPk9GmrKfjXxClpMjQCpXr2dzY6G5O4D/2ZlqURqNpXJ
lTokK2Mmi2CPwhrBgn1PJzRTtfl5J+oPFSCharwLGTXtfPZNuq21GWNaY0ukwJxzZZ1Se3rSiKjZ
qTHds6ES4iRtp+k77T1EMVGgccwy2XbHUAnT0XCcLMyf2JSZheWrfqFWQVot8jo8l/S7FmVGmGAC
/Tkz4k6WhOnogFHImVwbkjHUv2TvZvezUn/7qp2unnoyEscG1e1TwBhwbauXGQ2j/xzih5vo9DY/
FK8cHEQRZfXrcDO0h50A1T/MAWY/C6arPeHtQ9HR0K+Fqa3sboIN/id2+xE8HipvdmbA7BBbLM8T
oq2PCFnfMA94ih+swSjOgwMvkkcPB5enAnjAVp6tMsJW8uciTLgPTDpe+0PsbwJC3TNBb09d5ZdF
zzL9buyx5y6j8NYuJCVDovTSdGehfhKLo8P1cF8TEsHBNz/QK9OuM3244f/jAE7FDtonaXrP9oRp
Yf3xn8b87ML/kBS/JphtV3M1TqW1s1HvV63tbXuZI616q4L3460CZVwbDVVGK3z8ZJt2olIrL9v5
pK0wQyqmaQTzRlfUGr0PaK1AmFsQNfnGItMkC7ea2/gLrRk2j3sjxIVKeiCO6rzaOPa7wFsv3Yyw
aPHxyFBDgd/BH0yrIaEq/w79/oI8YWuLtnklXpSh/NkViMMjWK8TBhbcPS6pmS3Iv8yP+AG6Opia
qf8L6q1A7atpidqwSm0iE0nGLt75h57tVlC96PnObFHwG/9/ridrj4LEA1VrR7zeUK7PTIZMcZqw
GtEEc1+aTF4Ijpo3T5NNfaq/zzALVJHGiorHjzBCsvhGDE6GKNr30H4YEF3y2H4FjF7KEeWh3bjJ
rcHCQW59QQ2XdFhKm9WjQHPwEdQlIBRQjyZlDbHDQQsuNcFosfAZ8jrXTpY9oh4eGOeTRoOE4zNL
xYl7gMUMEoPt1j5SRSZC2cj+chGW5D5wFkntlTlKWwtX1udCWZvbSBc+Ev/QODZs3N7vNQPONn7n
2aX5eGq130Ml8zixyD6bnfVLCNa9JLbiWXT0F9V9dbdCRCJW7VWgMKNLSimNfXgWZl5PAhU7oOIZ
iJ5l9Kp9EFIoGtlYx40L4DIO1S6JskCZaBjA81g1TroSlcf67Gl5cT147TiMnN/xGKd2v72bDfJd
QJDIHIfJ/+Vfpxk9T1ZqgJ975UpK9w0YZQqm5orA1a5P6DMevMdx4GoH3G56mX2EDwfBkX1M/KPX
0GCSZhTSg5VHgYW6wxI5rJkivPM3giVFaM9fXi1nq9joowcPtDay/BIigm3RtlQ+H1BlQFqxK0mD
LARD7VXz+nmkDgbJ/spDxZJgB2T602WPV1Qx2SuzBi70X+v3eJwZB5P299LixHvy1bkE/n70iW70
fyANdxCriuLKbXT/2xGzrwrcgAlEg/7/N+mU48p9H6ewD71cmgN8Fldj0ORUyyHjbM8C/BHjFXDc
yXF8vpvm5g8IY8BNH3Rv5UW0kpAsfgLmZrxm4610Khbe95l/JAjMUxQ9TwZAF0s11WAYz1hzPa3y
7PAOmMMORnTwut82IK0EJlveKDN2I0e+q3YxkbjTBSjDH3BmXWaa1hdYxkeVt9VS1CCabbbDxJ9G
HbdYxJC6mBVg8lCembDe97RfY8i5ZJW8gSCyNIQ7300KgJx7+FFMzMJsQ6+qqeR9kXnOCD/PzO+4
Bbnpj4DKHK6s6DowqneDSJeRgT7s5ObQ0QFNFiGqD4WgMKJwvqa5373DZF9D02Nuk9TuPjqvoBCg
ryjOUQkD14GZwMFLhSv9mIKNIk7IS5J/5KrIiJv930bMaLalfRxP3ae9AFNxRNO7cv1vOxMm2FS6
X3x8igNm6nMTxvglj7vm+JrgjAkCXb4VJDPffgWjy5IPOXsoYkKSnReRMY7DNDPUD5nYT0li6kut
PnKr0pCV23xQHUWUqjht9/DQDp11x1F21tIcN2RvRNa+I8OQlBstIPthewB17l3G1qKUf29jwJXj
Bog5QO6wKy/N7lU2onXyHol1SN++4YHoqoiPf7pKpow3TD9KZ+A+VEyQzwsXyR7/KCOl6F/S/wJ2
fvMaEqi7DLBuzYUPHVXQPWyePAQPUONjlhAmcDfJAFClXCOXFTSwMlX4SyCSpVhtdZVGmD3CW36d
m33nQ0Jtsg4CoFpwDVU/30Y/oIllUZxn9b3xSRVuezEwl5TUX3Wl1q/50P+DaLNRY7XNrQXrLEJA
3wBon7eE6EK5H4gvrhGxwQYHb1eoxnr5LGyEobOOGMkFYPnxst1ErlnbV8JYDQY89h2AjY1HEz2f
gRatcEZQaauJ1KWMJ7eiS/772BeET5Crt2oDEMfGMvmC6iLxV2RVc8G0OAxzapXkNpqu8B9hFZKx
sR+nP18SCm/296fZe2IZMm9BFs/u6UzYgFC3B0BrFH4JxnZ7LPTcGeDOpoYG6xlX/bUZ9ukuNZM0
nUpp99H8gBaSfYvuamocCZ9vm8CY4G9Vq+YVHMpFetLdtcSuwUB73I4PqZOJCR2gvI5tATZSgdfs
KWbrOBLOfzvZVQsUwagkN8z5egR71luxNdS+doo3nhFB0q8JaF82foU4S6B6c3IfA9YC0qWnt85F
qaddFkCS7SzDOqFmQrzf/NAl5CcoOvk3gcUO7x+PI6vaCquFykKjMEN7FGX7Qj/DQTEcC+aiqaOq
PQoi1VcetsfBBUHf3OfOga28a8eJ+3KNe69+lZzQOKQAsbYOEkSD2Xr3jBAxlW9teO+YMJche4Li
5osYsk70YF5rk9iU09D3qyw6kpvNohBJMRDci71CdYZhGzJXnQSR79u4V4j30+AQvsgpgUPrlNQW
U/DafZmc6HT1JcwMwonJx0Skm1TPI1dmXkO/BUPzMFPdb1zNYJpzLAz8yvUW10uO7/lMVNHC1aq5
MjdfWVV6s1z4Poo1NHfrT4g48MNqmvjWITk9tCUaPZQFMATyG7W57SSgPQiCs5eHcxkhoHlgVd/w
z9laCRTqeZttGnof2xkXZaQTDYqzSi1qK43YayysiHe8WKgMNubpU5QmzTR6PMPB876YVo/iPx+y
bekwNzWry2zhc1zgeOC8YezUENgWBQUqU11cwZTnqYKwxY/XcOegf6RHU3rkvmACsESXf5Nr8ILC
/qhJFCYwu7WkrfFw68droJfOa215wQrDJ49WB6IzddoV0vykXwTFgC7zLw/0bUkWtPKXp8XABdox
cCPn6xvCU4FISbiiwBiNAjLFWEH4lPmfx8Kg8EoiDTNGTl0yNdGnDZOcIOy8JrNfI4VFoAQnSPXR
61KZkRJkmeH44n6N/gl+BZngMtFfXjGYmvPq9k1MmvIkqARJd5LQgdEqTrjg8ZYG6fe+tW8JwIF2
NT38zsbEEn/67cnILyqPBNiK6reHyluLsRaNwi+bMyMB/rL3/vTTGxr/CLtLbVpxsnRpb5xdMOsN
zrxWHP+4yA6VPLGAcPAoScKHJ715vyZU6tS0EK0+j8htAOgMeywp0H0BRLzjRqoUc9/szDJC5jAz
alI4Tls8cbzRRNzgdXYS4pUgn9kwrNFEzXO4ZRywYd/IS34C+DQhEAzHIN7T7ncQbv8Vw6hdReW6
QF5WNVbX6rY68kWT7S3ugfSJrB4dicKLM6W7YhaD6X/MPTfI7FTyEfDcmzo6av7ZExtiMKawZ7oE
GGVFOzZK1LcgBt6hZU+GIanT4mHGcu6eJGdcC5NqXxtuz0xy1c2kYvM/uNJ9P5PDaGTMaunj/N2f
3/sQDEY7/X66/yO0N2YXZwEDRstDAzn0YWQSeN0evMov4OHevnSQjZ4p1T9+OSUh5lzturzwLE/v
0fmrkOCDAutHTVjNVJcJzbm2Zjx5Ot8CfeSmQnuEJtJKh6cHkvm0s0zmMYfcv5rvPmSVOSROiOCh
uCSQG4rrQtAT0gjMnZ9SzdEda2VNQMMwf2RTCigl1YY2bUoNXU7JRMV9uIrJyHkrERz/KgcxjmPn
DxEGlrz83B3to+rlMgGLpVTdzIs1R9c8dIqj0FL9MDNDXmyXdGAEFuQqq24EzcHemG0uDR9SF3FH
QYURy4drxPa0J0QdKYXeEBpD20IcZV7fxCqOkH0Vim4uZjZB/xWmTUXKnGxN5VIvgPMjBYC0N91c
Y859yPSfsYWPk01fGS/r2O+eawbIToh6+FuNc8CcJObyqcPCi+xDw3tyOdaXGb7dxOEv/IQxEQrf
RRFjKPzB+vwPbiq5zF1FdvdgfgZphVNxfdMmA58uaId5XgjAwI/bCbFcOcF45GWd3SDZ421Ill4v
H3Nwh7JT+dhox7DvPqnz7SRARP0oMl1evy9J72o5GXYeFHfuzPtlYGpL3GycBJIaGTsPUnx0CZsX
E96GEBi3v2LKk58LQf8PRk8X2cUogWjoRaK1bQ0g77Rb0OU8ezKu2wLyWuCoaE4z2U6gslquLxdf
f0PdL4YYa7yMeDnk55TCKIv2P3bDb5RruCLKPwtoefyFg2BN4xOnnxNoJN6+5CFmdRQyHWTNb6nS
aOAV7hkJtdgyP1y4DrtVXYqhWWfmDe3T/E24vp5V+NVuuoqAG5PqQc9yCUM2BM9v/rvz8/eaK6j7
fjnLRIMDjiZO10wVuNUo27L9sdnYYAf9AlDo5XiYotXT6gH+J9+jEdqC+ewNAX6b6fKRfyWSNvGs
FKvp5v6dtRxwpNUsNRrelNMxT1d2ZEmGiKkVEY/IHddsXKS4zv5pH9kVY9Qs4TpwW2Lrsu7r1uIo
WyOkOIv16LAWnLkRl2VY7h6RBeuobhQ6MeQfIecVSwhd5bQx0vF7v9VMFB7hVViQ+OwqWc846Epd
wGzsGYoBE+VZXTAMOrM6fJVFOX6raJR9hIWiyjXYT/AyIWVUPY9g9DpAenPTzRL+EWo30lUW8r5x
B6YZCJw/dJBewTBMwjMGBpMMDQnsqy3WmbijYKqincXIuCBJW2+NWtTvJSyX7hNnt/YrObFNMqAd
up8FJjQtjXhB7Gh24MhjakY9FNzMvlfYOGva2hdJxW2A3wW7JWTz3yHWM0r0SVTROKEDiHJSr95G
7n0umQBqIoi37GJxsfrdQlfWEJYz9hW2QnOwgZ4V91hPCNJqfh+JwAnTdU647qfaukuKXW6OmCIE
5hlPx91rt18OOMarysy1Z2kHd2f0aH56XJ3MNepXvIVxPuyyuFC+pbU6s8vcrzFar/sE3RUbBYQW
Ji69N+cMZoQdeqdYSExlR83BOwyKAF3Q2efeHvy8nde/u227ZNftMoK91k/dbtDZZDugtbNz4YBZ
dy8jOHUzr9M1GVuk6RBDrrPzTIE3WOihHTib0yrVNR1BEwF38TOGaHsQjbqQBT7tZEfN/DasGx+t
CjfpFEIOGEdwaAWffouSGuri8LyxdOVgOPDb8R+3oQ97gpCwZx3dwEvxdhx5nFL4HNd2PCtqcgbK
/Tn4oN5jFscWypVXb92k6oZzbatmDXQjaDvZoQsNhbglPfZ0i0nix7wMhUhjtVXKHV6xuoyWymOW
1QNWac24NxAgKj238A9jJXGoWw1ZHEQy8bSwJ0wgE9H1XKpq2/oewD32uAUhz4iv5se7fhi3W3l1
sWQwN7M1H38bzpxnAOiqvBMFfRyzbDEKIhuR3S1bZ69a2gIuSgqj9raGoOcjsTMzPatDp5xBK1f2
k9Bhy754hOcJ9jwFZVtLJFLQcqQZuh2eSSwqXTT0NSzFCSuP0bCDQ6EadhjtTj+dalL6shUMdn1V
/9N0RvRxtCWhCqXoN3+UU8aYv54+ew2/XVsuHxRRcgodNN3QWgih/g0l7edw8DCCP5E5TG/PU74W
X4PatKTtUT9wpd5I75nz9a0LbTGtkNTFNvWHY1+DFFj83N0NW1+xOxCScMkSCyJvOk0kg1mLflfL
cLS/3YQ042n4oyBSdbvuAjd+eMQcCsNlPR/LWJC80mpl7oRusMGNit8TabbkB5hRpLev9UJkNUOC
L4QAZB5JbbB8p51znS2itv//OVBH5ZO9vm5SvZcwNatyjq6kKgpPbPZ3p+X8GMIywBbxNTgOL6Tk
yAKB0asHpLJWdcxGsYRXQOc0hZ8dI2CIqugV99zmCPZTXtAnTdTdqnIhcYzP+qaMi6fV5yQnaYwH
cyp2dfaeLHK6mCL9L5IWfKTNDeyOc5fPzT/9NoE6yrGqIYKejcNa6Jisvpytj2PMC7jFYw8aHP+K
7FWID2doMLdSMTWYhQnb5DNmHo4tQeI16luICOrc792vQ0x5EnZ6fbNkhqSixQ7jRSqA0EKbsoIK
Almy+eQb5lMa2ADaMqMj4PnPfJ9FmLyA8NtlJC1MfmxQti7bZdjbaMt0gWaHAEbZG9YZA4UEcQE5
guN1rAM+8x5yGQAZ0tY8cucAcxKCg04E6sX4iYTiw3KwrCloOPEnx89H2LXI6o99KxIs2Sk55pdO
QfqySEji/+/p5lsbQ07zoZFEooneuQEkZio1H+AwjzUvvTkkvKG10RdTA0Tx8eI/7KWJ+3/GH1QD
usKRmrVav1455HNklazhx6cV5UFUFWldj+Ivf3oTZceGUGsPrBauIhhj8oSUECk9QiVsC2XrZOz0
gkaBblbyiVPrvWgjiqI7NgdufYi6Mxckg0KLnv9CV+24ZJxx8Vlt7bPuC/cg5kQvW++cHy6SqwMo
Z8PpFpQi5cRlhF6yCL0YU8ctiGxUOMdRfybp5IwqzLhsJVgo42oaJ/Iu1asRNBRoj0EIr0GajYDi
aV+YafzEmfqv0CIgos2+2jHJSqUdM1YGOTd1f4Zcec8aHk87AfV9e+9Tpum2ccGm24EV7zzMPEzi
yJadwOsrAmh8wob6nKGe1YT6ICCHhyg7yXM9ovCKn6/yyQVDIzImjXs0caAMT4cD09TkRpPIfSfe
HhcdVfsfIr5tAB9ilw0wFrji1oz9C/UdvOZB1tdDVO8xkRb2df+2P7IyBnPd/eYtJ36KH/2vcIxc
FVKonKsFzkPHVIvU4Y7ymwmAGQvy1saCYVqLFLQmjyf19bKywp9h51MU8krihyqtdcqxGeLL/3Q1
NAPfDqpKjLodsfJrASfeP/1C4mJBLaNh6GU5lnO+FL8JviKbswG2v3RD/NkWUQnGA1Z2r2WS97u3
FkCawKKFeXGnC4HYhNMIKjJVCl7Cy25ClNvs9nfA9FznVJ6ln7hPKOHiHulre5N6W1V6fDez0aU6
enIIcN0yt/F2/MJbV22SQWOPy1Im2VNKALkYMmVtUlyfLbScaCfy/9DJwFoaDNx1Q7pzRv6t0a+e
R9iItwtcSm96FlcwTjtokNb8NuuU9xHixP2RT1jxjy/4w3fEKNEadRSfnQKzgH5tndJG3waRCJck
HqZxZCVzLomzp1XDHyYMsTWkpew8peWF7fr2N81AeA4XxnQPhAtOhhD/MOWpSBY4GNkWmM2NUDvQ
UwuxrAtkzl2K1NP7uq84/bpK31WGERr24b9HddN5+DCQ5k8bTRGCGsr6Jpd/NZR4JjIDvrM3ZbiZ
cI0fN20Bg7/yhEVzQrxrzw5FhU+dfIToaIVnG1ZCKOzt8jcb18kWadq6Kt90eDzgRE/RvQEC/24W
sM70Fz9aDurXZn5EZsbxa1nSCVs5ln1rZ3TpKKkta8B5mSV7mI3qcGSOBrgGTCLbRR6Rz2JsH+v/
4+Ne714Ilfz4YBBFmQLsO+E5LvMZTn6G0YAhGR9ZtvxkY7SkePpyLUA8yWU430xhlk4Jd/9s0NHJ
rOMq4r29m6vbcODZbzDLFMnRfejbKCR8N1ixuf/rGq/4XlxHTfAAek7AOVycqIUe90VZcVbZxrLb
6lNVmCJeAQx/M27AqOrs6/8fMtSs/nHWdu9mIw4+Jn1dcEjERIHxVfdYYI0P0J9eITYs5uoYxAVf
jHMsJlpDkMS7iQAnBS1iID5CsC6q+RfMdbHxcLWjO/pn5er+H6aPpq3NM8UpaJY/tMl3S54qmaU0
qB13wNFRsa9tMZnn8g0oQzMNC0+jgJkN87IKUhX96xgrK6syw+HjVzMUevi3MvC/QIrH6nizqQ53
JsN1sI9t8FrrYk8iqDgYVseCViKN+sxuavvGW1UOqKYu5EZ7+1LQLlv2f9JD57ExxyQhASr2lFvM
oHFMa0QkVeUYWVkwGHNnNMbt/dAmGZbZyM24eCY7aCvwlSQ0AzaeTQHZQiaByUeDQ5z2CI7Uws40
BisGY1XJj/rnUinLbA+JB9wlteZkALIhJOVBjJOoaj/W/hlJgPtrmL2gMWN4HVJ0tV6bYEqIEO02
0nJG6LEGWZp0t3uQR8VYZkzjXdRfXKPAo3rHyL0Yy+KjoKrB2QQJE8VLvK9q6l/DmBFGeia+EKX6
7tic47ZAVV9VbTybCzIGHGeSu4oUQSD1ExUOam+uQoy+/6CINiWI/47dVNu9+4chyfAYtCKyvswt
12tHjeUqcxQIPmTF6AZDswl4csr11tA7pWsQ33OiYfRES3mLrvVyZkR3s78Lr7hw2vW7vgwAPnfw
aixa/saKaY8xjU9lE8Yy24sn1hNckLzPjR+5XOedSR/gq8SdxshPfVGJUdJPTJO7BgDZuWGgKnvr
T4zZvXMBBBACkA3OEo60qQdaMBkDOKrp/sCTXOdIZRsuHrqQEJ5cwERaIVgxzJjqh7hPkEuZyDX/
4D/HbiMl8Ada1SWcOD1JeMm4V7GOcs3YG5BODtN+uHAXULP2fyYXoCehsRokAqjXClezzb8/YWoV
xqiK5Bg3Iz+g5XxlncrLb2fjw6FC+IZUpaZ5Gd4KCQ6USzMowzE7tltd/Y1Zw+DnI9G8SOAqJvIz
mN78VymCQA8S946xhiHgEEy3NEH6stfX/Xed1t+7+JoVIqN+BlrmtJw9aiYuS7S1xZ4pbU/rTDOZ
BnPI4dxYf0mV2A9cy7xDok4cFO13Ux/oydocolrRodTZRlm3YRWY43l11MEj6gbwNlLQ42d7LNvB
7cG9QyRW0qnyo6+Pj+AkYVyRo3rEx+i1F57qxU6qM9FGM1FYGrGMccyKWGQuqY3umUFq6uoEDa0g
ICpXZlkAAGnF3Zs+4vRGbSC1EenEkwZT+VMJQSf8RWQsnpNb/MYIlYScz7f6w8D3/IBSP9Pituda
J9tkLzMsmy1uSihhdirh/DU3AQ2C/CiSwD635OL9OF3iie/frHqyHGAU16Uh+ZFHkfjDP86Kk4b8
vghAn6/AEkmq4NK6HkGry2qjM+iQAmji8AJFnc3t/G6j/noa7tRVGfxJytlKZAMilcdVy1bv6C+N
aFoHPcUnL/N31C0iY+8CEsM7CNb3OjDLdxIbE8timFN3iPR5phUXL0fFnjyIKbAxpooeSs3SYKuN
tM+TkbbFAL43jgXldV/oxPQOOBlSQh5wWJeyLib9kuEj4nW5v/7049RewzaabjeHiy9+TkMMd4pr
qTwXzdT105/RDJVOOh1i7wHcJ6M1lttwvz3xrONMNV/rNZPImgMDcHDlaznfIY7wbh7Cgt3mpN1p
at42inWNBFqBv4utpeA32jtci9UKq4dpt8ETH1+9ucNSI78Xxc/5AFc2bJYHrZzwSe7G1I6blXA5
AUjx9XzVv7xpHhpsA8vPwmCne9Ioy1u/u7FCjRG5o6jROYybgBsVDYsts8M97ukphJ5KH4nDaug8
nx8cU3EY0VjO+sR1WhbWVeaKcIprOyGoW9aRDDQa4nIXpKdniEAPCWuQ7q2nFD9YEXf9+a7QtJmJ
+orxnKC8wqfuaA42cMbtE8tlBvP4w4T8i7L85gDiLBBdTHHLAgprYy4Rm/fFMnKz1yQ9zGgpKoz9
dEhdb753Gpti71ZWw5/LBPdlqN+W/q4mVl1acoXrNiOXr7bHQacs8v0WrIgyFklQeulfLHS2qwMi
slfOEw7LN3HxLE5t7Sn9rrbue0UmLrmd9jjiB/JRB1aM5PbBzmclzLzkLLRQUPhqGhhzNoS2acI0
q6jnGIAzBblwe15P4HOD/bPpbOr1CJ66ErCdsSmuiGwZ8RbZIcxZLHogFyegPv9WplhtoAateuUm
6PZxFVqsDRd4urYi9jQCIKhs+6XvyDb3Z7T4XAQAOay/jRTnzFSd1/ud7ve0hXN++7+qUjueCAaR
MfqrVC7RIaxAc9n06YAYysOoiHD/kLg9Qg4nqq95TNdrlzzpIG8CGQWRm1z3Wy/qrd3EMYMT+Gbi
FhliTyJUvWy/zDlspPQWmqKpax0AgtfuCJwiP3c5q2HRedfHGIDOV9zJZPyXnzM/8TK+Xv+99GI/
QufYoFgAuigLMtQ2+SwxwOpmUl85jtOv6BLyH0szqihS/a6z2c+133RqB8xSEPL5PacswO80qbUK
EhjTcOMH7F5RYaPwzMbeXvZ/Tk9bfbYENVui4ndpC34Q0I0YDzVcTZkntVhl8wmK6VL3iVN/pQSY
JLJuYCYDnFifzzC9kZ8Ltok421Hl6LLn1uVM0EU3Oszto+/l6l8r5J5jVcZAn46/8DwBPAoo1UlH
DQM4ETviS101bj9sA+kcwOb1H9hMQe3qYPkfzjyITS681K7O7kLeH1z8CwXVwXvmuN3wXz2/ZuYP
I0kKH+zMvSMdzDEvNHqknpND4sLPHw3RjFnO3k3EBdde+74L9Jd3G623hfLhVc7r03RyqAgB05pt
KS0dpFn37h5Eq6o1H5iNhtpPxK+ipxEzFcJLzLuqtYhArNX03nza5S1Uq39tdB/f2CLuwttQt1ms
sbvAPoilERl29V4cVppTMYo2EVTCX+CilOjDRZT+DUWDprLLLYC4JObCRLVi2rZorAVaQPcIlQPc
8/WdGt+dYf5v1FF/eV49GEZjjuI1dTpMpzXJOOzH8OxqnEkDRs2DK9PblecrpgvVI4SHDVJ8iwTk
++j2IGBQ9Wk3KwEjbsSVKf9rzHDfLLFdB+xWjmKNS+OsArbhXhtShNfIHB+YbpqKwmo4t/Ya2AGT
V2mNehzuviPiXKRgXNiJsIJFaheBt4BUVfYk/RPNkkpSzLP2RVoKOmWAzhWGekoMpzAHHz5Htbbf
m8qJqFxZ0m78ZA6/ByvyEN7Fvk+QsQPvWOOOWPOw/yuVyEbaAXDulpykcrIfl9Yjp1syMwbAYpZG
QF7av4DC8FF9o6AP0QOvkN8Dx00IgO5DUtKXOEZGVescA4ITlBErrwyRQ9fvOZIt70snF5NA6yay
KIFot2JlWC3e+T4gFl5K5bgBFzg8ojZxgDYlPJ6cP94X4iOBntrTJm66LoTMYNHH/s5WZVM/l4A4
Z+1H8NlGTw9FMy8J6MkMfkvreAaqp4tO7IAdUhHwNHUNQjXxID0IO0PtiWnCS12yCdkrKQmFA6Te
scO86WsCos1Q3RgSbugoVdCTNCuczFLWkprwzyATE2tDotvyO8N3Wm0wV9hu9v2J6aBzG8udSNQg
dgT3qBcLxOvN6zRrZ5vbGRjo8EdIJAPDwg/2MwgY79c9btVYJF7PQVZIx1rqmaQ5mdXSlZsejEm6
u3/BozcdSJkgG9fM6tsOFO1QPG1n6fJMVgkGFjjxG9UuPw+LxhGEha26wVlWWhjVpidV3+EkuOBX
NQeEfe1kipTmuie04TvDFF2qxyFHirArC++rx2cBJUKw0F0uswLdXuycduMIS6zB9PUOxZj9mUO5
ANBGnhhLGvDO4eKoBkAknIywmmDHwKDdMhmj5+ckVNlQXS7YXTLUVKf1W9RRFrQcTOAG9I58I1ww
9uQ8xAM3wD+Zo9F1RqaxHvagmPmYRr0op/5g58rXSgI0Hj3J1MDz/C2zp6uX34euW82fRwDFfV1b
YvdVG3ZFMeTb5YwucZaQuHK1w17RypwP8Fec5N/zy/WexVkuE0yD2kjaHiZGubBMCOsTWfZuUwvy
lSbghBxGf/swnfVZl4Piv773aumy6pI63dhaXpi7HZZX+PaniYI1zCrtgctq/FcN3ZZetVdfbQYu
QDRjSYcmHq+LT1dCpneShhvyo4hO+QooliZdjhvVfOXRqQm1RuL8uip55JUo7Ot5HooOdkTiYBLU
huLa9QLXNZ25tv5a+8PkVl4/uqM5AE+DRvMj1q3kx93X1tVigmCO1OfeZKTAi1VKaNaVYEDcKcI6
eXt99cw6KIYP2PbrQBlTRLd0LJsQbjan/hmKqoLqpeuObxnlZzuDsP5IyH6oyTitPRE4B9lymhf9
V1yGU/mNdk8c0ZwkoWBJfXru33dAKtwI/MJNna8Gxfaf7k/Mm5gXQgPKoBDnVsMzzc3aJv3K6CTd
sQlqu7ePkXUGGKeoTFjdPE2OOmu3i8JMjBkzVdOc5JYwWY9OMBXRRdkCEp/59N1ibgpV6uYHQVv5
BPLZwQd10WD/MQ5zWfqlZi/T7sRFYgiztQHQ+KeHSYi9nYSf40eJzS70laLXgUJ+EncNWYF1DlNK
kUFrZ8sN4CKc74WWhhYU+Al0IQ9NBd2hp1sNpo3evn1s+IRQu6RtOygo1CsREBZKlte8rqIjyKBU
NHSvb8Nvfg9XvyedP3E5LlMLm4l7sAQEoQ+v48lBi84us9kBN7refskebyPQzsFCf/DeivjyaO+6
3RsgdA+uu3Ti5/3SWHmAlj0lgjESPqCXO7gI/V4UEQhrbd9Eyl5U3g6rV24W3ntinLMgFWhiOvhM
YrFZEPRoSSGBXx2ZqI2uOZrRbo7VePLePdePALUbcDzQKob8gKJHbLIWuSsfoQ6gjAO1AvPdUYOY
40QpN2MdevbEECw1bMgaQuSNvgSGh7BmpHCj+3V+FM+B+PM/8MPe0rdhs39BDBrAo2oCJciFasVh
SQovDtXvmaba3p/aL9uZ6TFnyxWPb76IFx5Ly4U63b+/25XIaQ+IIN46lOu08CBW4uIW0zLngaBb
PqoQOaYYwm8OF+lipr4YmAoQ16uL3U0td7FPc5AWSYLPEypkDtQ5ojKucoPLDCmoNmI96rqoNpnM
sd7e2cnLDIPVRBBzw5z8s95/yAgcc2nCm28iQH5IEGAYs3nXbdZVE8x9shQv50QmpyjV9YWj/1u2
8oeHlh6q9JOyrbOpCdOhhVC39JbY3w88Jd0MEk9dJlHIP9UxLZESy7SNHUHMmMIhlbKJBmDouu9Q
V5vGnoWsigK0XfUc8WlS5koU5Mvw5WHTmhwCocaUhrhYDHb+ZhRL7AXcFTySrcpdBAWyZwFM54E7
y4bxPi+ggcOrQ51d/MnCIGV9ZkiciwdU8Y49nNhGvAual+K8dqk6stAPm8LeaqyoxhLowNrdRT7V
6N1116caVj9awBnYfQZ2+v3c3spnjkjrUx2lg7t2emfIRkp6kNpDg2tcZYCXGzgshZ8mESry50CW
RZHgmz8DlSSglDDEu+O4ojR26NHmY3yyp5gN3ecbiOQ8L+hSkYG4A43zjtqi5o8+7bvHoe4EbWbq
cH2/1m3ga8EfrCUSHLtQd/hrLHrSzbn7v97YRFLeAkG2h9BVvKmKm3HDWXxzgyA3FwMmTmJ6Ohfr
YuKgJ6/o4OyniZvosQ61mWbtvZOfeMJKIo3/I4545CRD+ZV7OiyTL64wfFObu1WkGxasq5FtoFvc
ISoUKeTMHawrgd/le41DuuX6Uyd/3wrzwxK//JajpmaUYwqEnSEainPD+cU8k6Fq/fpBvjnHTja1
3EgIeCUktu2CxCh7owSpua2teOwFuv6KipW4QtcqaLDH+FB36lM9aUUheG+S4tD7QyV5CI8mSQc/
QytmFgYzaqciJSgNobCZBB0V0T38Lq1uAged2i/+oHyULABdyvDukpjw7Q1jQFUQTUhABUpAAM6F
AnaSB1rT8iwCJoFzGpBwLzY5pW7CwdIVD1h/SqBDwxRM4hA9GTzlPkAwIsF711XgAUNyX7bBI0IL
Zj+KRiRPQa+TCmZCvUmDpwpyddvr2QN92UI1D4sW/dnjz76HU9cj/VEp61p1fb3GTsrMatGO+ut5
EplxcPpUyZyO69SoD4BGmIoIBCeTRlKqIM466xFbYdPuPh3hLr0vMR5zZIleJ+Mv41j7eMDHmyoZ
zon4ua69Mf2BsJ658yJZ0xAidF6pYEvKeF5+lJg1ewmQ4t8/q/xJ6MFnhbcydaDJ8lqt6Lo2TfcV
mklrcBsGUOx8J+xfg0XeTvUz+E9KmVj8MX/5esT2592EpyEx3tsPcGKZdfZBSzCTW4t6KX0l8Xpi
xG/XzeM4JXyYAq+dWvqZS/VTyKdA2wx8sAMdl4tWKeBbj7FX+XwknfUlSG6TWItJu8SIZDD5YyiR
vBKSwrQWx7FTpUAhcB3EsUz2VgBhny+PuHD1daNA38xuuL7M+PORvIb2ql3zInnNSk9UHZ3x62R5
yo/04eIyTGlhgLbaZ3yADdk1BdqYVA9o4OvL2H91b6Iox/SXZpLmYM/Uy+TXwr8mg9xMGC2RCRqy
zs57pt0ERtdrGWYpGPPlUAY3f5zREUYw5ajCOgq6eMPez3xvPHjdi4XrfFtJ4mxxxC2Wh+84cnxw
HXKojfNWvg/7Pm8JjMUE0vj6ZRlyYpy94FN5Xg/oquBA4+B4XnbhXc4r4qCjX21Q2NoL9bDej/kg
hsrdO0e/3iuCRzdjmsWKgQv9pUloA4giPZIYFRVBxGYTeBXF0o+5piL2BmV4Vo8o58seoJR1V0ZC
G7c0N2vGyD91xVONTtbuJ+VlXAfH66Powm43scbYp4Q6bCGp9iVTUJsDR5JdmzUgihWedEySXCS9
uSo/jbkFRuuwpciTQGzeOErdDFDKrE62+C9sDkUDMySuLhL/ANsuKvzIzWK/h7FFDuGE0rmdEPNM
qCMlyPXcVgXqJ3EfTIswpPqzfSzh7ON3REMuEbwM5vJqIcqE8oTWYgKKrZPzFv7ypOyRzE0eEl+G
gUfXdJe1KxS6j9lVSF+l2A2ARqvT7aLAHNv1oVfFkGR+A4MBgvBhydTkyfDNXdm7Q2rFUpkfsGhl
h1VwB3sAwOcQNa2qxP4DeCAzz0f1y1rQFfp0u8CUScpksuWhzFy4rTlrbpjILbWpv6BwozPc6Lpf
mojoEHhQ8EdERoetvV//v6MRz6ycYeK3Dr+c07acXYVj4P9GJXQYD3vllJuQio6MDeVKMp27Cwiy
01H3Gf6trBs4L6I/oTXG+BmSGhAQCJeY+UlAeiBaqa4fNNbXg4SGWKbfylknQZMfIogq6hDaoqC+
4hpmgUyR0PBhB6R+bswQSbArSbm3XfQ4eweiwG7FCgEp/rIcT0ikQvIGks/YpemS+/ScbNkc4LCd
KkTfXLisubGJzCSHiYm3UYS0lv7q5R4Up0YpR8DtMO0FmM8ciEIwvhk+mrEzMszdUBYHOQNgvEWt
9v66A8z1VooPMPHZDK5njQSogUjH+q5CU69KsVuBESlXgGriX16/rYCt4SZPQDwkbUsr017YveCJ
pP2wbq1R2AIOItf+nbsFqMtJw5a+mtqEbsU5FIKGZbhfEFtgcPGd9rAS3cg39wUT07++xKzBWimW
Czt33+T79wD4KoPA0rfsLnboWDzaRKRBN5HBNDUIP8+Iz+sNo+f3ArrJJET7OkcM1vPD7YxjaVfw
em9H3e2J2dZJd4XASenaIZ7XRac41l0huU92KIPbaMa51s4r6wVmquKXtiki+n0D6Ogoy/O+XlmH
pG66L5JzXdwFXhYYAQ1hNjBY/r7tTDtBOVMV6oVpPkAJGNgvb3k0jzWxxYyvWOaCbQFG4o5btwan
ui6/RdC0MWevxQXFphNJvU/S907aCfGFGfYKYO6oVGSyi320VfCjSv17qv1adeXwvvI1dZKSYuXQ
oLF6Tf4gONdgjBUBeQ9X3/HSBW/UQAUuVi11K6ewArW91IKBSVb8xqke+veYIyD88+/F9iIx1WyA
cOMeDw0JpD3TrIC1Mr3wELXmXkKfwOvb1ql7Z7BGD0a/3witnVt1OJFNVc9n45Yrv+7DD/XjFu3r
iu+GfTtKt85UDf2bsfsb/zsJqBWTgtRcs4VltwsSkNtRyM6ybYZPb7w+NshOgta8SYroBgqLTZNz
9Kql0SwSYCdXQGJLGLml+y7kyWraWBxQvofD5JzZ6+1tr8tNbTT/vEmbQZoVY2qb0JVopbCOziY1
5WodA2xqtErc23DVZlMcobxVn7jZvN6YVsQiGoEqQNqBKbrDKx9eC744+okrmFrUHOazZJM0bRQG
VCVlu0wbHkNPpy5TWQVhV8nxwR1Htpp1Ux/Jll+1MpfJ5fEdzEF9H7NiqRKePIBTEee3MrADVZcf
hnMHq2jC35DNbGmP7UqY+88WO9jG/bPggWsT2WEFRj6xFJVn+i7dCk4gj1rVb508BiO3npzaZXbA
c/ZRrjS2zLiY5uxONILADyqPZVDdjinRXxrN/Dxz/HOU9LxlMWbF4cRMkp+S+X9rhqNNgOu2atUy
yqXKiDNpY0TDAtOM1B9VunspPFqJWdCu+u4X78l/x4pYTUZ3pXomeSe8s3320P39bESqy7Gj73y9
D8Rm0d+qQcjvxy/1aHIHTRqj71AKRWrbrkGVwm0BUr+sVfcOaOoCknGaNO5qJAQocFZmTlv6CBh6
KGlyAVWovl+LXgu0ipbWvVsqc9F/rCVmRCHn775KVaWDVIEHaKKkHUgjs9qJ80ZZzsVnUuzKPVo9
0qLwNZ9G/YL31fabCSLvow7nYhCJzHjIv8JFxPeZENzOortRygTV6sB+gZXy4y5CjFR5EnOOocYE
SVJz0uzPsi11RI6Y37kRL53loMRki5akkRxizmxHboP6a1mZQ5xfpt4t5Hgc43AtovRceb5+thvu
9A94Uz5WkcrPBIV7cgbps6YajNinqSles8aguG+RRG7gazTblFaOY8LxPQbotwTmN6rPpWEisqdk
AByVCCTdhg9JfDCSJPsQlZV1B3YGjsZsUVEm+TQuvskmhVA4rO8zqX+FmCKmnWEBY3QDb386IU3Q
dxNQdhV71j5B7ckUyC1KaR329o7yeyJvvjnRj98T7XTxpXPHfay6sMWlwB/bBUBjR+w/+kzxvomQ
JQ7Wz2kI/zCAgFh4gRPVexDDKh2/Oc+3YI9ZlUe6uV66WSNeIWIUqUdMWN6BzcjF+/yuJgVMgDoa
B3PJlSfdKxsxjWhdV+2cJ5s8Yyvw/hE+bTaPAN3tQ/bUXpYT2IRLoQHlwzcvdM7OybUWpg8j1vXq
bN4ZoLEl5kbmzMTAfpXuth4ZwiRXC3uQjtCP14bUGbjqEh8ZTMn0DU/JC2OwIIZrGvukxhTqVGOB
L/jTOZExseI5LHojHqONtSvkX4Q/s/jMarvHXUNqe1Eq+gYUIiWBKWe2/dOzNnOFclEa1jZS+nua
Gpr8FVBteucncm38frRFTwGCh+uDSzGie54vru+5U2yKinoBEADQcsWc6mWkDjoNkJmR8X+vub6/
FB3rugoZnAsbm8GT3K3tTd7DgBs4tlDEnHUThvxyfB9TtJXpEClYG5ut5VrdG0H/KI/zRyeSlt/r
POv4CyITjha1o3VXHG8KidkdKYjliEOzRnGGYEGE/X2XIaVciHzQWdOtDV158C0vTnDgkh7tIIsX
tV7qYEyFJoHrXifNHFSch7GEC/deXEXQdawGe8iVv+l+Hux9A/hOgwf+YQLAxtmhYa1Ad5YzBq9t
tHaCz4mOuDUZ5CNjzoJIgLXrJDMb6paoss0SYSH1conz0CrzPqq0FMG/Zk+y2tHRK6BztaJvUVUt
oyv2D7oTmQ7KGfG6kSWATjf/KOz0mzmG9stt7uyTzYKrc0ZP1MA6+rLepoQoYtL/lYonmW5isaYF
n+Fztk1iFYSwBn2YlVC/ucqtWpMgrGpu2xMld9eYjbxLvckP/TS7bjubQCUd28GcO0N3h4NFBo37
jrt7Y3rbSKBOjIjNngZiDvQg/HoBHWzCAgK2xmOCW+lk3RHx+VyyMm/MIyAFnQfcReZD3yMZpIYA
qZ+wADrv0H40WkIJxZsZHHCfhEjta1O/utiIUK824rKB2oViA++fLwHz5IHt1fZs5zPMmhC2zNbr
7F9pq96UmApW8F7wl1IhhDPvUPFwn0SHILImfiyqbumgnYhSEMZPv66drm68f2oerOLGmcq8tyDh
Kav+A2G8YGetcQBbu4ekdJVNg0o1mKZOw1hTPmXSFm8TvghoMzO9qWQcvfFujrD/bRcWSODxhTvz
JGxPdqu3wMclIUIcprXxf4/55e1o8h3Xc+4BTwUkMd3fIdQpKU6A6wwqHCqKUN0CO9LE2bwIUKuA
oRiH5EylwCnQ0RnmOCH7EuD+PBJNc5w2FefqcPlTBwu8Terl3ACthJ+iSrmK92fhUecwiVFs7cwB
Mc4okFMnKO6HaXEuZRvw9BfSP11a951qCb1ZoTDVOUZt/3xWWssNuX2hs4jP2ijBXvvOYrRZLMLH
XIXRtvsdM69GPDOkxPqjV73JilY7lHr9eeuEup4VeKc0s6N5olNpdbjVDyi+gzdf5ATJ+kZZhCui
pat9yH9FPipNDc/oR/psqicfySRqXZT1p0+p87pY1YKroonAoPENDN0wOCYeGlleOcT6LOKZ2Zqr
Fwn4ViAqZ7/btDV4RpKMuflK8CG+DVjBT149wjekkyXIxmlY7vxAlLUXj+LSO/24kHHGtE+RzB61
NGkWZsuwF5hMPksYOL53O6bQmoG33RqHnH4oKWH//SZapru8RzDqF9WERrgsmUR2en2dYTqaHhYI
4x9zU00X4kVZ8Wbw9265ZD3NXwWbaAdpVCF6QaJMv1oajUZOw9b1hMQbANPioZS8xR43VgnTpozK
hqNXOFmdAX//CtgUUSjrjizd5gJ5HuTLR8fWxxLPpPAFAY8lnTZ54OwPpSVR+W9sRIiAYsQhVUqA
XdKdiT2G8yP9peq+gzKlAUoCSzDblyTFsAJxITLZKHmxnirOlt1987xs0lT8Atnf1bIQLiZCAQCJ
ady3leboQ0B0umi+H74IoEAprou7kYHpkMeunSFh3bUwcCPtUdi4FvWqq88OpzwUCTO6LVeVFVhX
+DSPLEH26pq2INqOCWG4B/XILlV3Tu+QnFNEK17H5ELuHBG5PzcIZj6RqiqjKfdppxe4R8be4RE4
jpwNEpqtCYWSluuG/XGqsUs0HFlw7XAcnbCkDWWHsJapX9hp0Go159ROX1kMsmhjMmMuwGvgrRhl
NrC/xaRN0ITGE4uQPiN+FYd0GjKEr2tdMue+zBb7htY/3HqI/omm9GfC6GcHkw5HUsbbgbQ1+8SR
9VVT99ksvKmHbHrR8dlEykoiORwMhe+v+ifVMGwkdjYzpY9Sie8koO3uB9cy7JsE/Pvs4H8o30C9
TcEHwpzcEgLmlU9n6pDKIgoRoDWKD4/ta6isxxrC/QkSuafwjQG8xod6ZVKvJa2gaOo7quMhH23t
CSnuBWjH1dfiPm2bHtlFLGWp0xl/cEsZ3etvQI2B7lXZJQVugS/XWDjkGTqToRS30BXtG9s1B26i
Ek9JpfTrY9rlIUTfiifkXrN9B9fEH76upT90d/ZFiN1MUAvsSsqkU44TGEAkK00Qh9vhm6EgtT3L
oErQ1AiOv8Keb1C2g3YSO6nVeoOxQPokxsevKpkO38N+ZEbMcb24xaBJA7W5kgVylrOCvJuaW9Z0
mTDdMa0HpBWDArSrsfdySlFcKb+ON+gbW0dQzaeDgmTeh7uuz46UiVDVYbpT92bYVkyy9WWPBPmI
upcdRmV3BxY69ZLzCD3aYFKkCa/LW/XPZupyF9qlZDTxCppudOOKWVOVVNRLBLGRz1iP5eZK0uCU
RF/Ul8HRmO/5OGKJ9zjg9Ih6uqnKSjVOcqxMMbn4PEOZXarJRiOYTgeo+R87AHG/NEBeuBYbFE6o
/CF4t49cjnT9cVaTzMdMWiutnkV74t6HkYhR6d7puZ6CCA3g2h8FJig1WZ0BhnRAKWZUvTiH3Ta8
0vlQhSghlHpwMD2w+IcuRxgevpKe2lY3fnu5ZZztga2rXEju+wBCGwZ3RIDUP4L8vu3/izY+q1Pf
0HCdVGewLWo6+OkOdQrTm78k89kOFdWbqPCERT/jTII6UTWel8IMZTva7JI5TByFTDKjCUe4m4Td
v65T916GHRWK2bd/6kHMkLx42LT5IMQ5fXoC5egKCeAi4EHCTBnqkSEBDm+rbVIgl4sGz2zhlZem
wlEY7ZMCFamox3ocKcM01i79yZdk08riLasfa2c7Rj5Jplh1CSfpDWuw6tP4jjptTDCdgl328hXi
7RjF2BkIhUaMDi79vYUr8PY0sNIEWon3mZpueEy1z4Sc9dAm56JOFiYdxDcn1uzKunby5D8hIKiG
PZ2BSNMB1X5TsHZsJj0/Eo/l3+hyYKJe/NaIQkUvaKNyti1xTJ9uyVNw2PwzWR3rYnOJsZN//+3J
Q42WNeSdqHRBJWbYwubW2OIzwMPqr4s4tTu4glMTnwTtlduaiFxqTlMPi8ZC3hZsMfkZIbpVGDFQ
eZ2TWvslGUuSGX22s8RhbAJYX/hIhdclwoDbZhE92hdSV8UYp3ScF5MAXxJksySSZpMgQeufvpX/
PqHh6V58iZfTmqJbYPhVevsenQlTcyja+BoxQwgd6x0AHSz67BswlzG+dt/DpG6xRDmfwx8tkcfL
yMudMsTrJoChTlHkpsvqfAGkYQ8ulhOy8UL/dzDLEJHojSr7lG2DghBbqbfje4JUPGNlVM00ohEL
oDIGNbZk3SjJ2eT0ggMe9BnXQ8tUJA+CoXGVrBwiQ/DKMD4oXmYlnbq/6iaSpSEfqTolzwe9uo6A
4cdBy2Bbt8GJVcXP03eFNNhGchElss8iJsrd4fpc4zSUlrirMSXRcWGjd5uygfhk2gk0DsRW7JW8
8jGH/bK+tnTTy4AbjAgcpwfKQ0ZdPtYHs7LMa3oi6XcRqc+3YpeBcZKuEsni3LUKh0E6bN2ongpH
KBgqIsFxFvcvOG11zUuyGlTUTyw89vc+2W6j4/12CXuzl6O4T9bi5j/gP5pXghIanb8uhVYhlWAm
Twh136IVqB9Tee6XcakZHKv/VZV8N+oFScfkyl0pBtW/Wqgxq00CyqXZKgj9RhDu2TeK3vMpL5sf
RL4Tv5HbscdqxFOchpDfA6Ns/QkjrLIdSHhczJhnHXXipjSpuCS7NINrfroR6hXCT2fH6IEFLr65
tNjW2catHvs9b+aG6Ct11maYr/clbvcXkoDSb9zRNb4IUedcX6mJc2do24e2M3zR6lqzg1X8HAiF
lmxfCvMBXuktxZM0RO5Gt0ZVHvSXvNdKjNm1NGLOb05Qu8S3BcheQQqQZiU4xjsIzX1GcRoVIIN7
onCQV3gh29o5PVOe3zIUg2GrLKwkwOuiZZEfDWaVAJCg5oP2Qh+SsSTwNhKq0OSQMlkqaESlK76k
A+5mQYIj3FjA2SRhhpdR5/VcA5AcbQHE2+am1907pnprZi2bObCtetypW66mobWBIlOeetRvChjK
pclqZrhfNBi2SKX80leZoe8WPV9pQW0gMjj6Is2Fk02ACgwGjT8FHsHFWJHiV4jpiGGTFi4crFgs
1m9Sitk6lYq6J5HG7B4NgBOnZIx2APTJ0qoH/GnU3JbqiB+hBS9J+zL6LcVBVvG0wWHDTDsB8BYb
9yZe+y9twiR9otgS/V+4NTNJGbwvfvEiUYfWVCsZghvZZAeZNL5R4YWL4Alh7qC6+ZwiCJiLHCR9
6bzUmRrVyuFnDFLKzYp4YERVnRCJ8IxTb/o6UhZ0gPl6fTeA2JoJqZsyyU6XnfWGXrQAsbQwaKE8
1F/zduFe/nYKtz5gVs2He9v5HrzlgQbaeb9vKJUqjK0EEJ2j22FegMtaY4GQRnAcMCWwuJTjpOpP
NR4BinX3zVAzZDTNsHiUYdE1Izw4dqYg9H7QTT8xz+05+RJYr9+rCWMYeDjhmlafKF4DdAOv9W8v
1BO51eMg1vNn5HoSnNmEFSLhUulOn2Vvbz5a3NfW9iBJQ14JICjmefV459KUdjbfeAsfydvAbAFC
1Z7ksnc3gpu9Z6Veuqz6YCJsgtvnGBPCk3QPeIvB53Kou+LdMRd6MPmgQHv1yIAukeZ0PdDWvit+
0WEfm1Ciy7lXd2/WiVdIWy24KjvP7tb6QVPGSGtEspGK8o8tY9T1wIUyapGSsllXGyX9JOe6F8yi
/rDGaWzb9/pw32JsVAe7eC4Tq1RBaW9xfnzEmotI5QveVop0DuJ8nALzjCdPPzsmhNn0DIt54FYr
XXFDd9cWyEbkQ/Z0eX4XxetyNMT/ulI+JG+lcofmLPLzv6mC7KktKH5XFY4ARKXnnGxOmJYc4YGV
9TflPMjjoMJXz7Qnbt29hZEmj6fXhhlzJlESGDqvFVPAY/kCFsnDQcqKUYUNAbrxH9hHZuMEyhsb
Jw/g0H+sOTb6aTzF6iBlxLZ5f9KbV0BL5wyLfFfyqIYtTtrwcwi3jnOahTzY0e3A/bBMCaOUiYFT
qdXrBGgrWp08khJVpiL+ULGXBBHtPIB4RIbukdDZU4Dl5q3SmMYCDEFSSQ0rzObl7rVmbDuMay0T
Jbzr2lNXVu/gZnuOdY9zqpbPzkkuzBpswO5FumQE9rzl/ahl/Ox+nqkUedQBFMiAuj++Q5he87A9
4AmpwEPGyLDrFpU7wui2et1UhOU/ptXutoAednufyOv/GmDocsZT1l8BhWKJe0Xp7BhGn/QV3iM1
qbVDZxzH4juZan/wnc1i4ECFgl5T5kIzPYW/HOxcXE+mMHDxqyN6x/+qU1hK9kQeiR1yr5bydU5V
Gkv8Rfxdl1IL5jUI/kz00zPTGX1QaVwOOie2k33I0AmWdmZEc8Q1931Le1203ivtk6AxMJa4FNLr
kM6oOmCATRnB1tpVzmfXCetSZUIwRQ4vB+5h/fl0PMcSQqmOm6YXhDgGyGj4trK/7Hg62cLgbT7f
JsRe1t/XcAh2OzrUclERIKHVJiWD7sGaLzvODEQIHBLfJwj8UYRK/oxfSn8ZjBoHeixLZJBXf/0v
3JxYfQr2zHCpYyfHneSXEhKx7U1u/ahKz+4FXkKrP5O49EJsN2SC8ZUX4m+b3o0pqsT8WC5Oymel
h07/DINM0J+7/N1omMJuU7TiVnACd0Z21Ad1v+8pS9hWldYjdYCWmz7rzKOUTs+8Hol0XCZZ6QYn
g/xol0XnZdctfZ1GUGiYslpYanwz+y4G4InJZaf8NiZF/crpktmvmPcN3Sxdf6lxigcbR8G03cp5
QCq8RpFoTWBTGNQXotvip6PjbVhX1W+7k0z5bh9CpIWcidkqdCkCT/qNYQSTVIPXFqkBlmidiA3W
s0+Bpbn21b1JTFDittfqE0FxkdsQdYT6JA3GuOhffwhiKzhD1K88G1rsfhSLflold6cETRfuuMqT
MzSCfVTF95xWhcS+ZAodrKssybfuBDAeSQ0my7hi3hS8zf7acdhrCK8hd2UqwXRkjt/puSrsaFIY
DGwaQXjnQfZ+UpSXlELS7CeqW0k1soJseYBSzHwMawkdZq5Haf9PeL/lBLOqZQrmhY59S3E/C4tI
2kyFbuY9qIcDL+OZEkvtNNaLK9UrItYULvZy14tHQbPI/BI2rELKQU7DGXubRC+OFGzw3IRH8baq
/MP5++JTL9QQPIFcoKwgkWwp9BMzLdIPhGS8btTD6x9ijJ2Zy4UR97NtkkWw2XxgYpm4LztnuDWq
1D+Yc7kH0TStg9GxGQR8uYfL25gL3EWxhEVe2d1fjoQk5F/wSLAoTYeFrtol08CGQ/oPv2Jr7T8O
XQcCOIaFDUVnVs/Fw9lYs8i7tD4aTNA8nPPJh1LGbh+lWckyfYDkilasmHaZgbxybrI8+1Py1QQ2
3AN7Qwn0V1hBq2YBj6LD/JAPXQzGYMwy+/ETNIPkLirHMjAQ40Ld4gsrQMOx8Mx5MJ8gga5isH97
Mv4raYqNGWvE3UYAlHA79bPogDMb/a77u8kYwMjNuuE24lRstUHyCp9hvhro0ip/XL7TCInYPIa5
6T3KgKamnOWgMlq99DvuCsbh/yWpNPq9tYbzlcVNzMAM/mHc3Wc2IjgfnXTjZII3Rhi+ynonDbtR
TschjS1Q8iM66GqYmiSDc/gAv/GtKvcGFQ5DpAsBq3KqDkAMB8+2W9hB02qEXQFt1uCXkBlTZa8+
jUV3MEq1ojX7ISmB9UvwvsU0oEq7JcCHWqs37fteav2pEUasP++bPeDUhF8SKfakJXQJMZ5jBv5R
ghpwxGtjwTL5II1rARjVCkzxJHjVCoC7hKHEF688rf4jCDZ8KehXYp2b9eG9ufv9fAe1X8KR8AbF
teQIekJC/N3t6pMz8fJjVsThsLzssJVTxUgk6BYXaZy5uYxjTLBUk03QL4T1w9fLTqcM1riTvmcf
vObB9IGFrib3AOdTwWaMqRQBhO7BQKVHP4DiFNDtqiHU0MAOXXwD7h0CLCya+1KBIrPs9pcnbTMj
yVhWcQRD+QAfQPv+tL80/Sc8gOcoFAehUYpiUBKZhvrrtMZHK8rAVpv6ZR9mPM5xoAp7OSHruGK8
pzOSk6ilyS9R2v6snlhpI99OVcPIKXrDagNTSaWRlzCnakndRZHua1ChdjTqegK2oHEROYG8pq7f
KiildGGsgiWsJtp7Map3shNt7YhVc0v0qExLVh47NvtPy+R4y7KlgS5rlYFewhNnMj8DyQck1HpF
VNGQqEnwGeMLhrbNvvwmJzM7lZNcX3+lh2ANt1xRHbHI0eLBjnPmdqv3nmxJH5uSxw32/50aFSwB
yNzzOPEftVtLTkn6pZELi8sOO2/HjdlVMDkmaJXzDY+vuhdo6PijHgMI1DOfMSuqWxayFA20Lzho
r/HsvAAt9auOD1Kf0fNTqZnDxH7GXhw+w1I813IW1oLET9eyDE2zL4HqdGXfYAkYHlcG++oJjkRQ
CzhEaKB49IW17Hsm/9C3JuGeycSqMoCgvkELRHAN6AzpTZXryTtUFCWBvllsjjmIuHAdf/SRoYSj
oMTFLlGlI/ykcgLOSpxl/09wwaJv+w+s5geH5en9j+Sv01p+NaWZagpgqP/jVBueBbgtXa34p+bq
zWCTIUk0LddoDhuE0Njlig7bexa8AXvk6PzdUjX6Z6IfFaR99ZrR40PmISsqwCgXob8IUCndEABc
5/wDTitJMbKqyXcn0qJUtLOQXOnW8phXMq7u9pktfY6rLrjgNPTR2/HWXsSNWiN8cMXUsPsNzY+Y
bGTJu5GnX5vI52a10sWTEEHEsoVNOJXBSQg/Z0gTKaoFFkr2abwilK0QHxqNF5zX8b3BRqn9Zze+
VJVCpJO/flPrZBWOvW9e+Y4OHf1S7NM54yYoomquaI8OUT4GD/0Py4a97qSNc1CmFICVSzdEkUNW
fgAeMrDzSqXytbPoAYcWDeAi8cAHsI48ntzkZDSzsSsx1maMM1h+W/rjFHi3N2AJrfjzTe+ZtEYJ
7ql++AjEqaiyjx2QN+MjmPrO06O9Y4ebRppPfVXhLRyM1JWFHSg0VsbHe33uq9HLOnTROeo7BOj1
B+MPt2OJD8ga0LdHN+tqE89nWTcGwOgsGJro6yf6o+VbTGgHX8NPd6+bksK2DxqZeWtRuBIuBdeg
MCv+aBokKyBdUee9z3sBMmLA6n3oiPOQLEV4xhA01987HhB37DBeFWDIrWUuefrWD+1v+Xtx93FQ
c0DFMu3l6LQXeJxA5HTT+VMLkiVvarIE91DO1os5Ua9IphMl+1WNSroVIFdKOwmqjrrYX5mglTm6
t6kefxSQMoeEBYNWMecqcQTC4alvATKeZNQRJNxZnPH6v1DzQC3kLmvGLnBMKuyXrFXJhvAzTsfM
Vj0Xv/Yah3jlYqMEN00NlvT5dloVVws08ByCGg5rjftzu+bvDX7gsaL+1YTarRQeguw6zkNjBvZj
VO8HnHnpau4jtR2NWjwL06ewqTYhOM/PLk12sWo21mgwdsy9uGwETK4FVECincZE95ceWDKDjA5T
cTQ0xklXwtIRbZdkuEsM/AzCd4qk11nHHDQThwOJFV46jdluayh4rnbcv53JXUPwCv3HUGqtTBmi
0LI5NUISp6Db12SxBVDqbB2b3//cGaFFfpCfTzP7BoGzjz4OzXudJxA/PzwlNs9fbwzAJNFJMKIj
j+4PbuH60WV2kE08wuH+919E0Ha23BsEBGgJnfv4cxTcmnSL9gEYAhyNPn9hl3hTyJOFG1G9LQeZ
9+cWi7PNR+JIbFF0IziKYECMQAhjGId5pgigBJ9dPT7jyQ3LKtk3+2J2uqWiuEPzpKthAoc4qKmm
zoxEbRTAyChqB4s8IL9cZXMyYeU48yktYgOU6LfD80gQmKXYjustNd5qLmCjTVlR1ddFcen2Mtme
VtbauDB2Pibebi6K8QCbSybJSN5RNw51OdzsTDP/W7KlC3ORDgihsrfYXQhjcU+y4YhSdqKrK5/Z
LOtdwUYFe+OZNBjgHNUJeQ2Uxw8X8oJvYohFnrS/TgyItYvuG0Yx9s0kn6VWbyEdtdiitPMcdZvR
PhjkKHCUdP0BAswld8LeKi8jgIHNVT2lZJnPBzYSys0zz4qPC+W5JNnxIbW6Sj6ugPPBJdkyaJyD
QxgXIs61SdFTykOBqC7yFpAUKuch6xmQ3qyctno1PRro2tuOnc3Vi9QZFRTmHGLl9rtb5YoWdfjb
NlgNBPseACmChqPZFugn4S/1WkA9bZ1ynOQKFfuOcIiDzi3VhxjlKOGHoH568Ab41CPCBrWGLR/R
S17BofLgKE4kniSYY+Qahvzi083vmq3Lu4VBBTO92McXcq1mBrVR3XwxdbJ72OVuop+vBMEHdcr6
aV8lfr28uBcGg5Tz8Un6g3/82XGlkhBE9K/r/2iRP3tnkPDh0Dr4LxOO2egRN16A19hdlPmvyIzj
0VAUubPx+14NvDRvnr6fuuhIJ/DaX+l66/+DQlczVHcz90Umhfy+JDWPLOl0ZdFlSmq4qhrO+Knv
JLENCDF5uxjxgKzAWGCcqDR8hWVWIi0K+CSeA2WxMH0TNVIUcZkZh8YKWVsF3J9SK9QXx6AqEkaD
cgRy+qW8gZF+FSvZTnYgfH9awvXzyb8mZX3JbLl/rNsB80umRwP1cWyUnZ+MDI+UCMM7/QsmodEJ
5oP55/kpHPlb1Lpp5cbKtTLDHoUuZfqEVIvW9HBy7z7Y0SI47uuXL2fd2Vpjgtp59ePiuU1rGhE0
GW6LRk5KbjSyuwgyxZTA5tHzi35blOWDB6faFjK+xfOndu9fUgRZpu/zlxkuOSKlRo72NuOT3I9u
HH5SkzHRieXOdVXIacecBqHnEiPj2YgQLFXylUIg+7y01ZzkkfkagGuaa5qTTxvvInvVvlCLssJp
I1mxL5bVHhMtlWO0W/GrBN4Jm/OzPgq1AuQXYgy2nAWMIK+8vaAO7iuHAEDN6Ee5fILmNI7QWUaX
/fg52Xgh5Rh/S0QzXiFomK3Iz+JgeDhafCdRG2bOy+V0GmRuQoi3d7p4dtr2jx4xeNOibvsA7jIP
lq5kUizXPcTwWnSKa2zYuKHTmsYtIIAHIcvUV6awkKIUuYidSZlLRkXx0SW+BHcRkf9tpgZvuXbW
ZyVP3vYAo/l5ZtQ+m/p+RbMU+muzjlTMuoFe0So8YhXVOyDTe9WFTnEPY/AhlEUyNJeVSkaZybYP
e9Da/UwSo8UO9YmQvWgnzxxwEr+F7xakEpqGd3DnsBZhul+iAkFHxY4MQC38qqSUsU9yemv1X/OC
f149VkXCXExj2bxlFiTliUgez6AjjpoRHzB1ZFJJrwNMZ0EheXVDlDuaMI87ARS4n6RGd3LXmgsU
gMdy9hgKTRRBQhEGMtv1O0p3BV9tuxyZ28PVT7wj10RTf6/sjwPg/SoaWdv9kF7GVCoq70Fu5x18
MrfaVDbDg9UTKtX24gxlQ7kZd4ewfsX68NS85GZeXKTkJuiHnY5A09Vexyzut6oB2F9K5cf+yESA
6e9OnEFjCIQo3oeBoNUH7Te+DCcw/plXq8xUVhiEwbUN5L3DXn6q2Lj7jNDY8pj6qFAuF9X5qW2z
FDgDJQqvEJnyTmPCgFdwOej4wQUZFBH/RgyBp15J4c7gpkr8mXdiW6qud1x6vrtZ4p9HidUXh3dA
/Y6Xz618bcuOW5IZnpeF8JgQdi2Vk46RTAj0pNzTANrhCbcf2OkQxAxVOwlPH5ObYdPbL3EzrWJh
Hd3MpOFQQW3d2z7WhtI6rQ9dVUlj9kV6qcnCGgI2ti9nQTd+LCZWFrN6QXdRMNZR5WaychTH4YK4
eGclNO9EDMxr8pduR0cvZaHzQzpYMOVT4Cm4fNruXqhD5kbuffTxUvSUdsBo7nUKdjGLh7etqWed
kxRR6EFaB3tr0h3Kgdnqs0DH2MxEHQVw+fu/0afUAZl7R1gnO07RAN9wVQ5dF06cEPvgzVfyicz2
XhWs/xPQo8HAZOSUrYvLeSdpIFhCvIIqbHbetEGtsS4E0lpsPaDFkzWKvCIgosaSADB21gx6okWc
ED0AeyWmfbPJfB5TPECFN+2U+ITzCUrHQnSU7SSzJEWSnWMoqOWO8viwV3Kss0kuAvm3Dm0742HE
7SyxvVpOu/+OoIz7Z9EX2WcQ8THP08Z7SMQXtestheznbByv9acYndaW1/e8/C4pOqPwLOOzAY/D
WVKe4v2z4/xN8Sd6DgqtBpw85VUcCtJnywfejiRh2PVaa6zoHThBhdGPZFan06eMHG5o/6RWhn5H
kvxSncqKXrx8mfKr+L5BASHtJtgZ+gB/LaFVmgTR1vaZfFLIH8g4glAKatdmAgOIEgoHKEcFm/Jd
98kTnLVn5TsBL+tdUD9UKp97bhS5BZpGeMJHWJS4E7pqtRgyrYdpRis3lxU2Ty5QQ4UonkJHeCml
UYvyQNUyRjea4kTwuaMJViS5d1em66AhmUjm1Y3x5o2pibZZhp9mn2jTswg7ry97Gh7Nm+ux8viM
stK21GtGmGWGhLGIyCl3QO7Z+wEV9yQaRWV5oLOHVTmzdXR9kXvRgiscixFVnl9kp5CmjAkjyHu8
C2RJgHgjQEIhXmWLsZO1aDDWVEPgsFJTH18J39yyvYNHfANDxDSWypbZ0e95G7G0/aC34yixUvWw
zkGSNnadiFJebNFk94PdPR0if5cQL63DQJGcFGb641DVGoqtquk64dBl0D0hsdGW15+pDK8un3YV
lEfEfeKAgQXdOAGsUxwvKpKi89ivxryH8eKhG2CG3icm64/OISnbrxTxIeYPMzB1feUoMQzy8f47
1+fdZa5le99rqsk8gDCnd5Pload5kq4kSSFQEGlNx99o5PIZqwT+Jbv5LGaNBC/X2dQ3v6cMSbO2
QwBPb22eWlrfuRK7WIiMrYphPZPUUUnJMwQthttWjL3L8kddPl1TMILb/1kmbh3jGC4RJBxox6NK
bKr5A4n9jDv9Us7C3PcSrbnhdzdK3RTz3GyBoVuVj2McNEnyxPwqaQoonhCHNFSInaSWvNEg435S
Hq1WOPzLC80U574BCvhWcwyei5kMJ2TzZJffBG1qv8Jgc/kBXLJye+vZ2spLFKADaxhTu/JTzVa/
G7pIkOq/1F4AzcttjcAixl9dD+T7vXfUf2XXEQaTHhWcgFtVVNOIXj+QQG9R9mb3r/TWBowWhol9
jRnPsaKMsTymSQ/PNjYfoajVz+C8THh9yc2NdjZ5BsIIlHnvQoSxYgyqv8qkOJiwQFvTR9vOhYZU
WpS/IDJvT6PZcfSKBvsAHSF0o03J33rbSt4XJTkzYNKGZ1Zj5sC7wlTONhNMCQLGeCixsusYlzkJ
xA1i4N1/tStfnVxc14jpUiO4iDQd51DRKJhaPylMi3vY9DwIY9QvjMB2NB3j+4ccbGtuuOktX2Ai
dwW+XwYCiyVIPvM809LMjI559AN1NwomvUvjItEX75CfwYe2djyj+GPDq2liBVrqB7cZuUnigKuy
/4isYq25MVeY77lvpRMaKPzODlW0qEUwKCrA6azucDQ+JDCV1h9arZF/XoPA19X3Jn9SQpdKnAAl
QHdyNKrzvLmdfuy894tlaKYOxZexSVKTfzCdOowM4SbL5rD1OVrDir+gnwNN3i4hMkoZ1tnb/cxc
UiaM05SEEDKT5EV2fr2SHnTY4msJ8VXADskfjW5fTTM/KL+dn1T0euvryKU0SFLXeMRIrFnUagZa
rqLNBLPBISTf8wDNclJXSOOFjHf90soODWsxXTvqYtP+uRltdmWXBrMR1VPaioebJOLpq4kTF5sK
RBLtNvlhcwgdhz//JJkkTqqSSOJyMRC9ny+IckLYN3j1Z+7yRlW+4Ey4FhqY9+7L6oxWQTYg0SNu
CTufpw305GNvfmbiuxrw5iaadHqxQjmVDzIMqRQQpUXnYr4eVA1PwbKIisDdNoKkY6My2Bc7RZbT
k4pcteqYbgNuOpdpP+u9gJpM3/RLbw3yQ3j48CtPLKNVqB0CDhV6o4MGSZvAmlZmFKJ3DH/t/vnH
/XRgWJx9BXSUqE2au4bxx9FVoeYD7KBmDqcB2Y4zzk26A5RmUVREPaJaE/co8rId0RnC2uSgcZFp
vfqrS1aZMiQNS8WaWhS/tUrg3exEzcL5LrPL/c5KX+4F7qbZdifnBJwivfO6RtUHDvywe4ETkeNQ
IiKWpCcJ50tOyil+galxZRw3l+/v1DWatZmpPGk4BjGQlb0fgzFgtUk7Ug9Bp74d6pjoAKd1BcaR
C6kcgFj9tIEAQjifXFojdO83lIVu6+wrCUyKBKI73pv58d/Q9ehq1lwIG4ctxxWh0eHpvUPljOWl
IzcXkwFrVdy/sJqUqq3X6od9RbPZFuvRV2GlF/IWLbkG02bHFpH/XT9MZjO7efeRmiAjVFV51T8q
dQYluEoDCWO7S6B0HIBhELR4cEoYAbt3EYp/gD26Lm71tAD7JZlJx7/YBUdJWhlAXJJhQeVTioYy
fr5OHCk3rNOQxT6WhZaLpxSRSAtLYQXnzPU0Tn79SHqvyuE5BMuAnXQDgK9lthXJNe+uyg1XE51I
OCH+rhICrFACTjqqSglMuwn8W4Wh1mMtowc4E/MMmoI+v8JNGcrhzIR1x4e/NvKU8wdmbCl97Ch8
kTpxkrzv//iuD66DG3PO9ZCccx1z+EwU7qkd4lxcFo47P9zXP0rDel/S+IClWse08jio1rHxhFX1
PMiJKChVzfAOjeWtmE2ww1lK4C48pDbvIKpDY1d7Ljqt/Std1+MHX8A8PfGXpZycyLXJ4j8Kj7ji
pU1ptQVUluikVbzHt5M9SluIFe8koU3/S2tPUKHhOiOsvxt/Iy6JzTfjOkASV6qby2KnaOa0EcBz
8V28tXvcM8eSEXP3nyqlHXiBOZ8ENWWdrRjyuzVQ+xXl6ifHMZ/cfbHwkoVm1+jfouOuuaxcdB52
qFl6X0IRLuIM2wNpX4FK73FVNf7MJDPxemLa6yx0NVX9bLS1enaUsa6xiRMddOno1CmHUxkMQyMv
225EnQ50+UWbPgmSlOYAUglY38HOlSsVivG2Yu2MAnS/M2ZNRjFHaiigkmEteXjb3/PpJPWZwLEa
29UNcRM5+ShLP55JbprEj1JipdpW/xK3g8lL8jg0TeD9iVHmKLJJlo67XE/ngpyHsf83Vlk/Ct8H
ZubGFe3T5uFZR/YqD0N5dWxe73OsUBkE0/HR8qh0bXYHVZ2MeKIH/lPwK6pnCD+g/VzvUFLaHiFk
UhqikeQVjQDE4JKl1X/Wq8bndyuKS8B3YmIB9PzspRtJjQS1Bh9PaFUOxZWji3pF51TQYwrafuc3
bAgcgpM6QC3lvbX6a12r27vDgRhmezJB9FJKucRH4THZZQzbQP+q4BKrcmORn463Gxd5YJU1OpAb
vuMw2Ytdh59aCICQd5MXjnyCOvQZRLPuMdOPFBkAgoheECYJH+0nfMfTmntEeCqeuY7kDNjsbbC9
Ds0cThOFExCo0itG+xBwLn9VkvAOe1rGc+5IVrMoW8OJE0FDci3KnZwoZMXULG72shpFUTcwQ8u/
z7psAa38yMSo3xCwJ9y+1J0uqM0agdEfP61IE4RPkjHZUztDnvfNPfZ78JgNpqyCiXhLakQw6g4r
ByD7RpFhalwB8y4bbeJmjGMcoOb/R9ePbWwi9HShwsqaPXlrMZ3j7QJNFZ8C6Vfj7EsM3X4rro9t
xzOMZHcQwLn7B9mScAKcB+U34tW+KmAdzTWfABintnleTzKz7BLBONlP2AGQbUhI8d+oRwk4wkyD
Ili6zOR5R82QUvPQ8gpNpsu/YBNNQbach9gq4TAYKAny3qSfn3MzfRN7ZpZzvPngyPV5gdozTUow
z73nGedIP9i0ipb4sU6GAk7pM65g3AH2iv2T9UkbCQA4N7ql8njphTmtJM3EmkBeQf9UWKMBu49p
CeeoW39zpKbxJnbiVXI4Sm5ix1GxX28C6tmFI8wVqzhlhjW1dWKs1hYetLpSbLVt7jKIHmSa6tZh
RT5BRGYmhLveMNXZMuVtEKjcJDqS8CqlX68ZgOXpCaniEmjrTgpEsw2JxTLYqhRZoX5CdiMawtYF
kJAHuzIe0+1WXwuYtnlmmVFOz4XRmG/phtqGRwfjTWRIvHVDGWjbR1wMwXep9yvZY5+N2AyfDnUf
KI4d9EYjlgFAozQMu5RvjE4UkLybtXLJ8UiDE7NYr1FtHX+VU0ezd087EJiPK3n7u08PaOMusFP4
fPWdza6DbfQyoV7oLIKbAMua/9r46XOwKro6HcoPgEDx5hi2ufi4tRrASsWOH9EoeRFHF3Dhtm9d
Tm1dU7X5jErzfty/zk3KuZGpu5BOjal3qnODqhzGEEBZfRQXpDZ5JOEe1z6QxNxj0TsjW1g+RAcU
MQtgooxiKRLXRVbdb0PClZP4l6Jm53ZAoyS3p4H83B/kQNP+ud+WZ5J5JSVJzzQgcXONfC+aTqq3
/xM5vmCbfbY9K415WPX5Pv0E42n4FEUrKtPpw03+PlkbtDYmdpJO+sL2NNa+5kvCpZjOvo8yV7jd
rfwsxk0LVU98uvDK1HKYoVQl6HDeYJrZr2WU2Qgc78170euyMuR2QQ/gn4sBL0fOrFjHb8/O/j8m
zvUhQTU+EDkv+KBIXoCSWlMunU5T9PcTay0GjxUYFwjJXqWoGNgL71VrhU0RvaPPIGFneZV7Dy7w
KiobVEN0MF8ckl4oTbbSo15YfLG8LQI4VJbeIA7sfk6Iqem+YbC+ID6JofvQ39dQH05itS/z73Dt
kErt1nRZ0F6CNEFXUGSN4LeWMkbQFJqEGl2rGtbAt9iN5b18vdnAZLxp91Gjt7sgHT6UTxQ23mho
56rmx/20Cl7d87C4gHutQOoMOMNAyL0FCo5TFmyFJEbo5Ld97GeQYKcYKNDMvLWuzmtS5avhzRXY
wk1LKJ+HCExf/H5rtX8SiaPLNZfwndkRwCToRTYYFr496re2U7kEcktewdu5/oQG3yCtRDwnoCTa
QE0zClsv5a75Nh6Wnwxsk0qkJQoveQhfR/+wZYJen1iT4IHn6eqWrerOOaJh5Cw/nB3eKxDt0RQ/
xlQ7dZDot3kDh1FuXTmSjvg6iIDMRhRrfC97qlpYi31O4VK4wAaGtXvsUr0WOII2SxVujc9NArs7
it1vDpnaRh4MK6hAQ/pNvlyst8HJMgJxt9jtPUzLtnSR2YYHUL6td/FP4zFLGCVbh2Ppwp5MaeG3
HM3wuz74FerpMR0ZUkkOILVrMtbLUIlnK/6ZJH/WOpUx45zDA37y2uZwjN34qp8GYwSmQrtzTE6p
Cp8L15O7Az9OBiBYdMAvahcLZC4nv8y2qgYT8SoNGtfWHEuylKddeZRDe14VRLWzlxvm1qXm9e13
RC3+BgifN7QgvdSaw6dIUAy6BB1GR9eBCYdcyFb7yDctwJr0erTQ6XAKxD63LWc8JXupB8/RSjJ3
4iErJyCOP4GdbfrciTByVh0Jf9qvgpN+r+Cj9M7NrwBMtCfTn5wtxYxPi8G8QOzQisJdMhmRpjdI
CW1ZWmtY3bBLuAYcz8bmzGxNNRWFygx1w8jZe7jO/VGP58UY3DSRjynjm9pU6neiGBtlq9PzlhPw
VL5cJqdYDrYABZKcRaxo8WvZQKMpnu2WyzMaHTOV68Ich5q//YAqAJoxHR9eMp9vwHgzJaNkOo6d
hL3W9m2kUSASpuxe3bP1xzYNZC61n9Ku0+h/g3vOw62alj9lJpzdDY+sQ0g5D9kYaKg4Pal3YgE0
C2DDDAEwf5PYOSYNAs8AUGKzZUuPvx+nGlHGrqKC3BLtmST7PRSp7LgAVJc/b9iLzAnSI6c8YIC6
4tutErVWmcJs24G2HvKlkwdA3FxbztVBV2Wc/Z4odh4gDySQIwTwN0Pmk2xcdosfxO3q6qq/82B5
0D0JfssDDPSwTyUm7ikTqaqqS6dckqoNSdkwLFIkue7iY9pZ418lLhUyFFACWxQ/9v9kTq9cfuow
5QJaHlXuxzBfqdccUOuWIx+fJXH7ZfCHHst4P1ODY5ctpC1KRrbQARv2lCnbV/QYM6OmHg4Izzgh
jJmqJqUld4DL/K573Tvao9uBuvG5xpbWHFjYSxUvZxcYayjPGV2VZ5Qu6ua61W8bxHPIEdQ76pc5
8FbPswm6qg5/lbHu/V4KQRqx00xVcx5R7oOfT0xL/+fJBPyx+Jm28jvXS/ggt4WYyHLqu1RymdFv
MhHmeudP2EqUwz3cYPzTplN3aSWkhYmQhuQYNTL+vCHWiRYRx6dwu8YnlZAeZVw2CqFeEwqjibld
Zlrdxj5PKuHbzgJ7jB/gkIAH18mOsKKfIDo+S1H1ezQO14BCH/Xfd29RWpFCxNiPSNWmfpQ783KZ
XZp4e+/tlNGw81C6avlgzgYHgoMv/vm9Ju1gc0KETv1G1H5BFTwBr1Pi860hYAv2SS8h9sHDAi1a
M4RsLlUhVZ+K4Pe+taXhHp14XiKQ1svpJMDaiNaqaGVmXyesU5eaBmHoNfK4bxYdatCAAU/gGdw7
Xn+zCe0ecvGTrdpoKEm0EqiZHFy9k5/TQsB18XlQQDtIxEd97xmg139aKbRIObwA0QtKLE5+NGZV
nN2IUrKjzswncVHW+/+k/hEggYa+eue47pPNJ631UUwU0L0p9C3c0yAAETE+1ZKwTFNu4p69jO1g
pSFB0X4/4r/Moir09HtoEtYv4SXdDavFDMbBN4YM/5Pq+yCFVSGUv7PGRuoRoktItpwyLyjtrjCP
hDm9LiuicLpI/Llnrh5ySVkWK+e6xDZvcdB2o+P2SWa+TmZG6WlWllGLQ6qztAcBxHOHFQgr7F23
/qLIwUg5eozGtSk4OAaYBjGGyuqCTCz8VCXWohEL3bzDVYijTHOF1VBQ+gmMxrPPB2++nZL9sUFt
Ax6NjEqL0DEROTobpoc+WEidz3brAfUfi/H16oUEVQW5Mp1EvdlrEVJI/w854szg3s6K7f9Wj4nm
EEKfZX+7ybR8f/zOEPT4ta3up2m/9w0cj0rXoh8IyJZZgxetVs5O5y4CW3Q7C2xxmyEIPQDtVBWs
WYtr03TIoX1AGfp2HF0/3XMajtlwO0RHynVk7cmY6m8AbXeW4TOmmDU7Z89znr+WOS9Xf7Ok+yT2
AfTw6sHdQj+QuYUNrRgBwwbrsK9DoUQjYSP5HBOGzGUMSvmTT67BVhaVGjc8m0XEjMUbtjEiqg8G
2azCj0ungOWIpeCwma/XXuF2rhQuWwprb7XegbqmtGb6fj4BKuoQcbeydaPGldqwywOE1+zZddxa
hdEMJjH2xmBhfWCjb2pVzcSFh+to3OP5ohnQMFf97MikjJHKic5TAE+T1FTG6WdLUIBRoRs8BRpL
+mY/buvL2Cyo22AB+HrloOIaK2bKCAjTFhwqvig35Me4bpqiBmXDYyNXoosA1Hm0KSAE98nCwNFO
EU5dZ2FU+LXVVJTKJMl+9T7ygu9fSF0QCGGJen0NxB5UJaqV2veSBIjTLyxxTRznWdTbexO0Ps9/
S6l7lLxV01zoJxORcOTyWvxAqUcgZf/RCY4d2/JJNO6wT1AS9K3g6vpRH+cVyGHYqgUbqjpoUgPV
TiUU7MwpOt4H12jgb7QlI8s8rshbYQSEZ9Tsia1moWmtFbFQj9t5k+xQWC8XYdOvrkDWtEMkysV/
1MjcPbM4cfezOhMGtJ9dTPPScx5HXLrviFVcJXZoatkqO3BE9g66GfLESPrePK+Nshbd/AoYvAI3
byViyw/6ROtHBvqolI68cP7K1R9GcaQHSaYrfQV2ZoWwYB3tYltLW3WRxekbSpRxdyjT4GnIZ+16
ZEovdIf00D+AVvD7NN5v8qXvoLd4emRkKooV4CLtZ014Ir0LQXoDgi0K5p8qnm9KJer01zoNwnzI
tAPwwUfXWc0+1KD3EbR1WAtHX7UOyi8zAiG4BNmuQLDq7a1TAd69YL6uojOTtoaQ58/CCvt2py48
izlKj8G9T7lE9f26arHhLflqcgGVu56CtdUT8qbBDvRUtdoAr5YPG6s41tE7zIYiVIpwCKKrBfvf
TfrIT/rtivHp8qOADSMZ4PF9tX7ClBTchZiptejLkgiFccJABdhMZ2kSO00WIc8PyBkUi5JHhw9s
ZhPI3ft8HolHTebl0eUTp4y9scTm9+vbahVHUnSTTaX5vVTdcXgLddNQ2lluPwj1ee6BKH/dxvcA
2yoeFAEopcTyNQZxmKfwfxiwK8hq9JsK+LGgZcRY+xhr5VrXQDn8b0phLzQvn8K0YHwmeIQLRvlU
7MOh8bZCFZ3/dD0yls4QLzN1Gv0WqClZIvinApU1Avz9ELZhMLolI8zTE7L8E/rA7Xdg1hC8VxDd
GWN8HXbMz1TiH45OKLQzDTAMSnYGF1nv1EH653jSZeLBRNUyjYVonm7YM5dk6aMRvY4AIqADn+Ym
I/xYCi6/L/C7CnMoeEenGOKSWRhwTfV+yrSfv6PbRZJDAMbGI6pjhz1JXD2LVXJBSshOoRchuVP+
stg3Ns86WVDaAuY9s/PETrneoRoQP62UO0TCyCsI+OmUiJdVqanUVyAQ+NTkQsGgdR7RUPEG8eXU
aNA7uRQ+uBgOXBCIYpOlDKM0n8Ty7qoDYp68G2LCc/jCq5KCHEdEp7KffokNes4y6+7PJpLKHSLW
N9pSV2CsfwsLhISutAcbwjxNvm6Eg3dSF3o0kfZXgsiKUuqRMflCNYyXpWfV+De/j7f+TOu5+yA8
1nbQgj3DtQvFQvPhoJcZCTJJyOMkW5CbDZYXB7dyOXjplfxxvr9FNiNzyS5uRwwUrbs9aanKceHN
rfnNOPRYEfcwIpDaeEilr1nlvZKkTcREeUoyd/AkfYNAuwrK6+9pq2H1UwSCq7tZrqex/FvAx/fx
yyNnDEr4PW6P/mC75p2+Cr0KZ9Tm++0RhBQDkf+5MPozEobe+5meXkubFa800sjsXgquX7Yd+93Y
CBkA1YNSdv2qDr94ipU1Nsp6RK9V1RKUGdLbng1rrozuQuYeESugxOBx5//4DQf1OZWYlBDPwG+P
J0qBC+j/QbLVpbk5ySTALqiSiWcICGUzpQPoK6r5/AD7B9tzq3QgrdAYUKfYnGQnrgvIxMIh6ljF
Vl8ZJTB2szy3x4oEYlPNLRtIg/AApH40RgYU5PmA7Fc8Cp7c0ArZosYxfa6XEGlXY6PAt2uO3RTC
v/JtXchNfb6d7L7Jxmjp+BAt50IBSDN1iZBUapvY6BgJQUZrPafu2iIBIkl21IwqngZHC60zzWSI
CTcr007cHsCvhCvGPkcmopNN3hexboSROBU8shH8WyoK8h7SALx5AVlNbdfBJphaLAYrG66WeGHX
VYvdQdjKVGpi0Z1pEE0Ozq31LC/a/k9l+Dnx33eQpZBRcxNFBgUM+Ug6nVuaLjuy5KAdrvMMFZgB
HyLIlYAochaWHbt6BVl0n4Lt6/nfHEYNqzFAnipQ8noqiLKb+LaWr6VKQLsnjnVKIcP7y4EkEO+z
DVDaqFG5XH6WW5hfLmqUJb1IWDLPo5tr1G/MB08yJJURkjMRQRp1h+tsUf6rrFrvf2ZYF8DXdDGw
N3BeqiSxUGY62A/aDE3BQaMMEc5D3VlhpEO/aHP4ea3dA/3bvPTQrLzI8dXJFpmkUUHHDvhqdVY2
lICM5vtw5Pz20XimX+ntnfXT/feiTs3oGuHJ1AI4p+wDsyc5DLB135ckgE1vwe9BofT7kDmf3xV4
kMeDVDx/bwXRYwQEDR0HZx79O1PV9x6IvPJoSRzaweUCdkz6g7uQHXvlh8C91hOEbnpQAcR/JEBO
MqDRQm5jZ2Suk4CpgyYOUVHAjHnO2JUYGhpuduVZt1hnh/j2nsHXwon9jy8v4H0yCNbwBVMjBymM
wOaILfGxUIUIpuhWgr+khEEI8WlfrM1U1MQ+nx1XeH1Net0GLKP/hCGrWV9emznxxSpFf6MlRFe1
lpsZWKMTowgsIsp7eo+8cPBuNiHHzKIeDoZXG/9LL4jWuMgrFj3bFnTqhP7t/YSDvuUDy+TLLnnX
DGtfl1j1l+kdgqzRc89Y6RqWjS7eEDBVQ8uxyEeBnniTKIZoH+1YB0qmZmwO9+BNpp7OZak0hyfI
qgMqQbqQeAskWILhwGtgB2GDLzkCafGtUJsTaKoXtb9IsJzRcrArism1+dKuHasAOvNBnSkoxvG7
8+2/khR4VOCdV0JFp6UB/yCLF1ltg6q3bsV17zXtlvXfqzptqx9WSKkImaqZpHf9WkHa943neaXf
1vKBtpTAiLcJTK6GZ8mkSaqrHaxR9xV0EnrftBpKToyvtWwqdvR+sPYx+w9VJ6Q3Q7528wlpBGbv
x2p7Tsg6vM2nzXtB8aYnxIPOCHbrtFdllz102ZJa8QIQ/HnZjCXYOWy5bGqqIN1OoFBQDdr8puV5
njAQ7ySh0poGQKtZttWxAelFxrFQYErq5hYTm7X0ECREI8EeeIJngtZTxQDqRFYQOujkouXGH7NX
ERoudS1gd68wXvvYDZ5/JqylVGeas9E/Os/xj05GlTcPWL+ICsOkf5wGyNKqJxRb7VKdadtvxdGb
SWGgkm4tH5B4UOrdfU4/XszRkWbU6iHPvwzZRmZvLpCTu6TNNZ4ee2lfqIV8iaLMK70fVDQz7Pjb
e8g8y4JfHrKQVQc4SKPb4w2Dy+RvXjAtm04RNpnbT1mmhyKeEzxAUgN2R6xTynLxJ9iHYxS8M5OA
rnOyZeuolYplDWemcKuEtm4CiM2N3wguzdInGahMB2gFwB3aEe+6Rt/mIQC810Dwmb3mYajjcQ/s
iY6QxHqMtf3bQfjaTc24v2bee1i+CNNzzAD9xJ5qlH728KV1d4IA+v9crZatKhvH3LY7JnUY39gF
vB3J1sMTG7g2OYylZl0h4qlPG/CX5cSLTxATw4Vl99FRCn13d4KzP+XFAUOTKc6gTN2nEfvQoU5D
UM6hSgW/E/tYGzan0yTyNbLWAWT7vB2VmlZO3QIcTWJ2a9rhiJB8hX61gw8vHwYVyFphOpZYHrNB
LMEvcuFqGhj6XWg1D+QOy2XQeytL89jDLKq3d1ttLKt2mhNFS/fzmesUmSl1l4InRp9cDjQsEL2v
DDboWw7noIBbL4eYLJaPaF6DsZLbTEYjZHRS9vSVJrGr5UxQcE7EGwC4s/LdOyH0KeYSRzXCnOeb
sRXvEzGD6+ep+3tlqeh3J8Q3ArnK5pA6fOpeA5XKCRqWvI6V70HiLR5HLmXsdWrvmGG5qpVCSe6g
CwNxQ62DXHf6fzgvJ5dxt/OhPRt0Pffyf6N18N7CwKSo9fbXl2HaaakDvVc2JFksHfkI/2MABZ5g
ulqmdojbuyvijb8H/UadnzDxcAPOjBvG30/xm4a3TfZ8ZSCB+BDc1xmuBy4m667a8jlk8a0OxiSM
6UJklsIhkX1dnZFe7T6C5YFIRu53ER0axVhNXGaYCabmiShWb+DSpmTlJzDuz9mDlzU8MYHJ5HJa
5cxoYfBQ+AVW5CABaIVc7yq7CPZ6AOAwmYJRN6Xo/G1FoKRNn0DeunTdqMGal3Kq8HNXXJTV2n/m
j6F1ysucK7p5b5PXlllVsDaPLWRpydnbljv6pwagR0/LzntF6/CcesObg4/kspIcgfqScRgjqscf
I0OkbE4pUB5oOFRIVXYEp0K2z/Wv+l6QyE+jE34Lsg/2G6cbw3TJBN/BpgjcMBRneh0elvDk9tmS
rPJamDQihiCjCqmLeAcBVIhMpwNKTcVX1MEZ/tyXf2gnq0N4ONGHKupUHCCf1+sBg2ESvp88Wzh0
EoaFACHYyjysnK9hKHk5xszS0XK34fWFdFku76QlAbaSCHVh9jidyVH736Y31t2G90csr1tCe3FA
0x3bu/3DH6M24PrOLgmduEefgNjpbeDzcVe/s+vy9IcZVCJQoTm6uMjvAPVqatVYZ0Jjs8rhYMgb
aj3vjDtDA2mgPNKOrXqYBzBAm2B4zFd9PEApU5Gcxxg7d1PpB52tuSL86mNP1qhQYSDoEHznHGG5
hHSnglzBcArFpqAVxi9XlvGEfbM7SaueTc07A+LkLxt2DAeqI6VjE9v1r0iLnrEGHu/JCeYRfX0q
7pUFl7wsqOJjXY631n7R2ZatCDyhP4vAZdWOW7lICKISoSiLUMCabHxuS/4d0aH/COgfJwjq8dDL
6EKpljVVJ6xHwhcmolAPcIGG2KsxYrW3wvfV0VJthnmWvx95fo85G6YdJOwGLpDHSTRGQBFLffzR
TW4eAZGw3gpSXV4IerevM96huD+D12eCjN02Di/c7f9/NFC6q1qNgksaC20yebbN3wpc0cUUlDLL
wFpqqZwztmKf0ITJ3woab9Tvam68EhgX9QiS5XIPA5id73NQTVOs4owqYn0qXDealqYMr0+RpNN6
Y0QXTC0k3b8jMDX/InTHf8WdfZ/ZarPsOiFa747SiAWyiT+IF9Eg7BMQosre5JGTjnds++HdS0jx
Uj+P1mGt2gN3xRxIj25cnqP+67kuuTobSTWDKM7XFwQkXBkkQ4ZkiAwQQ38fBVbIughcxB7og7i0
Sei14uqhalNTiKzvsD2vWak+SYySp85ETr/3Ns3eRTMYQkcLBLs7rKnaaW42oH0fRkOh3Ej354Ko
dm0wc9CKrXvXicH0WCM+ptk4yfl40I7HyX4HNPcIEjMCEjIImEU4lybemovPtvVTtuSlkeHq7z0B
JKVkTImXaLrncFKtOZFdnj4WRyiXzpbzeDSQyxVAY19kzhmYOp3Hg3AzC2BJLDVC53TlJtfE5eix
4IjwDpVa8oM/dxMiIQ9GPtblhD+fMYyzNZtUvKXGypnzYrcTEv7iYK9QDnhMyD/N0N+shHE1S8YW
hsFMazRE5+3cSnoEi3PzzLcI+3TdZjRPB2FZ/5+95r5PpPANr0ZxhC/ziPhsk9Adq/TCqVeOCLSq
8WGcSmk1RPib2QQH1pz54uRqClo45oMbamMFWVGi8O1bI8e+5tUuqnOSVHWvF8Pf+LYR9CwxE1i6
YWIopK1sXPrzsVuRTfJQovkrZhZv9eBS37GwhHSGtdTHLDpSsjs6rkto76Ik+3SZ3HY6XDuSTteZ
Sw0fAkTDR/HB5B53dCJOEqqLPRHaS4mn4D9wSooyc/VJWGrIXw7bqEM0O7QgyzwFbHfmrdr52aXo
nPACagzKu6IlsjseKbDXdMA0GwqNRVGfEq1+y1NxSCd9qW0/diM0QZjnHQfBdWBejBQTk8ZY4IBx
gC8JmiGPL73IXRUav03CLia+ovTx2kBiM78Y2hrCJBPGgfvNCqiML6UNo+semi3WuETwzbrOhNlR
jwgKrW9OgXcVVm9gIaMxo//cdXBfAwWjFQB088iGgeTUbkQSI8FsoFIFoY2buVV9HfYA+7c7OlAm
hpqj3WqJNy/1PY0qMBegpk8NTGuTN22gxit17lu5rhdI6a3aeZDCzwgvW6A2a4BtPxGgfhcJor6G
JUaX4EZ4p7jP34xvOGZEMkZQpP3hgKGiOW+qqrlEfSFExnOFjfBxnueGQCLUrs4C+6nX5a+lHSZl
6pa8j20IcXJm6Nrs7F10cLKrevKWSAcsnMl+0Yt8VujlS4EFTcw+hM4yz0wxEzCAiAjnLjAyLJqt
I1yaZvkXJgoayWRyU+4jCPJ5NkQBheYJWFDzdrTrjaWsNEpltg5o/fqRqt0+FahcPoepU6H1isej
ItbUHXIWi1sTUeTt87hPc3Q3j/Y51+9jGWtXB9vh4xlgLgzkr0ffdEPLUiiPJ216o+qt+3a3JW+d
a5H5i/EQWj8PpRSxkcsX1g8xf+CERFiNj7EW4Fb1DGHrPQiadmSKhcWigXsxpjSep/J03IkEG/w9
LlO7/WGNIBanmhpuFWXfFSwLg+NBQ3PCU+NQlGKZtrWK+6LovokAxeiUtWGyBKLSEUFW/5sKCFJn
IiwXnbo5uOyfG3xQCFHJwuCvL78zvreBIA3fIE+eCCZDKFPXE8v114euq4mRif8jqAjTynIKFZl1
p4q/9bdLyWZ3tKkzWykUbX8h85dPTGCEvDPDVJHlol1i4XLHE0KLEhHGcaGCei71kxRZ2Uv2Num2
tCaKsJISWIF1F4eB2m+KFEqpm/pC5m45vPpF6A7rQ7tqVhZLw/EcAGphNwgoIslav5w/x40Ay4G1
cVOBmiyD3UWh3YdeGHGdvrapLxVFVT0hCWbtn/P09wGTeQobZwIbeA5uWVnNpyUMv384f86HVgAk
wleICuq0itz/drToh2aiAkNV4Ciz7zpS6nf07Esgqg0Y7Eciz7ll8AWGOjOkC8kt9OotRiwfjUKW
qr2ncAiHTo1EU0QUcpxvSS7Xe8F44cyw0Iv0hN78pwZuNsyUzsbPyR69cVJ4vxumHD4L5Ilaun47
prQ1f+oDlmP8W8SOBC18DVTBzm5Co3t5nS2H7zL+XvuGOclPZPUM/07mfnMegEkMw3ItOkK7xbjy
9f1qzsk38BwG4foZRoGlbwDkaSpfgmU8DUACwF3Eqr9ih31/LppRjMubUKITJ6D0l8l07ELSWj5W
YN3DX4L3NPrQ+di/hqZMBHBdhStP9k63FGiD3cGCG+HabrlI+VgcoJgq6BT3XJfs5P0SdGm2jLOm
Tv3zzemM4Vtm4EeR+L3H5IrAh3OqYWNXZHjT1G4Y0+Wy6vVJwNIPmsdZsovapdVZCotsN6QFM9q7
Z+oXvFhIObHFsLlSIKcQhLwNNeQIphRkFtd7vEElSQHA5wJ1cItW9dwPUruxK6MgtkSQE8hsf7jZ
w9tw+VwfX1kF6Kk5y6NShlo5B3i67rN1si+UHO4O3qqIfPaqknCHuuZGmmnyASePLPQhMxkeNSas
YGcS+LmAMO+aYfSJ5YawjkBncY4eRYIKr8ra9ZlKnA+eTE0EyrxFCPvsAzgn9oWsPZhpQcn8TXx9
/xM+0ZI9Jxx7kSwVsFsK3h1af8f0//gFdIvJ90IG4ktV9rJ9x67lvF2gh7K/MG4/oCiMadL8K4Nk
vll5rBxhIq06pr0BF7m0g6u1xiV03CfeqTc012Qxkowuocr9tpUTK3fS22t1/OHweWKTi9DPZezp
hfEf8FQA3x+6Apahx5ZWLepWTzonGtYpNU1l4inCb9L8LGgd+uYs3qKjt3Y0rkm8i/YKqEn6ORD6
qLQERj7cynEYmkDJV/jJLaz+dvA4UnfGAqDNXbkwM3r5037DVoL4o0dCbIxr9R++YHTbbNDVWO5V
6+qT1ZnZQUxAqxacYRbnonmTteekkcH2mfgshkCjwxxuu7z6pdUWST/AeTwB2ZwrSOPY0O2WpBZA
QoBIb/etNLMizyqzGeNA+n6Oa2fvCYRcNEzLzGHJqlErrJLGNoTRozBy4pfKzoDRCcLUAbMDa+bX
U7Ly7DXPxKdOAIwZmD4Mo/j4FmQEf4ZdnEuX4WL7ixzUp4TDhcnj7xdfrZX81AK6sczVb8GkVG/u
TGAxKN9J/+pUeafn0Dga1JYR30kSmKG0DB/LcvrtZfm+FQLMaW40pHQJj8hgm0bE0LJwmOyOEX/n
6jCjN9PiYlX2rRArUqCOuhm7SNaATKpj+26LsY/ILAwgxPOPjTf+bWiw5aDQ+I8LBtm1Ll7okkUe
lLL4rsUG774DUTwpogOK1MI3lsCNlyol+cyjvA/eQvICh2x0wddiVdFZcL+DRiTm28S5Fi2htvk7
iWSTR4rbE3Ri6IW6SQumDj5eFM56FAWtfhRQXVYclxVZfeq0gEjqJi45YaiJEWeN+VhOfK+WVR+6
C6+/7Zgmi+JeN/T+kscXvHzFkay1Apc9rapi/QEtafw1XiTKOk99HujbCrrAH2Jhdm1oWTkbKLyT
fGhKSWZOVzoWsk6nco4ORkI8PZa1eW2KFOgbtKFju+wwANAYE09tSbaS6bdD87BaG0fDO/baksdM
yJQ30NqLW5+jCcs0B7uB2UNMQcEXEVYpm76MDhVGcgWKjWI80HSKE0uTk2UIm2w4CRo6rQLrOZAv
DVwqTHdXuRiySlQPs3gQwv6cYeXn5JHlC2DiK5sXlFFeR3/kF04pKndL/AAaAGgek4N7+nj6r18J
TNrh3IhKSAP2QzoSSMcYd2pPiY6CVnK0WhoQQdrYyAMK2cqE1t0wKbvfolhSM7PuxPtKJkGi0R4e
HWIWlSwUPKhc9JjLV2qrm46mOdkHig1hA7JKbOaX6LW0O3OCWlU9usFqyJS9suhlSalpbQS4RHRL
xxLSREtTpRbqEODsA3G3HV34Vmvs4wmvQw4J/pUHvEYfYmjkn3dNfABNpwuKdaqL/qKHMtNUDbBc
wUFKBATfwVexvi5AAnMjejy/YTn4NQm20mFUwU63jUkjDi2N3BVBhXa5xClJB889ypSqho26OyiW
Iwo/Gp0AoEf9UbE1uXchqEsPQlyQ2g+dLj8zwwwKXXmOsjFc+pO2YB7TKaTwTJ0Vxm44fROl+XKn
Wlopq12fMB5ZwiPENmC/ECqEzYj7azZtpIwDJKyilNWX3vE8AENPU7T4g1+nQXKFY9jaLLKhk/8J
MyaPSFrjtvEM2F1RhuhaI21QJEo1ho4UQt5rM/TXEneGocOXQpR3BgFAABdCjKez2/+VwED//8Zo
v9tu9cxzcsR7Cg4YuiYkMy1FzIN9l/1oDy+6gcUDJMYfBmKnzmYFPPHY0j84mExiRoUYYNt0mV3d
sOikIBnY4+PwIfK8XWh0DAfI8kj17Qy3MtuJUuDnqT6H9SeghKpAYqazNUBXHWvH3W+K6hAPqmBi
gpHNFDEhd8IWDZqZYWPG8wmB4VZ8LKBuM9dTYBntSdgTnJwrwIwIITZA8hkz/TNRXBKrq/ctvRwM
fPo3UhRtWKfQZ440t7c6C5xG42Zbhbd1y2Lf0aKKnsCT6Yqq/YcDhEQUU2J5ht9Dh0T47feE73Zy
ze4j2iXAna8APbBqtRjyLTjFW3CldPrC0mTxSDQuXnDbWbQVQBzkXz3tKpiF8wQvJuA+9yw0PyUY
Mde8LtqF6kBpLFWr3JY8N13YvuShYCwCWLjZoSqsQ1SsqYuGcOKFP77cB8cpVcQIcbCm2AhOx0va
kLJhvnthU08EmAdzAWxV5u0awzRuedr3gB+rRdYHqHy45WLpVrDadT8C7djP+qUbHHUORc8o/Ivj
mVu5BnCI4rbpamrik6vKv2xgf4b2WjnFAUmHn5PV8eBcn2ieaojpn188/0Wy0Zt0SgU476jWm+Zu
5Oq0VySQaOge3dJQeO6wA8qHsN8r/nmqKiAwqfd9y6tpRmU/jNFhfRgloeJubMoTwoef6KlT6Xn2
ZIIlkK//T+tfkk843r9GCFzKL3+7aHytjvLkhr/88V54bdZh3cb9iWD1qKYPEImGKNVNj9vHYpmr
ZKQmn+LAxuzP2LTwxQr0K3e9HUEFOLnFRgRY+N6xdg23MdVj/ELc1ywhaRFPOKL6vNvy9yBOwv4k
OwyPzSxio2/D98tY4AHoG0st+ZIDRJUKifmUl2vqPL9TlYgPixErXIbltFJt2KF3VPgBo5adR8iZ
5KAkJG02PkMyplhqeaxD/t69aIgLi79t7J9gNHYHGUrTF/vle2t62eq0nzOVjeeFN2Ehg7cKYGVT
2AVq8DEYQTE9olzr18cKWFPnj0FQb+iWPSYjGJ0petRKuc4M4dZMIylUey06QD5Bqlzq4Yk/hUNK
l5MheaNccsvN2YIGJBwxUZ1s60NUYmdvQYha662WiHGEB19aHHbFWFNCKAIvWmT1q1fvLD7FXgzN
Y3PzlRAkQyKvq7FAXTvd0W/QiVlEbXRso1UE32jAixUPWFoURWNNWBsV9NOWKx+8tcQJ74MS/UcB
1t9Lm4liWp8H05ImGIYIhTK/yWXKySsRn/SSP9uCStaQ870MOtPMCmhOGtbTzchCwy+SKDwBlURG
qqxHuj8LCAWFJt4pBb4Vkc2PoOc1wqIO5bqajTs8GHN42oZT8AxFrVcjQSNyNXOF34wkfpFbTxsb
9gIPQJR4QREwGCea0Ki/wGcLW1v9W4QQGoRrb96cDkkWNISJOuVymLAWep0/iUDRj1aBTDYtGOHk
KbtvQimnHsNDp3AAnR8ZJQSHYfl9SHqbq4SRI/tBzsGkgGQTKguZZo5OdlTQ/nzKTiYik+Hmu9Uw
/8SqSWnhyl7T2KHmPManFck1jQ0+LKnNzkmLdBWi++MbcAUd2HUIdCQ+3Zd7w6PJO3Xd/4HOabci
N8d7R1rlYpQOp2G49dCm0B5q7GCYC/MuMk9rb0YcAoKYZ7Qt1/Cs6INRJvUPYMZD06xUmBOPvX82
iE5ay+jidlkW4+qh0Ka/waJL49qU9XUkuK+LoqrCMyYionEFp+yUgrl1rD3UnDuZ+VXNQzwPEbxf
bPhJaf55rdL7eXcfY92/+z1z4SS84ZoRzX77JsCnMKA7TiYzG5Trnj6Pvi5hAetsO7r2/6rh6bFa
/qV9jqs/52+9vwGz5FwNVsnsfWjPPjgoCgzxcI4YPGVkB5RiwS5VRUdB2u+sYCXytrY+nhLaryCn
ZH31VkLS5cRxQNZyPf11XUq3AH9ViGM+Leu6WmnoGPp836BRcU35NIwJdZGcBR9iu+7Lz4yEs1Wh
81HqMYWlWDKrWjkEQdUPxB+EMs8Rpc4rGnnCC6WPyjlWQBPRFVzTTNHwsObZJJ+VAYosen7VGMro
HrS6hduvu1d6G2ETejPi5HT74bL7SESsBIeTb7MlFE7ip87pPHvbBczgxCScYf3m3C25J5n00s6s
NvpnkqYZWiHOU48VYAE/MoNTTq6QQNGg3u7gQp2Zkuy9ODFQBYkl1sMluvyOnhCGVcVKNOiSFS28
PLiT+HTY0LuxRldTQHjByvzdRA1sQRcNSwh0IRrlzMrq1ghaChCcCJCO9mcMYoSNcKFOGiOPcsg1
Bj3XYLgLsjcCbKBP5MiaGPvew3iKnw8l4sFSf6Nucx2T1vH0thgI8iF+gTB6UywHokBuqQUA5YaW
qj0iLNDyMJhqAWLGOHpdY1KHoULERLEqKLbeJYE0zwf2Uw+pQBnUL2uIzgx9n6k/JLmQNMKlavOp
ChsFfqtz0MRNll8/NJX1bXbBe0Ixx4Gzl5r/C7fOGZmFFNXRr53vZ+tJ7X/SmiTU+vjklpAvb7uR
WwiA9sqFJW11ESilxa9YiRyPKhqGsnPbbE+I7IIeP2ztylwjjZzUfd48P2ZJRdVvQVxk/WVepwIj
7k+Se6TpLDJOsBfk5RxafMRWvh9pRiLq5HaJsdHUc0O+n7sRXeICr5hb3km3FXAmJVt8U8nMF/sK
Tko8LYg+93Qg/tnKWwaJt4NJcCPxyyiW40heC/IplknLKL/yyj8SmxzkaTKWoDALHekuxkzV03RF
4zhUUFHV/jPKaRRbpKFkvRPZdU+N4BSKNkqNNBkZczUZelv5unTi6X+anyV5mLr23hIn+4uNHaoo
g9a+iLNPC1FyuHajbe9XqUUIQC7hnonvH/cGwggpE/xsLAeZjTSLiYTpAEKia1MiJgD4xrPV2/NU
np7jk8gk4P4F8t3rsQBNpPJxzW+YY9uUFN8qfps83rl5Zx2YK6VbfNagTQfsOq0PVEzozwg0D4GV
qCvP/vzqmltpXEZCSkm54XvMVM6NNJPAgZaRPS+mA7LKebqto7423lSiYAXv2Hve9UxCIB4k2Slq
oqEePDICJoqPbDF1FYHC8vXCS/fsnROQ/7CcRSRxdeI8TIBDUaS+CUPYyZkJU+VE2TrWiENVKoFu
CcR2iLYjaP6FJJNuMhb4vPuVE5ljGc7ABqqrv4ilbLqe179jOD3ZhwjPt6CPgGo25yKCy8HCLbyd
JfZZPW/4n1QpbvbabaY3x7Ci5s4Y0phNsJGtA4TS9scKkRkXEWyKW6TuOnaSlyBACQuoDDK56HKk
NxQn5Qw4izRgNClta8mlku1xBZc4pVl4RxH6NcLrfVaLADiGF1F0J6a5Lz8f0t0irR81Rol5Z2A5
IxtIWE5eIzB+35YsFCyGnkNXs45HwNLWdoU92ytuJXjcvRp3VpQrdBDrHmHfifYX1K8tBo/S97bn
6DGeLfXP/IkdI0OeTY0oAxonOk1kwkAzp6ygmyJypI/cqncANWtmO37BjC0/GeGftH7XdpuH7Cfe
1N4MM//I4FFgJU9b6UFnhCiNPl2uiPodrNSZ2NIFsAlj5ilCn1LSV2melWYlt/0yMSEVfhdmi/xd
RZ4SxiBp76YStifl9SymU9VgxkpSAZxaaX4V2lzEFpPVGy1c1F8sSORkyevvFjLHcvMK5lzRRwaG
N/BxRNGheLGdI2Ae4ZBaEqnbyh4d3UR4NTnG1RZGLdDNkaGXR+vECB4PzsXPCHQdZJBgFHeSMaQA
9SP1I7byEtVe9hqIKdNJG3kDOt8hdagvH+LvS/SEwijhtvRLqPv+VeZ9QSQu5dlnOP757cXLR9/5
L8UKytOcJviDVwvcCien991DspsxphEF2+NrrtfHMcm1wDsJ0yPa7xAJKaKq3jq1nA4akr0t1E17
9rNyWGZYrfa0mxqIeh9lsnOf/mCTnCOO5kfMYWlM7nb3BFPRIse592o9Fa4C4nW8rZFWX5I0Mw3t
kQwhV2HIGdWY0Km2eJeV+FT+nmGC826ES8inTur8prPFWgE1IIwj2db7lijcuDBEa+0X95aEINVY
joFzlxRBUp0WTudJvjTw7lER3E69h5j0ZvEuHrhhNPH4TvAJdsiGamKGkseNEOcjROk+0s/QI3nE
YRqBI60lqwgQ/NneMvo9I1MKA3jCcCqS76UrCtIBknMIRfbmF8XGgjBxpcyyD8drjRAmAH19zW5m
Oi9LCxaVJVYZN86RVTJFbKHY9WVXz7grq4hnWx7tH5l2hKGMmyx710GA52C7gO2ErkpQ6grUtvWi
IDUUA1rDopoigLAWNSjD3j8furLQqjaYg2jToN5Hk7bhAVC7Bg4i+EgxBVSAYsV1B7NxOcuCbEaA
FH4Xkxp9C84K1MkdcyVwaPV6dysbQRUPmYFLmCZUG6VaPq/9lG/jZVJq7V/CE0KRe/DBHKichqeY
JryWE2ZM9NzrIvOuW8T3pfDcj5cLKr0hEurfkT29mz1ALYh479g4vIAAMA5JD23bGuFSXjV7wU7k
4fwd5EhrNhlZPXMQ25mwoOH5YzIseUCjOh1l/BdzDVF50DFRk27F45uvI+02nnuCIVfeov4TPugr
hnOFKgHhrZyNR/hPaA93ldeB3LqyAaAS/bmU/wf4jBU9oYHxDn9pBxyNrkAXZlv3ClwyCcFjTQAy
U9m69N0zufUAQlCV106pvq5UzYHjBvuOyjnfp/z7jhUZivyRC/zF5tYLZY4sjn0x7CH8vCMIfcvY
YrqEpGhCJxIpMFZA70H+gW9KwLYaQXPKFOu6slRRMjFHnYIWBn8clpSp8+t9qZhVe17bOieu2Eq0
Y0OfO5b7BGVzsOV5QpVdnGjMf1NSEOLYIPjRQdLpEi9l7x+Znt6ratm+cNB7Nljq72SwYOjeLtG9
BsH1OhYelSz6hD04oki5x/jRVpKI7w7EG3/5tVN6p1x4kBFB08tyrK5xs1hNxbazBlMrKvjnmKxf
WYaj6dED1XLR3a4sudjUFnUGdpZXV1KxVVrYVrkykYf08w/w/JhLQhTIUE+27DpBVVes6Sv9By/P
79E5inswV4shn/Un5CZsfdfaRMWN+B/LwdYdfj/ZIZLL1w3GDN7beWAvIjJ9QPcyWPr82biUiya/
w4jKH7SlkDu2iLBM/iuRUunLtsVGVJ5vl+a/FSDGTqRzBuE0OqBp3bnCpBsx5tuHqGyfW4HhfSJa
kHO+BVVXqE+q6CObihnQG2SAoym6AG6jglR2G2Hcdf0bpMSgTEaPTItSEkWc2Q5yHL5U84bTujwl
oXu3YL3Whn3o5A2eyeFtijNY8ndNUzwMsD9vYmlU6UnYXS/lcA8r4zSNPWe9JhOtgpaWQwEIyWnZ
bbcz+9aUdbjV4IojW0GlJz1XzTtk9Z03cLlG1HNlDDRF8+aferghrQRZrTBQ1NQNEvw685pkIoj0
yzlezM2wnyD5fXxWe/uPR178LWAzkwwH9CX5cO+5vpZ+46pCK5+huzAAzK3PV7a0BBPgqYBHHrdR
DxaSAHEmVATqjRsMDB6KiMO8ii+vCczfXkGCBwd0p8syIrvh4P6GaalH5Mj+lWKTyxKtviPQdhm8
4Q/dVCciL7MKFTtCAdMIKB2aNvNcDW0txdMmM+xpn50w0SVNnF/vyg5EZLPR7jUfX/twikRBr346
D6zhklXZvOOMnHdwIUh6WHos5ERzMX2ufogg2efXUFieBeLcY+Ml2nKpz0WomvfEA7WSUDdauyW2
1TCCJM9Xr2I4Aw0C+dIMoVVjIPkoIxgVdEPIGYsLHsPPPzyj3govGdnfeD9PVO4gUsMRI/VwD/qT
EepHrppL+0BxQpz69ub3HXY9wwh/lTGxBxU1KFoobVnI9CUirvmPGx9DyD2ykzww0U4dGFnVs7HI
VzW8DZ2167vIm7XacmS5SBs+X/5G7LAMMQp7nzIJimUOk0q1QVIhBPA3Drgficpuo0kUknwPOVYd
9Q6JrayTA3YrxU22JwUw+ZihRs0gdv9REya30DdwvzQdtUhTaQKRJNvmm4cZHuK/oSO/Bj9TqeRg
5oBl0zyZSfWEcuM02/ULKSNX0Ng3txXUgKI36wNlpjqqBenI1++g4xMAr5bcpWMViZk0lm0aPaDm
LusA4Lifou6KDs6mjup/iDyH5GHnvXbOMlVeqkZY6sISzk2jDhfLlZ3FBtHtiFhzv7MnToTNq874
qOg1xf8Ib93Q//8EBY1vxSuG1qc4V4cVvfAvKtiB5yqjfBjNPB22R9SmTvzQENZhITH5KcIujd7l
8HEWXz+Y6z+mK3dYvx8h6SzlrYUuOmZ+E3J/0Fj0bOFPnLejTAUHEvsKbMypSZki8TRsVunzR+8E
DeuFtZgLociej6nOsd0AoJc8JRRt6JZ/5d1JOQk9BrseF1XgK5UzQY7x6M1KZ02ljbA8Vttl6hS2
+Zq5LOXvzXXImRDpFA8vqkO+ihseIq0G26Rg5LF4d4LghFlK0Z/qvRUBqSp1esirVNnoncQ/wbcE
uEYZLA152Bb8qIXAEVsaTF0ASKd7JPtkLNajS/GfB49PQKAD7BZ0JZmov26VlLYS3uRngqMjHsjH
eB4fOmS6ygr2KyXCkcbTjCVB9UA24UB0gd83foR5ZBEhDayQstvEN9d8fXFzf3ZG62vPZxaEPEuK
lXmAxfM9q0no+unmKAwaXa+7FKv7eLf+YNuaeWFzUMwKSDm/JU2euJJfLySGr8VJnP2K2ClUb21T
GnfXPzzERHdr2nzRtzdDKXT0Y5gGwigVfGhggdhrqGqjLYRp1ivMvyflbnRU21sdc+6aS2YZ5tsr
VDS1JpOb6dvEfLs/HF7Hy+jtyABHziGrxMivbLU7mj1eSmjuTSvJwQulvZ6+MViA7JhtE8IT8W05
SjwwDRPMblKr34cGIEM/BNO8c+Mt3jbkE6XFh9RlR4+LWEOK900uLRu8ngpv4I35seZuEAQP4GNv
bG3+YuFHAJkbROAbbiq3KA2OrkbsyUdUNUZfQKPi+5oTUbZGew/Bsm12Ym5BFR1cSmEEDC4sd5Np
vmSkr7LXdKcYTdw/OQW7VntkOGuIoIslqzB7perM70sQEOuJ/Q5IVCO3LyWdNuyYxdLZqXoooDtK
2gcLe0TXQtabBZGTQrLitUAuDABrSLD3mGV7j+GJ6hlXcfIWd9E4HWffbUpW3ZIdkIgmVH6Uz7Wd
Q+AfMQXD+KlY5/F3mpY+zZYZHGYcGjT7lryvHqbEtdo2B5WnEaMsOB78ojfkMu4BAjmg6Q9JqC/A
a8ioDuIq2TdB18bZx7TkoPhVzZAWDYP29hM7BgggpocRmF33P89SNkRFXhLdcZisDfQ9TfIu+pHb
4jEWritjpxwA5FXzM+z65iOmhmoieQk946L9bhbYQ8W2yMVwxy2cRKn+lpdc6XyqpzcqFJAkC5YQ
EJijoNFsy960g6N52tb6/k5CNWwRFCIfzjsANWSKMU7+r26mXy/iz7hMHqQo4rFVDSpHGH3mnXIs
RRSJBvFvy2/OP7laqIyc5hWoEKkdy20dEyWm0CFyw0tp4hALRP2ZjJZIu4Itn/NL8NUf++FVv5u4
Bva+mItiRQxdvYhafzHlw6Fa3t6wpgTvHOqbcyXvuhrpSoynDqNygY6X4y3i6tqviVFFkscisw3J
ESiwjLT7xejG/S5vbCfBsGDCPcWz1KLoPclmXJp8HUz+644p/f3pByKU4qw5Sh5PDLDZy5SFh4d1
kfvM+pZwJaxoQRJYhGkfXzoXQMqkw9hk8xnk2R6kSIZVETejR5FXHsnSL++KW3vYDIZiAIBP5nIo
QsdHeb61QAKjrcB2Ysa7saAAg1Wymi6MZcIosXiJ0G+GtiDGKws619tbwo3HtzihwNz+sHeOZ1ps
SoJJzBns/aHbCWLGwLFwcjpukN9TWl4wSfidGAb7MYdsOGs/NqulkmJY5MPdHjAG1U7qoP6/4f6T
w1hY3/HmpQlr5TCHmQDK3w2FyQSsjejBHgSMQx9d/jUBcWz+F4htxCHsvI1s3BwvCsrhJsMJy6Nq
MyufN6fzZ8r4KfAsDao6fHjBbG9DfJeNyc4Yjsqzm/ErRYy2hCPCAweX4vP+U45eIYQ+7pWbJRE8
YJ98h/TeW3kquJf9sDwTgGu4C91wmyvceJdSHQ2Ny6fCPCdj1sNlDQUKl831ikVKnXdWhpQa4KkY
VN8AZpKMEzhnVjwiwxlmuixFnhXcj6fbBD31SEJ4dmExsp9Uw0xS2mUhZoVKPESI4yZBymhEm4MM
Ous+dVEjz+kg76uerhEpKLIJ3FpQOXTAMQvGVCGcXqhBYz+xYTvMMTuqT+1MjTAStD40uggGBthI
r4bKVUa4dgTK/IrLxDuIk3sl7dwaOxPPmA7iNJVJ1xZQ0veHlFu5tRZuVJKp6AVgeWlj+ar8DFxj
S9l6VfqVixRymNPboYnFCoXvsQ6ErtyG1qbfXyNX+zqUKmfbzF/VYx+1nhm0JWD9gFrXOMmD9TG3
ggAtPzcYa3qVxOBEMG/d9N/rFmEQIUc6ybE2ZzVPLhQ0KAavktGz9M0WkSYNu2DIypKqSMRjVDHJ
04GRSNqFQymAGiqxcQw6c0lK/qZLTb2/SBFruBUJ/Kw2rYQ0KKUKOrCe2g707p3HPPX2dA+IIuj9
rWDD31CFJlDiHDFCVHAnyJ1sJhSaBUhO0qeAZZjJVgLS0hk697BMk9I9ZWYwrtqrkLKAszzlk0jX
I3l/11GCn71NScRio4W3INAao5usCyxEizx2tPUpPFOpCBNXHZe6jog+6G5S4mpdkgjSHJogPT7F
LgO8Vh0DhATIFeCUqnAui99bltZxl75sYH1JVupZ+8tlrCJR7Hn5AFqJO/TL3rGGG193A7sUiVLf
tWRbF2U1ZFVi8Qc5RNdMfx16w1qqgvApcJHTJX8Lh32huPkaWnDjIo7fxgle70M9vmvmSuPilmO0
tjljgzLqgzWbef4hn7fhImjQeSf1PDqRJ6hEMhG4DpigHwHecghNYavfPosKv2M88VgUxigd6sVc
C2gYoedx98ldTCrcQ73WgWGRuadvYDMhVH3xoqeER82wAbBGkX1Sr3zGekJQgpHI7MnndRr1B69Z
iJ3t1K4TW/Yr5qqFtP6TWqzBP2EZxsiuTXXLomD2a/ueuEt8wpTCgST/wblWGKtr7tIILQlJjk5v
+FlG0APP9LAenXjtXQxC4WIoFTaG1st44Fyqi/lN3Dzg9AF9dsOeTxhIl/zMXfWrR9LakpNx8gCm
XEy0UZ1Hpx2+zQjve4TSB+13fsPgI+l6e27pNGwt3LuivfbgOQiFkGvmF5Ct8e08G/hwkuUv4yCl
IUB/PkqaTMVkoupRf/mXeXTLLC9zo8fbeAG27oMijap1xKxnFscNAhoL6vTMOHZaS/+3clrjAdt1
WMtJg5Q7K9Rrlo05Askgp9ZXv2PpZm6hGkIbjFhfIKtr7tj/zH/Sy1rtd9RGpVHmMTm/jnvu/9i5
vQX1DNEYnBPbJGXp2ptun3iapU3N0upeS1esVoJvXsA+k+DYZPfzPCbVRKHRM7VA4k2M6lsJJOtm
kCWzJJnkdu9XrSGBOnrWePcAbmtbl+VHzUaMi14+LJnP/ZpzzI/hX9NNhU8w42gdYcvuAbwApGU1
BLGihcsNDVqSG6txJkU8OYhU3XM3gCtggnrwSWPFVgy8iSFY1HEdc0m+RHhkrq+o794G/kfTofNn
AVe790hftF++/CuRXwy2gnaXT+jRYsGi9FhZvO0q1Y1w82G/nPzaoYt+gn3i2AeUf0U66iCcipZv
8PFlx0B1YwwXGCHcQaWg0dAAgXJuLPvyUYQgf8sPkMdeMOyu1V2p/UilNKJ6fDUniQ2nAiSqZViO
3NVNhmOayMrLbjRBCCm35UaBCZyqVHv6LO/P6Xo3SBWnvR7qoRBaOsE1xX9WDfz5nNNv05k3ud7h
AWwIOByw8WdkT4TtZ53cJzHAe8xufu+QBuIvBheDWKOumpcqKnnKbpk5WzSc4pLYPKmg7AFrZC0z
vs89Is4a9et4M/8MZqRjid/H7y5e/DdQdqu0N0Oyf03/1/ldeIt9T8gkQQJt/8M/u08R/FyHapnj
AY2Fr7fDNGgslvZf8JgzSEEpSgyW2Xf1KEfxhzqkrlETsOvJQwt1SMwpAv0W9e7niC94sdnSKk5X
V6otwefZ06WjTznS4ak8ROUFAR0jRVmdQAVaBoYWwr124LFMTMbY24VO31Sv6s1WyCMRUItewu/k
8G03Wts6CBH+XEoR10kjKlYKQKXnyo7AjHyS+PDv772/6eEdFw4xApVpMCaV/CjN6QhpCr3eDhHT
U3EJ4cQuxykM7QlZwX27AQ1JpbiZHCJt1ka7F41y5bvgrz+jCE8aPAQ/IwL1Qde2QmiGuztMjStX
GOCoTNuMNLKMXiFxRY4r8Z65zhP2kpwzS5czg6y4NLotvQRQ/LU2SKId1bQSPsGBX8cvSio02MoG
z8dKXK9raA5rlHFO5p2svCkOxjRadxZwc6q8Nt2c/R6joTmGmgxug0BlbuWyj9pydAiCLwdtEgcJ
jf2QvA6qgXlHo9KrxqXhcKsbx43KZYoW191xOu3y4sJRHP4Zj7WWtSMh7tICncER7XgJJgUWg1RR
UO80KpKSy43waOkOKw1Xv210OC3wZZy3kFECw1R9RWqp8j7JfjgqTIV7H+aTK5vUFrzoagQV5oMj
JLxFgD1Zpbec4NeHeG+JK2xuv0xgmAxqDgLeLqmVKo+vHoKL804LFp+FKZkH8Pt313tvKD8mUgyW
ZvKP0cLCbbyU5CLkVU8UhfgpivTjpNGVKeB+i+Te01bsPTRQ+Dlo2dNYnPaVnHNB/h3Mr4BqPeiJ
9n5FMlwrFCwUy6MZ7KXzl74D7E6oqNaouqYsIV5y2KlLcT+jbfI09M0oUn2jxlahicAoE/xXtKiB
YQt84tcKOpT//cjhXYnmPIhenpNWL1nnr0Nuy7eI5Vi8w+GT2GsfQnQGerv/chLCYQwjSrjkCEpi
AvHpiQIwVM7i2QZuiy3ohFjyBMEEL2Cyw0Qn6sSderZ2NXzxoRKRxYP8nqrZILWJIBO234VotkDl
6U2L+68KckxiHgmVZmbrriE3186BEjPVnUI2ON9FhXvLTHQfR5n4RWqdOL5dA57NSSGz8iHw9RQe
6Ifl9CZq8DNE7NXH3UhzIDdPQIuHY+fcvfY4jnxUCu+fqsvjj/yVyl9wxeerexr4Gkv6lsozBqe+
jssxNiYOGhegPVEzDZMWRxhVcGG4zdN6r9GfmZ4KJG/1lITeY+o1CPWI5ik5xZbF1nkp6y4fDuHF
B0TPNRR5KkIyjPRPi2H4a5AV6xKST7JbdGD3VFW8K27r4mpjXxGQvibJtXQflaqM6vYlNk3zQRML
BCtkmnryeqJC//PX5fuwLwfTL7Ipp/zFVn4NKXfml9yjT+xUE5ky1B/2dCnAke3zu20E4tfr2Z7G
F9qweLHnoDXK0tebobbE2MOinMcM31RcJQ5Ccpi2FQYi8QMznMu3DnjxRblBvGtykZn3P+6WEFBU
RLhmuNo2nJfifCgPXxQfakfcLOgxI+qj97qQUh8Hk8J8DU4CTNfEiNJlSMEr7ZBWBUgWbsfDH0cl
FfL0QlFqHD627nr0ey/GdC6B86LU5JDM98r9fQuNtm2WwHHudp2lOrfF3Ry2+yJN5n5QEG5gkWO4
ekvO5sUO52n8EM5n9Y+Vt29XbWAdUUDrMQu3WA69GrUeLxgZopepH4/vU3vlshQBODkm8lzJ4VUA
o3EKx+qDI/F5IGFOTPX32QLjB+Gywr7H64GMaBj5Bl886lzTs1isMWIdct6uqV77YLSltmD/STp2
NaUV1nyduacAB33ViPL5iOgao8g9DulKzJUaOs+ikjU63t7ryVJJq6snsvJAC00cj2boL48M23Y/
jTmAZMMnUZUMyV8XUhtwlybkwzTNYCaO+IYoQ97uNWULPWnCNPChbJIRk1lSECT9vESSC4se/MH+
8rAUOBcGN55+o68C2mJUE1ukA4GLqtXoycfnWx9PF0hZpBk5PyaJSKpmxFKNXM8kVsKcAOnxjUHT
ENHuTZPg4HaJPWfc4Vi4yVCXcQ473l/gcXG69/7JAgOA4vdSK6cQW1yaKpuGoRU0sGXebylwWz9X
F3CaIJCz5T+S273p8nU3/ma2pyD0o2zpcyaBHwe+j02DrFhFwNAAkJot045KkqMJRYimkmh1t43P
yZ1yS4+LRGuzh+02MbJgrfW/96WVpA+uYWkrwDAfjDnZ5tXVmQl2WazCNHyyNfNdsGPCEe2b8JZ1
8o5W7z46aVVuVoRNLrMhbum2ZDxN0KiyQxhqWAZlbXGwoRrlButtE5RM+WjrTsZqSDGLVLoIFPyq
qC4bMAJb7EThDiNw9tCcSmsNr+pKp19Ew9+7KAg/6TRDNty7TN0nVOLJNCUZLHK9yyrx+iHWS5b7
HDXRPr3+8XXZa7/wir5E38SWq9JOwWvxhBKksSVpcE4pb1S5EK/f1hYI75YdOz9olobaopEN7iGn
uyZTQavW+RnNZwaQpRGQrgsLUKFjwL0Yoz3ZvmzGbtztGmBeLx3bAuK/4r5LZcq5xe9L9j8tL4RK
V6Kefsnyaoe1eEWHc+JciO4PtL6Y35nkOQI2+x01PppyZqCSyC0oswrceE0oYocluSQlDc6ujKuT
PBuDs+IDkKjrtvXypg8X5NXU4FZ8eCVS/VNGFSxqBRHoE2bk97Fi8RR1dzryrDmAted7zgT5pScB
AvlSjC5YcAWa8VaBZfyjVFB44OsEsuLAEZss032NIyvRk8tMrwl5wCAnPNkK4jXddOlY3n/MEl9B
SYqCu0Ywd8tzGLKvOUmOiCepPK3xYM8JK4i57wD6/cNJTFGghnZBSposzYi+rO8hV18UC70U/wCy
pCHXI1qn/px/DmuZoyUtcxn26h9w5wjtTIFJLb3fvg/x8d3tq92CVgeNtcMULcSrrF6EUTcQGtRG
rcebAr0WBCaciNYg9pc6l8Kyedjw4lTYHfW/Ivdt55AyE6DqA6Bcn1Unpqht+jMOABlss5dzeMhI
mWpm1TnvrUMp1Uqp97XSrpYwoYNBBwZSIfhDcU4tIauWAPa+urAo1YyiMCsybYthxo3bVxrRwZ9I
Zi0AFewsDZpf2s8R29YqnxAtEmuRTO3cNzShpzPWO6Uwq0+uK+dsUiCPnBN3kkcjrKSqQzo1+fbx
n2W0FzbLMxlDxxSazZyvmFfhBu1Ee15sirG+Vl11D5RMS/f1PE5i5qrCAE8KD4yi/Ik07gzaeYvm
u1f1r5btlKSCOxgkjKhzo1JgrpFZmFRgfGswdDhA3TSWTEDBwGrcFafeenQeRvM/2QxpO4bG5XPD
pcqnSHH7QJpI5T0BCIQ6zBtyxZM88wQ08i43089BfWIdnvBoXmhPRqEDUo8eM6RiislCo+Jpzb3k
h/ztxPndcEoaBMLrY+nUPGUv1nr4ifqQzEEb8exNuAN7QUk9KlkadsVRuojbEzDSnOgJHwgrcAK7
URv5X2HmwTbk2dyKNAhFPCiTQSWkn9gte6HY1KMkmCG5Dtr6egGTqC483E8sUmpbiewbY8fw63I2
H7IPJUbrK6HQoXzzCRXk5yWxT4PmDBP57XJb/E2iYYoRuWdZlnL3I0mE6+DmGnJKehjufkMSUW/x
WBozKna/b0nkn7Pa/uGC4cbYgBAJ0hzOaVZgeQXkrRt72+L/mEAxIJeFljZD5PIrHmTpvJ2Uq27V
r8IP11qiiLL2yaNhyphfYKnB97f695KBnOSFDWp/F+tSIcDbHrNj2OZgujdyGEK5+mkoIwJaMmhH
W4Qn4LE/4cNZCHflsXBBvc524Iefe50A9BV/JHA2FvMn72cgXLFsymD1j2zKonAVJfjeK0Ks26IU
sEKfghS2+izA11tMVYm5Tab0W9Iqr+LfFjPjCxq9ftoxHIE3XLIGqXyMEsHZT+aageFNcXF83gUQ
33IsNSpD2spUB6E49NSVsfrQCxLsx9cJyVvTank9al8nqWpE6pUwDYu/VCcq13Cw6E3nX1fR+37w
QzcnznKQdrJfyVB/CimyirXnQoV2u+W0bSDXEvxO3v/+SxI8+t6bQQAf5jF2JKLAjcEe2CsiiMG9
0XKvbTv9cRaUcm8IvUaaaBWAltgGmyzVHTh4IPoQTqqOq/M07LJKV2A6BksouIUWfaKLWv7WPEpE
NJnoZydhQ8Z0Ad+u+Jmn5x/+u6dqsH3qFckudTeLw1caSXy0eGvtUkz/Ck/R40pviWjqZTNxyxNG
V9yAU5+3ceyh1XoQxLvvLnDBZJ4Y2WZCt8jgmYR1hS/UnqPcEd/aAB0D4OmLjFtAJcAyxkWvvV9v
6l0UVz2Uq1TeptcIEwuo+RrhWB4p7crxHJC9pC3Fjf2ACVbTKlgeNg+aSyZpElsCwWsvvSiHAYED
KZ+1z5hrPRqsUhR8M+YTJqea/KoY7QfPaP58EglDGFgCrC8HISw9BOR4BlODCtd7D94zWVTdcVh1
bWLXu7npZBMOQAHgKttEhrX6+fUxyjcmTA3oOBCC+6pB+l7griYtVurXUmDauDKHixvD1rwOGw9o
k0aK5vdDpqU7ChFMlb8/pvULyKaDsDQ10PsApaNapxoAAYly95pypYQ9+9lJ1G4gRHdaJeg3+NV9
sXEmjlv2nQJth6+maDHzs4aKSiuLfKgH1m3WXCj09WUrW3N8YL2sMkAJgrf/srAsS8H2NFqqnZyZ
EfCk9lUXIz5l9ovwA9wdNV4L62Yltwjj73QVyFlNxwBTTPqC/0FYJcDWtjNGBRBFyo5MiAOyofpP
lZOP0rzouassGn1qp4KsxY+XVJdSvZr0a+vbgo0HUyNvCnfoX6OiAbgkf9zBMW1L1s3lrd0f4d2e
Z3Y+tOoDLvW0tbvWPzO32SH5jpQ0i9h0YorehGnHV3rwyYUmpfdU/fE1fzfITzpK31AstUipNTOe
uGdD+10GRWKKf/rm6UpSpDQ3cc61CLyGkiBW8g7tSzuxd9MV/Q9YE6HVZgSsWkLlhiAor/nKOeN1
OLmwJQJ/lmpffSEFMgQFoKR/yvJdcJZJnipop/Pwr2WNQnFJMBOL75EB8R5qV2BUw/486rslhVxK
iDuHKuktvtmoRC+CCqsYfa23dXEuR9uPXbBmZiCUhRfwTU2Dm+AA6HXLSWPnWkhmpMRopUvvJEGj
CnglZjxkb15MgEJr0kotCJQJdMH8KzWDjcTzLP7xAWscSqlrRai+8R44k8gur2wnORLvTncXrbEM
gw7Frgy+eAJXhlNp5ohVma3OnFGjFABHG5ElkrlcaNJPLqaMV1KjfQDuHQ6hKQllhZHuQkuR1Eou
fse58e9aslMd3GkgjoYAdBvtDNV3MOgBkf2sf3jk9NHHi54TLcxbLFrMnTA5aSv3EpFe2qWAOY1l
+jbbwJdfQprowjPNN35G7LeuIBcnvLAjTq9HE2hE4mYZ90B94qNDzB7HiVMXGqaWPOzdEnI+znAz
gzitW7bfedPv1pyf/pLBL0xb316Ywgfsk+d54o8V3pu3V82q0ZKumf2DNJEfhrmwXslZr/HLduP4
idK56AawwGXpdNhd3+iJ8kC7HLN9QxQNSSyoxCDiauNdujFwS6gjh+OuPVWlrImd/kpOuyyz00VX
3f+xojDF5zETFegOFNbHQ0/oCcB2OZGzSS66RlfZ+As5y9B1tGX11nvWmRbJ4HbIT8aLw4ihsDub
iVRjnQNgw6WHCaXFuOJWM3jwd/RerUSi3icH+PaOYHxNBgcDHJzYfEBuHJKHWRJqIl7venkSPNnm
BzDHoE9lFSe9VI9+375OKLafQ4wiOnUcTyQ2DcmtGIlrOFGRYAuaNTpVPcsl4BWmXxyZX4ebyZhO
85dFoeRpXQvNmImqf1tV+3qcXgqS6WHoPT1YKpuQdsc8QfDLNH0KNzMz0S+Isb0ZmriIjK0HxaN0
mgwZBRBmNv7Jim2TzN/QBLpIw3ZA62t9Y0WZNlJr5UBltjkJ6e1H6nRGBzfnN0l5FkEyR+10Eyum
nK9qNXDEGdqPX3b0OjgGgZ7OpKVPyRNxXKBxdEY3f3mirg/Fxh30kU6gJTNhYGqEhQ5XbacOBrFV
o9o/6UPowxMddhq1vmfGcPOQJ/YDaW0YCqq4nMypd9ka63zfJLrfvPif7kNDcCOVCbF1+lGBLAzS
tyRRTZuMZJ0qCxEGTu2snDnMqZYZ/HWuefpc9XMsPSDpgaY+3HTlDnD6MD6UgmUPQE1EXyGYRXAu
JSzNOwcGlKgFlR8/ffPjzCHnQhRjFVtIf6zSPLEqFVAE9sxOdUhCRcBd9PPMj/wgmHzKQHmYH/yO
UWK4BHUl7RveDYqQgFvOQKnf8OE3TlLlLjcTLMoRkatkhvgh/2ew4lh4JpYj6X2I9+3Pyg1irpve
hcJtzu4CS14Wp2jjDtqDGA5ze59SxcYPOl2D1mys+vTKETB4iBNYBgvrCW/m5MsQDFi2vfPe7BV8
enMyuh9PczSVlAgwXSFsFDT4Zi9zYIArOkuaJN/hslJohWqIncA3C00ugHIpc/isGGxJK8Sgtns1
bLsw9CY6LxEHxinaviX8OJXG7Wfsqrxq1Elp5rlxtStn3A9C7OIKvo0mZ0h7XoLk0n279C02XDRj
BbDm4Pad5njA5kUk4AHo7unZINhT2CZ0fR+oKo/jGwHPTVZTd40r1fF9sF7gbRQWgiIh0yosXAZX
vF4wzn5ddM8MZhBb51lI3OI4zMPZQNdcmYfk4unFfmLzKm5k1v7mJAj5grXLIo4iF4+62ovFzoQo
DdylYl1LvKxtByYa6oDOyga/a8Sy9O1W+ufUVuPs4OlOdTdX7W+ECziqRMyKtEQRfep15tIFDgB9
yPKGa4Q7cYReuGvQoL7bA7Tg6mH1GDP36iV+LNITrmH9Wv8qQY4btAz13Swmuu8JdEQKxdGAWXL2
xRa9H02/hPLLmpog4/bRLTeNyT/nd0DpsYX+fYlAU39qBn+6sFetP0TIX8RWOpZ79j9LpKRGPlcB
qKcbuvQqGMog7oqG1x0i4Vyq1XrISQ1KlYUxyfdfxzRmXhwBNApSxZsY5aO73gRCI3Wmog965EC9
HwgCrgAbEHkBxNIphVgpmG5+L0fXLhJc/e+GEXe2YTtYhoXuRFWvFJfoFp6F4bMh8XrTVMNUMOP+
CJwSaJwmgl8nj+jtpnlsOws1r9/QbFgt9YmZmNuu/DnYbpl8UDtM1OEvn1+3oxjaT/gpJCNYXHcX
rsWvK5RAW36mlL0q6DgJYIm6pFjfF5ZwNS3Y4XdkoHx+cu72HfrTofD9wenf8GuT8s7nFZZBPpP0
X5ClLawbpTSmHSpIIFRnbWwCJp5xIxTkfRtRM5VwEoyfluUWeWn/Q4FpuPpFD1BNX+33t/dQ+B5L
8GeiakdNqHQ7be7Ikb9KeAfJq9WUgsyG3T8T68u4jLuRxpDBZxl074/4KXPk3Po0bLq8Jbjdpz1p
KSG/RbLzwol2aqnexrHow2EQJTKEcsy/uuTuQDZe3gLm1NRDoTGbgI9l+UauQdhktAqlQmnfruJg
BCpKcB3z+taWM+TMkd7gxGIERKb2VowSrCDXKaIwSqoe85Kl6sTOu0GnuNyyGxCD9CryvMWfRUlY
aUyMvIaARC6FcZdkABsk0ItCRiT6b40KwGt6fbowVixvPmMVxSs747JGULmLD+SV+LyUqTLbNiX0
LXdFh19b2sSlCA+Bmlc4lcdMqd4bj4CMw85I3eIqk5MyhzkObFerZkM9JovoKyPDFGrojZ7HpCIK
PirWHZ9rolgWr8u+8UDgAJfqwTK7wIGsEsSVDOa/iHqebVdPEzFuL6ywz+c2SMZu0mdqqPmVQWCl
xwGzTS7WNKsogQaKgjsevJkaMzd1cVJBotwz8IuRUnaFG0ggMrkJSmBq6V4aqoP28bFZZYGeeD2Z
ou8h6LMBwy/41VuUvD8u6CqSIJT6G64JfKWCSw9RFByPfwIsENT7I7yeQOBXDcsiu3cgWGKE+SOY
XDpp41sCbc9MW8QJlOlUI5Bt1EBEWcE6oc+fobCIatrVeeBW7H3gLdXUwg5bEnTnB/H9SEzuLHvi
nZAp6DINW7A1lrk6nZlFKzUuXlRkgXATLwwJQcZmznrmJr3tR2LJwWDGs7PU2LSikRddIv1RQPWL
zJdAv524ffTozZl+EOpMkhPu8Xfei24Hq1JPzV9pqvkRY+3E1MukUvPZg0JhRIevQYI8JHXwed2X
Gj1QRVuIpQxYCvBS+4Mqbg+fUdsxfT5VLxZDd00f0er/dssD4q6I3g/pLwJ5z8+1JoX2eD8pq7Eu
RVxrewRQSnZC5KyO7re1B3CIk1wR3x45KmTXxJ3dLlXv4tTz4BaDvfiz6nWpak6okbQhGL0nvapL
FdTw85qspEqrUdnkXXXwjGtS8xcZpww6zAF8+oLcDvupScT1VkPztl7guzhEC9neomWI0Cyl+Rex
rCSHAOscfuIddsY1lfhSNwfpPQYRBJyBJ6y8j+sSryaWo1gdlewg0MY7IpgBbQsiiQCAUk54xMmZ
W64q66bjkzR8T0t/0U49zUXoYy+ImLYhfTk6hmuxrbdd70x9K59ArwKjF/OYjWOusRhC4bCuIl1P
LHbOWe/7VO+QwUX7tZ9sECAlKTtEUu8yLN52IUvEtQqvx3PHSjVKAZLopCBDCQs69VIxeBjQt9+3
o9tz8wWGYnCQtaYcJybzfrYJnde1Xvc3TFqRFyQADrIiC4rg+EeH9cjSCiBB2fl6LkPE6p+GTQIP
IMoQtpOZ0FpXqbEOmfIMR1oLrfeJIcL39o0B5N4cD8J80MsRzHYTkGKFAc+l9hghcXrh4vCbah5h
CH5W8WvC1kyJ+4YQfNNt9vX8j+XKnxxBJihgn1h1zMAIgEdBhBQ1PObCME8ftWtRUip5nsyYHXho
wIiMNTwi1MV0vCXV94JOzde8pfzttMSuY1bu813rb/feeK9J13b0PVvUWY0ij5DeK4sEBU86f6XO
sqWmy2k9wdoWGh0FYMILqUVAIsTl5NRR8EF2/HO+AeuNXXzpQAP4kI6cfHAzQDJ4BSkv6PfU+Ozn
+VyjJjHip+bLubBYOWDSBHAOyK/U8k8J4e5p/JeltDkfQqVFQsgCEwy/mtQ4bMSV7iAezpmlpWhj
r4JHUSII3EA3bmO45stzGfWQD3YUu9VfPeCm5KcGV3xDV5kHwzLz89V2vl52XWbzqK4EAs6eR1WU
ueZ5IrvXbJC5YOrFhnARwMOjsYyaLyUCnwV7Dn2D3L/S78kkO33iqyPBMdh1Oe+QtDL+rEdFbsf6
JepjoqQmaWgTMEUvdepQobqCoUIuErpyEjYwdg34IDrhHZKhAUh1Q18vsr2RwdHrjSl9hRJIheJh
nJ4mqaAS379BOawE+5Nd8upN/LmevyMU2xTuvrfms/jbGFa1AiytKqM3DEDUbq0c/b87E9xXA7fa
Tu16l9XifHNMPZajjzTRK4ZQg+zO/6IxTwygHNf72ZSBGOhCLYtW4fVb8WAkP4gaKB0f3z8eniwS
K1GzY7zXPPmlCGSvqZANGJUJVLoQr1Bsdf8Pu4Z2MuioE1cuIwiJUxTKiVYsrW0VypL6UXQWemzu
86IPQ2rb3nOU3gMCvaiJIJbcBMEqCnPWmTO14OjROxP7qKdfnuUIT5sxHOI+7yEZQpLPlDkTn073
/CiA/zDJn0RyE6FATZB53vIOFAzCqpD9NJXT/HoBrDZu52AqInC9BM80wBCXgARbBcDa4j6AOUmm
wtJDYcke7t5ZGF/UKX+aXn1XK9+0quUTGVVxgMdP8JQu0q6Tgx6y/fjd6WMEW2Wj4Q/oMQH3+zDm
L/DUsBhfQE3bGVIIjYVUcNr8BN6wQbntm/ZLwTbdVL+BA4Od2NYHCeHlUw2zcNccQDMjf7MRxyR3
gwdj1tfoRI/N2K3WzI7O6fOOuyzypxx5lsqAghy/BVmunnw6i7aMo2CDjKo+2T8k9V1GxiL2+UAa
91MKR/v22LgA5C9taFtxGGelpVG2M65HSnWEDbtVEKavHFuSn3zMLM89a6MKetLoFDK1AXYrPkw8
EBLr+fQDC5YO+P79nIZ9WaRnGAWBbjzgAfY6NHdbv01FWdzdWEINcSuX5RS8QwrfZFHcbRAQCwOf
vo+Q6kgLBE+D111wzcpq2k6mI0A61XRno4T1aqQxHzoxIFXT8qb8Wnh29Y+T5hqMAp4EoRmMjTlT
4YeR5KumZ8XSL+sUHIIeTlnKPvYU9cV31DQp7j8nmZUkoRIA46A7dQTxg0IJJy5hz9H83XMcD2y3
5FrNzW863LP105ByB/XWUegpRoq8yisj66si09px6ZLR5Hjm1MDHVNhKw0Yns+S06SAzflZBm64R
9Ip0Mr4M7ifix1UNcB9dDn2LunV5+z2lxZ03jje6dyh/NVviV4Xl6WwbOOoz+gxt4ECfkHkTVTF2
ZJo2xU10CzGQ6pk80s1orXnIeEWhQYcHNdwxwGV2Kvr4DtxJ6npyuIvbhw2Ud1AczZONUPrGFkrL
beB20sJiOrPmDORoJvGbnPWd/GeuGWCI+4qdsVuqgIVLV+I/d34Zs+d1gKDsJzGg4DpIWesF/fuL
UB29POzD+gLgqXjByXn0Pn/9YmaYXhMJqSfMk56H8AiAbFpgy4EURR26hhm0tw8UctpSnEWCuwcJ
fNiJ+yHuz6kyDvn5aBJfH3xacJpke8hVA4RPhpom7zPEvcRosyN5RjbjdGlM7Af6wro9r08A4a83
0r59/WXhhevPJU3BI6UaTN0GAUnQ6YkphSdULIAFktbzW0nTwpXGI2bTQRdpNvEFcttqn2qbmKAP
LXSc2oNmhliB/ydp1bwi+NRw/iHgoAXk/qcgZXaaqJs+X1xBSgYi+ZOecnNEJm9DOqft3EPtkWUN
NwBbEIK1juHxhwaO+xDgtc7o97Tu0GG66tqzhanySqyvfWcxvQMY4LaWmCC+OaIlV/pdUIPK/u/4
QXGzK+3Z6+61wiJ/J/UB+ij+M6so+gfX9n5KwKr3ZHzNGpacwfaj+iR2sxhn9MUVyhX09KHSfsJw
buc+/V9IO3kMFBBuRnyDg7LhJ0lT9g8rGvgv+zIvguO7rcTdfgafo+6hlzYxUANDm3HG63jBOLUA
ubmP8jaFvcZutRrtHiO4onF0t3PTuS1bIUe8gSG4TRK/HhNY7xjcHh8tv/tmp6fcKorJ+uYdIOwy
zd4MpRGQNKcktdmi81jApD4m76Sa920L4OtbftLjDNYlrb7ez7WfgyJDZpO8rxUKNOwqUC9PVYYy
sf5lY/T74XjlehNMrvtpqyKW3MyG4bVAqLLqKXmkYtsa2zj1WjQuP9WdJpT7UcOixpUF99EHL2us
p9hzr93QAlfF9+hT6mLLwahPSJb/oICDFj/68FUHe6xQ5nYqFCTPcVrV52eg4hnP8BgZgPCvvQk+
CPscCKrOG4GFmooyHY1SSbQzIGyZe3OViv5cxF6a4mQox4KLh5u8obRb8tVCOagqhCd1/kJNaX4I
AXLQXrDMcuZ0JerPOVd7WUj/0QD9pFl+reh3kGBqrWY1h8ZfYBfBf1UrGCo13HcP0qlzndMZ0RAy
hB2+cRqY3KBUqemqV+7Ew1M6O3SCg6K/2FMmfdrUFxXmD+JeJg95ePexSwELhOXg9C9hDVJRLhgl
YugWNX6s2e83aLnoGp7L0XoRNy1+sP2lY6kPnxdfJTH0K5CmTgjwpiBG7MY3He4i+T+fgryXdnoj
vdizOTsKGuCsHFXgXq3bgwk02l40mdFVJQEj6RAj9YFEaKwSIMdjmVhAtiesNABZt+mI35kywN7f
/kCzvEq7mLK28RhNN3b8owFnU4mHbSNdMVNDUzmUocDSQW7jObWMxrK6ShZwnxtjp455OiMI3ufm
XDb5zb2ja2dDAAphnUmCCjFDXFjIoVPX1gpFRpLf512Mpm2PUymv+EQoqsJfIYvOqV7EBJaEK6Uf
YGNrnZwhQ9e1jcDegLNAV84GVbjZX+n9pID+gSG60sa9Q14Yui8YCNzdNbVa5vuzlA9NCN2f8I86
ssXlB0M3lA5mY3/6BrRUadmkIONmk12UlUngWkee/jk0CU+NkjcxGpr9+5zNL0xAeND280jqma7w
KCWWt6j9q+jPRXIUY6ut7GNU+f/KowQezBuyYOCPaQzhZ4K1wPP+Jzql+pxWuKyDbXmMingUeU1p
XDhEWwUUUjOWyRDqxcyVilvvzSJmUnkadayllJmRe9Q0H7us82LCN+QjfDJL3J6uwSzIbPi8m4/f
nrMEuFQHBdZ/Rrkmm0ic68Z44VJEVaCQRXRodKMWxR6SCI7JpymjiXq16HL88FoYnFxLDdsTiXlI
EnbdOiQDCwOA8sdleD2unG8fZpC2H7K5f4BeLa/AtrHLBANAasrpdytygTAz0aLYMFuw8ZMfE1mJ
DG2SJvcnmrZmu6PX/J2oXa/O+xk6Dj8T6qCMIj1z9cfjfpz1i9fRmpWN2LHd1CxrjvQLi6ZzzzfU
RCVf+0i3N4SXYrO+i0OERG/3CsBDFUxSFLvtK82xmDDWZ2LKAHLilcceMrvjQO2ASKRD/9zms0Tq
SxddgtWtQCemnoKrFEd+pT9o9EPciUFeRoib2WKAteaK0dvNa/W6z9zH0A/A0dLURDzK/uA5ZHa2
9cqPUYTOGMll6YYZTHYaZ3DCja1uNHce4Xf0UgKVCDpNYefK4cwcGKF46QLs9HXciY6jIUrF9AYD
IkJ0CDONZQlN1w9D6S4qh4fXjCKKcXyB9UsZ9YQRIZPuNVbGY5UD13vNgwDSkeqOR8yND9cFkDvb
nA1sEb/6PZi189RmFSKNQwB0dSOZD5/AE6rwjURixHHpVZwucmPQX7W/9Z5W/QedTwyYvGO9Taug
8KGZxIzEpbLssGRIIzA51Cl2jtqFYDxBIirGe92rshYnmbUeL0apmQsGSyxQJiIOprfqbRs95iEg
WhFY3X+UOrp50Faa8sLK2zx40Ym9h0eE+iOqhGF4XLLgiqP8zXreTFxyYpVfuVk131GcWVOFokSq
IJEAqXIW4q4sNhMcnbIWDD2gX0++iYw5b4mH6gIbkNyW13CHCjLMtzNjKP/oFLZvjJHLParM7tYA
G9gr/SxOmWCGLgcGhtbw6wBLyLmZwYIOx+QyolrryXfvQENPHfBiLk6OJySiPSvnv60tCdgYAKY3
QgvvXH2dtxi0sR0SHPrWFOSd9QIObWFm5BITp9Imx59a4Rlc1AxeDbiHErpETxT4gGzyicznWG5n
deGe6yeiQ7rPxe9WM3TFgo5g8WuNNhYwKxGloDgDhomCnB8VFUg5Enm90XLaaSdEXQYIZvxWLZmS
VV0/X/oyzJqZZk6U2Eaqyy131EdetfKR+VQONOvUPUxwX72+S1Pii8b/2sq0iZVmBHW6Q2JLI2RQ
3ityzKOdtFshbrhEHaYlrTM5PoDjA+KtCJDD1BdXUmuVtmqgEo7O5SiiBkVIRS4gc7SSrbpEWgaA
MCKCtGqEpnhyCGdtzxFuIoDCIJykoKu/XwaD3VY4rMNjzW9tJxGLhyflI4iRprPri5RxrttU5veo
KG89CaopqaGkpsU0nJ2V+QiRmQ3GjWU5XfAb70fNt2OOBHv1PqjoGUf6o2mDrzK6170YV9JhDDmI
o8VmiEIZ5g61SmflSVFCed0NpSPplKH8z086JhXPqfY7j2JH9xwRS8hLCv/ncyPX04mAUWt3PgSJ
m/K8jeM+ZWfgpwnMkMSBWVjjhwXumSvOKZpA5niSMPjJMRMPI/J2G0z4338zWTEKEcEsj9etD24t
BtOlaeutVlg53x1sDckHTn+XxJxwJa7Ei966TksIrff0VFky9ZL4qeB8MwX/dzOCMrdOH0dZhT1j
ST/+L3A7ew6Se3HyT8F4w+ZJ2F3sj6bVGyNTqEiXZHSOOJo7QvN20pr/oBbdvLN3+qTpmmm33wQe
95+kWYMgLkqXUVIfNTj++jOWKtYoEjCYh965sQXaZBIoLGshK78TRMVYrlckgolRoyP+N/Ioakna
nhf+WY2wo423Kb8mp3pWnomwyNvmHwSdUJcxGNSaBf48s5Nl20WonREEqxlFJfexOOHiJNHI2DBh
S0tu2nr8LCkZu2HsFLQ1gxDgDxcuBldKKZ9RlB4NRoJXs60nk9IxbLXWqulT2J81bccHLaMTCDNH
MHeadXD6VH5U24gE05GCXF1SydIVmq6LZJMytF5rv+c9yMUaRnJCs7TBQPdJtd6Jk6Wcrdp5pQpY
GY8eyiF9TmXfk2/0LdRAJrya/dL+wWwgI+DLah/QnJFk+0t+Mly6Mr9ckTlDXSIVYTHNU0/XXW6v
ZD0B42vjPvFq9uozi1eZDj/JVgBslat12Mf7EhDRQRudyfjo/tpgyYUzbbQubN6ZDVL8Cz7RWev4
xcu5N8PqGMChmdBSMA4jCU6JjlDEoNGIcFnfHrFtfda+chFp+BsAhCwCBWg7LRAeUMpekACBMIlt
tlwMAjNUO1qopawTpMpICKrXIep1NMs0yMguCX/PYSlJYoZr3/2WHqw/6yvuLAxIA5TaUgi7ltxM
zWanYYYh+AfGJXE95zAwyrABBxj+R8NM2gIEQ1CLPYdRDIVduJ26l8dBLbqFsbCU+9XKDhsKNOUr
PlkQrKzezuyFp2WbCgk00ETOQXow4rLL9Z119vrC7Ozw+wJIokuFq269oN0M9Wh85O+FUB1pmFq6
8wynDos5BncQsUzfEWGtNaYqYTJ/XDYyoH4R65nNFzqgLMSqzSAdox3eFH8rO8SCbYeN7zOXPczB
vTzpMuGOonu4J59VK3dAorto5PPovBu+4KIe5Q0g+pb7PtyRCKhotbdq1L7LWNlb+sWwg23/UvTj
5fTlJKm6Phwfx2T/Z80XJC0emGm5YLf+YSE881sIfMGijy+L0oIALsX4uJN3bCBl3YE05ESx+xdv
CwNpstXKH2mWT2LIZxgtN/yxtttNUJgGCkzAQ4AR6Owo2JlXqLNMl6lWQfP9opnGJVCcLL6lnDLd
1kjyeFo1wIOTL2ejbgPnTv57MQ0IyJvcStJymip1agJDu5IfPoTqxd4Bmhtq1430ZlCz8h9VXRgg
MBnaKXrUCnAcW4oGPEfX7I9WK4+mzP8bQIX/cyR4BK6hT6z1jd8KSUP5BHHv6a2ZlIEbN66Saha1
HksRh9Pq3+803+ncj6p44a0Vq6ywEPiqpMclHRlPYI8q/lB41fl73GQc/EItfYpdO7VkxVEOR6TV
VG1l1GjTerl99UwHKUrTyQ7jT2dd8tNYNInEhW5LV3EfsjfSncBn4Qhb/OnIvKEGxUNTrdEGPTWV
J7tw0ml4C/j5LcZL3x0kpGVqnNksOPKrf+OSmKqpbrsFwc3kUPgG9Q/yaKAZ8hpaYVRsrgtth/2w
Gm2uel2RqOebU4qHCtCbMGXaDWZvX4Kou15BOHxYSoR/Ts7Wd74VWOdNDKWk3hid1oTMCX+oSZch
y1i/s4kb/45Rk+xNuMrs6Bvtg0Y46gXHvFR+RfxHLsuOKuMHFgUs4PI2NIBd0NKVkNwMWZTDr5os
ntz4HFbuANGgakv5/AOgMLDEx/zurtaL+tj0F5fgw71zevk8IZrpnZB3mYSBG6mz3UfEyQWs+h6j
/0hh99mn722X6MDPcpDxOfRYSqk+bE+yWFEUqcUXlCxD/8vIplB5PfpY8mklbZVzZbKFqSdxV5Cf
GSMON783KqGhCceFc7q97/ppLZ4b5K410OOxfegQZLI50tAusGPd8MacBGOFyZQPLgq1Sksk7nCO
ORDznBXT9TOThKh5jePuRXTUOyYRGecv/z0wPzGsRlfw9EQc93tS4soGFFGfMm8oj437253046Dq
zMXGNGJWvMrEoAMofBYOUChkPxEkc+HNmfM3tJRPVaMIdWh75m941cgP+eZmdHbDBrYQhpWkLsqx
nip+OMDc8x+sOv/7rbobDlZnzHIZKlSi1O26sdcASfbGt402oiZBbn8rIxtCxbcTEN1wQbIOvsiZ
UsK/0Qp+jO4vYv6BHKHUl6aZWyQK7V1g9ADfvzM3nkxAJHOvwbUIiZg+HGHdXsWgE+lUzQP6xG55
DqtCqumvOWdVIzrMI76rHWBlIWWfFe0Bb7YPHD3gvdUipqXO67/D0wYykMd1NpMY6iIPV5W7UE8x
gggE3wh4XvjoItPRbhTCB+i+kS9K8KD9kuJ+TWHH1BpYuKPqvjqHWjOcmmH9C2FBkG2xjY1pFX8x
WxBzy8E5+h9fhIN3JSDTaS9iSaap8JGny8ixV5PBhJgzNwZIiFjy1Js/KlXFwHc/U8P6mGxAlfr+
+jhirQI7d5zSD6uJZwwnwEcuRr9CeUbal/vCBx0q7gFDyeVDTMoCa4TRfNYU+kiN/0eZV157kJ36
G31nL69+EwGsEzJ0BQMDER7knYvKhURL5IzSWiP+sZoa3vZEcW86J86sSVymykyKJqC8ukzCNcvi
yoYmQJckxCFQYRaN0X1hKUXOPmF9VTZLEv+Za+AMXvROZgh87AbjDMWGKAxf8HBDnVo2rpimAQLA
Vh4Ycr+qMdSpdpayfc5f5Gzr1OJCSz0q9hyqSh+d6hbS4H5vlILUvHB0xqS29KccyeaFgdrH8Oii
TjaB8TfMth3GZJ2f/AO/DSrdbAGMol4jVhV5s2jBC1iR//dIF8PxUydAWK5pgz+YnUEAwq++GaN5
8LM7OkYhLJAI1F4hSWk9Cn1M5eoefpopRlFqOC5+ltXj6eQrm2MJVHcyif5h4mjVoW0ROcl8BfwI
Lvaf2s9HOndaJu9R42imDug144JvxkfxvjY+GuDsQtht+5MSgBj8CcK09tqfk8A8hujeNb+Qp20Y
tM4IzLe1jzkLOoVyxXCZds69b9QkffO2JNtsOxxTVGLRXP9x2v1wC+3btuIXMXprwK+vXcq9aUkR
iZjGRfOM3KCipCB60qA7ATj2v/RG2MZJGLariwjE9lqRkAxm2GSAMEzqX+erVt4nb/nbWm2wLyg3
kmBXL3EigcIcxaIwHMWAUDQG661meS/YZ3lTS4e0h5fgMGiXK/C+rMXqI7qUOWM1j413WVWB8WnR
vFrpxy4jpDZgb3hOrjXpwuf4LUHX0bvbbcLTCuEbOOl2XC7iE23UvFLKDfyhuE9wXW3UULyd7zbB
A+F+o2/9g0D/exx9LJy/GimGoik308bK+mdcvcEnU8MPz/GipeQ8jUEsm/hu6jonBHxJEkMKAZpY
zTE1vVhF1DR49ZACjG6QMzptrc49O14ROgJNo4dccMRWDB411WVB/WEIzKS+yxGhqh9PzM3h3K2G
f6FkOy0H4d5MFz4qBd+4emGc6QoWy0XYzbVECOFlM6+m+H+b8ljeWscx1ycfyZ2Es4GaByqjiql1
+tsGkzNd0RJn6Xem/eMMAJJnhLoZN8aj7czz+XvJPIAhZU5QQg7PgDM55FWA5j4JyzpdPEBtvQRF
X98GtGX5Uedfu29Usj3qdiD1juDnGNDn43QGAjKBrCGbsDic/6BY7EMGo0JJ6pndputd7j6d9yGG
vQc8GgPY5CmwdiHoVo6z5Etg9RCWfyNJ2ZYJ2MKyfdiZ7oAS4Jp/weE6I/U3leDCH7cnMVIYzFXF
bQG4+SeGY8hgZgemxAFoLCL8b2uQoEoU16eMffPMyyYIt6CnSLXMorCOZDFQWg5SBPdsNQqkfHHL
JmK8iyQ4rMaRlq5a9/KSgWPGOlMBQCAbQvxSZqXhWrTjjOQZy6OyAxSI7xmm/Tykk2Pr95grbYTQ
9xbP8ndfvE0GxbM4hOSGrmf2BuIDhn6APDa28thDSQWdgf6OtfrVDx1/yZp9ElvxiRETLKfmgIzX
SR/72tx21GLKUAi8QytY1pe4cSMyVc/XFoZi8yI/3C/g0CeUdLT/4UluPE5sc9yoLebOeLW8m690
wcYQn8B+kcGf6s/ah+XxyT7nmdHSbIzVoXHpr3lk4OU0c536R8Vzx6clPkaAk1PnNcI5H5tdCBqY
lgzdzNhlJYoS9t+jtHPtn1pVttFmDyQ80fzyIUesbYOOO31ayE2Xs4+s4hgzqlmaMAE3Un71q8QB
CDEqtI0HuEaokf1Isyre14i/Zsdnu5kECps8YYOR6VFtpBo12rca7J4NC7jBCL5+im2a35oUg4hd
iyVm5oD1bZQqLjLnXtUEAqOB+WcPSa3wphXmHzzirG0g3D6peZ1IuxqFb0+E3nr8T3pwD5fMF7Cs
a2x8R9bCwB7un0CiQsV4WP47l6ju1kA2U6eFg6ZsgFkFrUM+f2Kzmy/2momUGOchLqmeXE9ZSZ8p
yV45fgOfCQvBQ7x/7CGedpY0S4BK+opLx5QMaf/NIVP5LGCriokJLC7eRSSe8mlKhxxP9yY9yCoY
R0fWgAm5G7Dl+HSviBFOmeJfN3q9NviCE3InaUJJACk6E4HlzgWhVqcK9XAg64HPmLW+uZV7ZRt8
uM9bKdsQUIlADmGrZ1VkUTXGEqiq93zhONVpqLec7Uzx+8BgV52DOFc2iaLo6FSJ2fKD4uctCsiV
/qUcxuikvuyV3GV+lDRVl/PbnZ+Xd7YZDhmOURQR+XuQXREZnN9pjdS0g3Zutt+FEzvqHbv6+IAy
xV6NFdMlU2IUtpHfh7e9edLWWOJbMT7raT0gdhEiyOA9X+z47vSh39tT/ByZPCAZ9iQvaY2HfwSA
FyswoZtKzCGwRjpIV+30jiIw5scl9a2O+k9TCJnHWnoNL1F4ekFbNseC3NBZMXH9QWUy3WNR0Id3
OVJCQYOlhQlGzVFBgZiA2AYbtFYz1ihBbMX6rXZ2oiFJEMoyfnFCVD/FD4T5HCSKdHeGjLoP042M
LZeRDEwsxGMNC+k496IkZioZsW9boaZc9BhcRa6pNvskH3CR9OtaTBvrilM0sWgr1HB85IQj7CwI
Jlj3x9UxHqwObz82pE1/zrItKBxMoEIPbAmx24cLqlEN9GEY6CUoOjv87089HHW//IK3cwhR3cCx
UBFE055u2FsNfuLuI0yAlD8EMCyX8UJ7YnIEGaZSWAU2enILkM3NdKLKyPjV2fE1to/5pF9jkndr
/klhALm82xdxN4WQK/GxmPzrLz6DB0JI+JCMP4phLuiQj+/EvXUvNS7HwlihxMf+uPDS6/8M4A/2
IAEMfngEZkXIYctqG7jO0ywIG1hf3toCh2n8bMq/Rzvy7Lnilwy2n3Z2sRJdc+7wTLVndG/tWSAm
Vx9YspsSYNs6L2ZHEzYMtPV5f0OhpUjAX3luE1Z5alsObjgRzWtcoJpVCU9DuFym3+bbCifoH5bT
a4QccSosf1md/7dIclqjsKGRn3gRjsR1i2pXp+f1akIX8U/xYbfjAW7a59f9tXdjnyag/dS8Khkj
agVL3vsr2O+DQ6WWoqsSFniOuslfYOkeoGY4F7XD46w/icB72PuNCy//BH6DxDVDJBxwzbh3Rbaa
TJS4wY68OOIAqUpl20dNoX/O875TAcZXTo6us9dguLW/AXfdfnOSRFGr3fVE0YcLTEExsOakQUAD
jct3WFij1uFHbKglsYGqoQXHRV0BnXRMylcPjGr2ApQRyTdaWl/c8claOvMJIiMVyiFtTrUqALBH
ipV5rjYYkqfQab9yhAJHk2DtathZ8jcZ7sA8hMbkj5dBSUATpVhT76ImfBpjSzQklSEC5SRMPM6E
2mLAHI5chVg59r0wblXmiB7Ci/0AvRjoIW7PbYah3010VZmI5VtCm1R6m3oP3Zd7YVkeQ8HZYFAs
SCsUOd8UABCWR8iMg4zEBzF7U2CyiZam/Ofnnwhmc/d+wWm8oBIu/kU4QxaB4n6QodiFpyBlrV93
Xg+ds0EIN6IuHvn3a1zarBj497MESwivCr3JOaOrwAShEUL8rjsBjB3fxIaIeB7356W7S2hW++zY
+khtTiy5gBb2idP0satRmmkWOAKF5uKd49i1aFqbcgOswbkgWzahjnZVvt1aaMKsuENAzleUykxP
8YZfHJOf/5y1z1IGjrPOenGkLZmhFEL9goQvmlQFmXR5wY9X9YUPnJvUXk6+1FP9u5caef/8tZyX
avxMvbtRChoYc+MxNNJhYgZQttMCr1tPK6k2pf80pLaSZ/oOnjcr3aXhzp+CMI8T7dQf4/UXlSCj
UTjMiy1qhzTFzzl8cTdKslUmpQrqMlhiZWRzssfiqC0Vs1BsMw633bWYOSB9Pt3FxYTjsJ8WGTCC
wbG3OWVZFl0DLI9JgENs1j2/p7GbH5Cwp6vM72cFhUy5ckIlh4oc1p4SD4U4iDmFVHfOC9RDueUC
6Ba5BBscQxlTIT71DvESB/D3JD0+7KuXMfMxf2/TQaiczJeKZ53G7RqAoYa9u+OdhUPoP7mxeY06
ckXSOnzMcww9XOz/9cW+IEG3acKrY0nGBXrJ/e1zKV9zTMrjKGdDDMiVFLDprOkzOeUe/bykrn6n
CTKc4QdiTKeuH8UigTHkE8ZfFQjezaWTx/UWsi8jnXLQ2elHVMpYoU7/bq+fMHCZ2dEgt9FE6C+M
Recg1xN+GkqEaA22y/ruhcCJBkQ74xmqyCZfUX64h+EjwDmOfrSx130jtf8nKpdzNsN9/jt3xyFX
Zs4DKotGaD8uUHpqEi9Z4NlUvAkrLeUJFqjFtOiCCBnnu9sedPFT4+a0cZd/oZd7rqtduZ4xWz88
G3eUisSRotDZxUapPUUMA6GiClQ1ncnJkeopORMVO3GSxUbq9UJ8/pQfdm9Q+6Yk+3ii/+wot+5J
zGDanwh+RyWrsUUgVHD0uIX4hd17AY/fPMu/5Ck40vMfJNfv08NPIY5eFM+WqFLblij7mUM5ceM6
qHYuMYqaOxPnsAqY+dV+aCJ8SRucDzyiOYh2ZxGrtq2jlDaKeYp3SHPRzQBjZIE9zwjPcN9pEK9e
RqrxE2/4QJH0GvmbkRzsWawobwXVFII0k1VSXTxRYe6sUaUo3ykEDwvc22nfCMhrWvxD0vTpdIME
2HNSrvl9sQq1YqSmsVhoEBOAdBlld683bmMiwcMnIMJoZSlhWUtjgFuf22mvpPVMz34os2k2JQ4F
Qgv5ZhVEKbY60TYte6PtEBSuFezWIIPUlGj5b9CJ8k0Wzo90ZDCgCH3zR4pAaiiUVhdt+ovRjvK+
07vecYt/3YV7KMEwNiyVkRrpJID1+aUwl2HNtezS7AO6Rj/GyMWBX9b3gFroQ8AD+b4YuMYdflaj
WnRgGlONl8wysmXLIgm9MAq2frWsQlqzzTUMkYsakn8r6649OQP0ziudRn64igKKUdkCX2q+75dr
j0lAyUKv+QRJLkiayy8xyxY20Og9kJQtCYG68c9kXmqynWH+qmBmhMUKmsA8Z7jstcQX6hQM8zpZ
gdnl4mfKzveKZeik36xl9/ppubqJ7vctvqoZhWjRpNcGGFWowxyuoOBBEy7kioqUnzRlTYRaM77A
Dn9ih+DGbK2q1rwFsEpCi+Sq31A/KimSL/TWHD1YHv+iFbDOa7snLhb+9Q5VwN7C45UAV//0K+ds
4V1tywSYjcOB8CNW3qUVTjJSDWnfhGYCpKK6A8wDyk/IyncgM9DSs63uKWzhANy5Ydj54fzszF71
jOp4niKXRLI5g6SaHPFnmZUzqkmLcE0ZSPm/hExmLsMf3x6a6SQ6dGTc1eOr5KF6X8PH+TwAqFW8
KlJ+YCX1VdArNGOt2XX3/t5lvu1No2+uXzKT+DXzfpqWOUC2wovrbacrcZdqcCzAjAkOWhKpgJvc
4BruQiZhJU3WsZDmvRXq3crcTgDev5gkZgeKuvMNtFRxmrIpZXiJIS7O2hAz8B18toDBgWU66hsF
PwuOZ82/Qq9HxcSmzmH6536nv1SHIjzWotTlsghXpgRPldDy3zp6hcKPdcNYSlbFEpRJmMNE0Cv4
MqOCZKksA+K62+npqsYfgBew9xoOQmCQDqnSnXZSjNn3uSZvOWtMo+Ab7yTfzrkIK7lEYtwuQS+q
nZ8gmgPTgU14aLJ0GevDgQP+fNf5X9Ey2yaTivnOvdK3JDWCVG/+OnXO2y6kcb1v/HOCzIKnTPBy
GfEjVMS5056ZRoziXmLWQCDb0OH3X8EflBpsCsiz9HfXrp1YA54b5TApWVkQPK/oCe9coZOk4KXk
P9e5xOvwZuIlww3bWgcHohpB7V3riDpBc/HsoEIlCcyEQjzlpCYl0knfVCW6YBLSJPmL0OwLW4d6
ktyXtF/dumQeCt2uKSJFE8vbNg7n/npZRCsgVnkpZREfm3q2cwM8FNFhr+nLy2K++Qt0fvYpcrEX
x8Xbm5owmg7wx+g4jinCMRLEGl+/2GfxnRohYoUpMSmaLUWccsEcMpg8066w1AKUrkvOSDQKHCZX
JPn8AHzrinRcuLdRtvqldraG2uRU8XrfCk5Au7bmujQckiLWmVgFG46iZ4YjpWJFBag2ixpqlThz
CMbCPIO14vWmAZzc38FFs0i3qWtOZk5EX3d7tARA6CwBVs26U+JxKOcPdjPefvqShdhyalpGP3cI
naepLo++RT/94R/ZtPrtHJIFnIt9W1V8i2xu1FFvTRD/Hdoib/hYiLbrD7av0jWUWr6QDWXqnvTc
Wtu+bMMU5R9uvyl4zo7p8STTh1JO2iCM5rHEZs7XRUhOmMruTOvcxwGrKjrm7ALoou6HQKSTds8J
+aUnxOfUkNW05/M/pd0bo6MNTQU8YXGfauSB1eT9yKXfHIFiw8Si2HlfCHUjhOV4stINUumV+9Vk
w7RjoGy8dKHj1pPUraWe0hpWRCXNsZvwWwyXhiNOZF7+NzYzDdgntiIrVeVUOaD4vRtQETXKk7TU
Q1qnfU38/VI/oZJJzPKlRpbBc8PAm+GcGBsQ4zObJfUc88Rd1fpL5opd7vGkJP5+qdvBjZYNUkDx
r9HENPV/YzFqykZNs5CGpi1vaxxA4iZwOKA4Bzahw0uLomqYbZ/Dsw9PSI1TdxzCAJ5ywCFESIX9
q1CfcLQcHgdBRq8KcaTksN9QWBzzL5L4QLuRfkpftcWMC3se8b+2V7KD1SXxmTIj1f9NNeOneinY
4DSa0De4nopiEfXkh8tXxAgjUS78OEK9jb6GXB5gTS4HTchjSf9VryljSUN5EKorLxZskDQ+sGIr
xXeuigm4mtLi56Fdsy6rHL9wfob2yCIsuDhKOcinAf7eFocC3J2vhrdwwpVguhVYv+/16kJx9dMp
ZOif6gMbiMZFfyNT1C4k3VULLxmj2ILdhvOcJdbpxcy4I6F0IAASyxcHVKeYfyAI++89lbSt/wKf
XFWWUWeRGVgrjUf8QJMf23a0XNhVvA362Eag49nBeE2CNLviqAirTDyAniF+wmfphaskoDN0JPyf
rtkPItFRGB5pJjtWsccULeSeqi2WomsGrU3vbG6yLS211toxbk6yokqZIq9uqiLj8uJ7HYB8tJ4t
oR+CYaQa9qgmuHS4/GlOhzX9FmHMRJDBpIT7yVhkAZX7KQZriFuZbQJU05Qj6AMHWGWWWRl/mG4f
dVbEe49lo3F68/DEaVTvtK/B7swuVxXKqv8PJtjPUJ72uXv/Z5BG1aXzqvZ2m2e6S7onoqp1XRQC
u6JzHdXiEgX0hbR02f0qEOm3xlniZRexw87RmlqXBwDdSWE03knlex7RDjSnSzY9zK+FSFwQQXtV
P/qazZTmDtjpN/WHGJdsnbNaVhUCwGhqfv7H8G93gfZgwp+WER3VvXYGeIZ2K58n8cCR07m7Ck+F
Ojd5n1i2WPANaVf8IKrda9nnkgemWAyc9WdkyG1wx5a6kiKBgJPJWUWQ3Lxi6ZsjtY3DIq2CStNy
HtqKBGO/Z/V+zZ2mbDl+BHeOw4ViOZYVzdXSRPCp3o6oJl2c7rxLVFjVa8CTFl27U+GhJFcPfMyE
X0WTL3JMDV1XDpbKaI9Hefca6QDQX2kHE7YSziHGV10uUt37K9RtaJj8+05ISexKEla6f2zPjNng
sHOWGp/gQMCPka3Ef8o/wScqOLbwjBCcVB5imQkeG8S1OIP2EmK1SduJwkYuTibpB+jZpQifQ4ZT
BK9YsQPhHJFiIk/quZqkPgzcKzhjENHGTeEAdVuUbNBX7FNDVWfetXA/dVPtumVmXTTWjmnq7CWS
puy1ZuFXCyX/CmKw0omsEgmbO89dJKOEHE3mFOwvqpbNaMo81Lfpc1AYJJtzGtd6sQKIZWyG6CqD
R9nM4fiUVWRmnq7KQPCxWzBQJOQvdS8woGXqdSpImXA53EpibiGPA69XSKsF0NBZDbvdpRmHDlFv
qvxzHQOqjqn3y3HWCQT4CqyndtYvo/n/8tzYaFzd8dSVMH+j+byzxItNEDVDvPDmkKX0gg/YVeuE
1aM6fYPzrko6fnIis8kjSbOCY13N0nGjxhSbHIpl9HrV9+5ViIo8QR+VyfNoMgbNAH4kUmtRIk19
YC2Xo7RwXgisxlio6CU3LlUS//oX1aZkqY7odgralMknrN2zadcstkAAgxtAUJIzL46bnf2Zusyq
Q4CAnKasWq1rbJbCDHyskFHaBDfQqLxKOO/cb2tYhRfdpTb/FEEFu+88sRVBIMtoFvaDgQBZL82p
Xd1h+2CmlA4D7t6Rw7tZN19A94FHnOVfsfsqtD7UmbKlx6yxYPhWR46BgT/zgRz746TcBh7uki/d
E/qPTMy+0ZV/Jh1OfKZtJZoTWa+F3YBK9NewNk2yZ2/UPvBCeDj0jNy2J3NTeEn6PXtPInuKic7r
x9Fs840Uf6TpwgaP701TZaFSqx3ZZ8fEWo610IxPeJzhkBGz7S2sCQUXtWNT3w5199aBSBYL7bXZ
2JxuNzlKzn1paJu/ACnNXPdq0BvtUwp5zBYHT7my799lANGYIlSCkB2UzUlT1fPkDV47nqQsXcRT
7RY5WUELNpNbbVeL5tua3SFCTcMnWPsTafo+Tvl9AHn7y6ttIdbIK1iG0E8F22PxZsxGUqvxO7ea
S2PEJZUCNw8SMmjDx2x2IV3AnNmdwU+k7Dpy1T+VLPfC+DGZNVr89osNDsmbLOHAzCaNYMI1mhb5
VKte/IW4Ik5utVgFc0syvTt1mSPwFkp4CJvaoi6iSrzXz4DmQQ5o1zPIBvCxVOpTutUQudNTZ7cX
lsN5CIW+1xW89jo9EtMXE9PgpTCJiPcXK+3IQz6RFUxO42ZrYTsVpVmcwXCStP/QbDCQbMOtEG2z
/rdGEAy07/MwUAKOA7B4YpxXlsULt6CcNSxIxRDhSrA9qN4TCk7ClmmmTYUXc6swPnah8YJvy+aI
PrM/CIxW3JcaF6NzrghvPGqdytMRt3OAX6bxR0XbUXME7mtixnxucThtN4rStNEn70E15lJmEB53
5IEOEj2XoVoZBAJQQLoHMjlN9zEHldRD4zDiwXimbeZkwmPwpWkCgIsNP5vw0M4Ko9AS8r63kqA2
WRqXV5dsGeItdWKuGlFyyFNcQq54zUOLvon0lxxAva0DXAudvxlgFwN/Zm+c6Up0WAV45UVsv3RH
JcmgSQNpVyrHv/68oAS2EvsOcQ3vjW5iGBWVoXgmYSavYcL2fHVipzH43emYfR7bpawawxYWVWJJ
NR5osd0b7hzJQcL6qgBdp4y+z36PgtJLJYOnKRRknq4m1LPnM9FVhxSx0wr8DhveX2Su26qNGhf3
7DROubXo4qzQ3im/Yjf9/bYvjeHWiQ5yrDQ0lt4ISncAM6FtcynyUu172djoqAQRhp0QLKd7ozZt
vg0tONxCQXqmkmPLz6RJQ2/qnsnjCni0we51qN+ugVMvvu3hZDo/XJJJzl42PcNFwVwpaRxHT0vh
67uoOFMaUI+XIRh+8TRhB7+XNOAfp9U4EVbH8frdZFV0p1q4bBB6tqG/cMVrJ4YXPgUJ7nsMFvxf
5KkPeviSfkmPB8dPkVsxII++EErGxnY/J7R8kpBQWpVYoM2EeenT2HNoUxL9NCi8b5d1r2G7Kc75
7A3jiBEzuC4Cssz1tfTT/bTsQ94dedw8j96aA61JaxgN62sBELw3KQnKmCauu/PapYshanyGtNIE
e5n9NGHELuf0w5Y8AUDANiDvKFQwldTIbnxEpko/poDKB1Ye/OujZK7PU3cLR/0zTc0eVSf0LzXi
f0AYhKfCjQ9pqX2pSwx06d8n6sQO2mMMOdw2TqYpIZvSo9Xf2r5nsI8c7+Ax84cVUrimV3oNYHdO
C/B7UyUusdaFc0ERkZpM94C9gqvtuAx43wqGDucMaX8Ya+oOdWyJ/Geu6ZhtNfmHJUYxvjWkdv6d
jZnYvUsxAO8E2p6MThrVe1S7jr2r5esLabDHy//doowVCsTxfTlO/nHFB8pbNUskuBWQftLVJI4n
yC2NMMV9HY9f4yHMsRjcrSA0BJfCP6dNzZpXeE0gbXIRCExbvehivGCDdu3X0nXkA6rGY+nP+EuV
K14oPoUUECDaEa7mcNjpHO4DJChmcCwgFO7jRCkmfnBH/pBZPlbtZT03XHHoG56rzvAPQPK8Dhq4
pxl554gA99dxnaHbDO0SarNHjP2kBICVhUlP7ahRgJP8xpO+cnhSNsxXGsxPopgj6Hct4rXouAvB
rcNbEaXWF3rFRJjALIvxemcIKV9T6uYt7Q2mseofY2qhI5BcjO7E1LLMOH4Wt+2HlQ5ba0XXzrr9
jK3laBaK1H1mtaTvvuXBi2otv7VbCm20KI6u3BDEn3qYTTU/8X5ju3O1jZdnPigwmsy9rsbv0wPS
TXPsIrSyRsWjOtRkZjn64quL6/AfgcQjfmjSMdWd9LPyJk/l7HX0PJB2dj6bbegKG4mwUYF1DBSC
CEU/5ta1/mR8Io6Yk4+SKeR86TQfFZFKnoj43mFB+7CMT321ExYHa/vjyRPzF+TEdCSl2f0MkQsI
WND/cNc5tAHZBCDPABbS3/+1GsP2edzcIstjt36SujgYXnmKS0FTuLTu4zJ5if/1qjvEDtCt7/Ni
tb6bh4lNuRvZLIc2Ph5uuZ9zyl24YTVFf3BfowAQBNW2xmvLZ2zzhfpCMeZGG9lIO0LJAk3ey7II
KBXU+ioJ2nR0OVXAO6p/yFe6L+Qn40Mf7DOg/Q0Xq3txpb6qLgz9fZvjzUTdG5bxqGrfAO8wEdKi
JT9c9k0u/OroEZjSa1gA8Frew+Ujajoi+EkZE+Gg04pj2emSq728gKtXIgwsCiGSRmVuNK3ZXv6U
1MOUm0NIFAbE7nj4zG1JUR/Wy2VNFXBRpIeyLcWEZ9a2Xk9m82ihMsnNYAR10ZWwIjc+Q8dei2wZ
oeRJW/f3p8PQ49CGtEUPTF+varoGEdyYZ0JeQ4RG5tV/Sq081oX5ir4ryRcf0MqF9453H8JjeN9P
E5/+k0lmcz1XrW4TeOsFZ9kLpAP4moBy2sOjwFKI1RTl2CPLusf3LJrr4vz6thmd9sVTQ1GAZ2yU
mGkdHAmyhn7u62HBTLNtVFR7IY788aL5GbtXkx5CSZ/RXoy887vwoDoJuRdehX5fptHPHWMXH1+Z
JAxcazHmT8JxgxvI3jGfUfRj1ty+5fvPjCGCCDLoWuYGKGHbJrx5vkLfLnrWdLhAf2128yOl3X3W
yGCJ7YNZ5ATOvv6c6509vFmZ2XA8Vumu8FwO7kVIUoMi+xJEvVNKyu5qQJ+5W+BNiD8TU3Wi2yyc
WmB3aSVB+B0t4qHVeE5htWZWRoXTVopm9I6AXYRAcvBEaFNeuhX6yfXN4/1xto3voAZEXzXhfiIq
l1p3OIsPcQ95pT0FaYUd2C2AMXmLJltT+O7r4RJyLh4BGdgsMiBgA3nQvt8mFSpHexp70SBvLc06
TkPBPOyB/Uc8qxKRt/dYkf5nbJj3ANDaWMwHZDRsxG5f+b9pAOhSqKrGHKIJPHT2s3YWxsJDOGsW
gu1cm24EixD0HD/29NDX/+xMiwNmiBnPTl4AFssqmEla3PwewIDIi3iNMqTtbOENErgsqP/Bsm5m
UESeGeZoJt/cHVUlsLFdHVsdLZWQOOKPPS4hXlMVymCO8JRiRAW/ss4qQoWb5Ub0dCxuANfW4UqS
nkTwbcW3lNy1VYgctPT7J/sObuJfGhDd1wP5OUl8GkGztH8QU6wsctSAhXsEHQwiXRD7K7i1ZtoU
qxebJQ5wOf34/lidrfJ1UVrOFqslkRb+pxHKfMmDTcvBtp32MVzYKhaeD56k5/NuwKfTk19z9b2i
ibY1OvD8nNfL2wItwBFDujiHGm4YkQdmnToco8g83DYXHDK8tDJcJIi4sg0Mv5DDKbewNLcMOZJa
8AXLi2DnL1PzPeo2KuBjes7Cc6UjD4nC3NkdDBeqOIIB9Esw+rWsVc3gAjh+V/F0hsWeUm65S2YG
DvpLr99bRtT+0Kb4eV1VgsT5aMdpcTSuT2QtQydSZD2DAYSnzeLF7OqmoFqDm7rIB7gj7YQda+LG
nWeDkVhfix7j5+boSPk5yPXSd4H0QrDERrOif2I3rLqltik4vT9/RYOKDvtZYEVyP2rOQiqD1qFm
DId9e9uZqPjTFbZmziYQ0uNix9UgkdkbBj/AA8TmjEtpb3f6F0G0qSMINrTGfd36by+o440A7hCi
cOMndFoZc26Zz2c8zjLjdKtQ3nPdhwEUxewRD5bG+GcOIjFH/Dwxm5Q5LHaHcA/BCT5/79iLBIO5
ANohYsf0h1lFvVgtIHxuOYWHwxay8Ux1YsRYnVTQa+w5yQYb+A2XCCzaIirfOIaggQvJXodhabni
1tGBFf7FKMwyXzZJES9QsNyOmduskOZK5W8golhaiFaxjkpsaFg9uxyVRDn25tyu8CcPEV58Cj7K
bh2wdn9viRPNCY1MgeVmxH0pux3o5Xu0s/BzSNY69jeVHbYA6YnPOZuuY4Er5fKnM4Fg+zZzi51H
OBlNZJKYBePkMCMVbS38K6Vk/d0wydmhE6XQ34yB79t73pQaVuJl7e1Kiij4eis8A9hYfazbKL24
OfN/42RRiIPN5f9xCYdszR3qcH3Iy5+U5N1C3xZKP4w5BVLTK1t8FhNz3bgE8WCtuiI3lPZtba+q
eVJAsNqfSQFeLbs6msN7HpT9w0zDhEDMGpmPZ0sq3QeSS0jVmjdZcIvF8osQokxZmpcrx0yNTpjr
UDCJyb+3j5s0eRzV/EDwJsFAP8rjwBNjvSb31eG9GkGzJtk1d2x+xPtbNf0QACF145ZyPAkX/7nU
5SHiTfEVQQfIH6uTrnDEJUNGML7Ca1WF7FqcacSrxjIC8FAF8xZVfKonIPzrlFH+Jd7LNISei29x
sdsdO+fjzhKC0H+5zxgrmfsgGlHpJMPlufV3riHYxDu0NkejF3yrpJ0Q28phS4MV/R6oHnyRzoCJ
iR1t+XyoblZW68c7bYSyKdAXYrZeah3GyFsluYRDm8Hkuh8RP6/9UM6E7LlLNmqg7Dtp8pdPYlj9
etLTViTREnOjIFOYMsgGVO42nidQpmJMVZx0qMgv5gJKKApk5cz2HzLlZBEVwGdzB+2v6bNbGDo3
gBzj9vUXszvwFTb6O+n0zgohX4JrCIvqw8rlB5ZF1rVlIODBiNh1qg1AjlGj4tcq2W+Qol+a8mvN
0de0B41m/VKniCMuVKzvYcDk7ONSkdqdFtUuPbPOT7zZuVvWVQTEGB0eWgY/mXEPetcUZ68QOSid
1ruPShtSDm+1M0hugnCBTNCqRjPFaDwaaLZ1OcXdbK6p070yylnbHJsTU0EodWnka3ApRbVDPRN2
Fc4siwYQ/SU1f/Teztvd2IOWyEBV8lc25cqPqhpsl+3ECXkcvZ/o8Tvpz0Obt/mQCe2g1cXdjaJw
B0s/tUt41yV1n1gmqXBpKQfQNPqiOu+Y7dyQT55iZ9cCCyzBu8Xja41ggNXijeja6pBqBLu5EvyU
O/I5uBOxrhmQciEupdzy/KMcKc4rcIMBBW+nU3VMV9gn/dxBJP5on+8/JI2kO9D9fUeAubuxLo5u
MTgNSfLXl5Jd7xmnzbjUSTyi7B5KPNviAlqebSlkccu0S1PUD6aah1y/lgbeQKUuqwJbWhLbzSwz
VJEAWdjfJ7ZIrSyXTTg+k1fTvkVMKnRDNLAZfnRghCryvK4QnkLz+b+UtUHkURtYb66++gwCN+rP
ddr8H7Nd5yErlSj8LzZVvX9oL9b6ullmsC0/FwcqOM7ld9QlTXalGYO50vbAsmjs9o7hYul6JEHt
VZ9zgusmztt9F4yj17oNLpXkkr/8GXnPzU7oK20LIilng25g+Q3aTY9jY4bu+R6gXXVNCAUUQGFN
rcGr+c4jlgxjg7RSHr+FevvMUAumQkmeY8gsqr+ycwN+a5m/9E5Vd8h6hBPV3aBSDRVvUn/us14h
W1TyeV+tkIm9bYdpZMnMmmx/6YlJ+org7NNy5MHwpMbAPEXGUf8Iz7qr90mVvdAeOXKj6E1u7KEI
b7jqR0bHmB9MBH1FSnvkz5P9vr2L64UpaJu+tFvsZlEeOL8je4DrRFamTtU++VXg5Tu2yTTlSePL
Q2pvAUag7noWNeRZnjBp9j9egtVZMLil/2YUyrbfZOdBD5AxwcUgl7g2oai7op08J/6ZSEIZd8rr
J0g/+8R0WXyW+gd6DjxMea6/8r1TTrhhOHzeN/r0xzWk++mbe5lETPpWT1Hv+nSVDaRzAkR9WrVJ
dMRaoYMyYgr4tmUDOsER7TIRKff1Sm5amFpjMp9MVjqa/68EDb5Y2eTlk9xKsmz7ZVZu/bF1aNRg
ktwusgbvUNDQNkoixFnRInr8SFdeYO8gu2OaR4ag2hJ6B9Tp1CV1F6GZ664IfqHPtEQdn1carEEr
jeq/Td30S7xquBp05E7oJ8WT3lq8l7mda5vGJgLleuoUFAMqSS7cj0nN/YvDXSLtrNXG7z65nCa+
7y3JU4ONgcoc6FPlVHDBdRewWK1zAqlubxsmdeFQwBWqm1RG8ds0tcaOFEX0bdmVlyjEKAJdLI91
vj1TQhPJEdR/oLR9BhcvVAOmeQUUdqexqx/UsJx+H0RIbtsNmDJF7+Rlb6nySh6/CxOGMkE62H4h
oe80E3NvZGndfdDtUfVXIVv1/JR4Kwc7YIb7AgMcUgOMmPa2pLlUU+l4t3wU6tcPvDGDluSNixX0
ckZah856JMb+/Emqbt9jxh8Z7/pqc2OoakV8DgWozjrrl1DX2+i33DpPshSPfKYnzZi4OpSrtNXR
PEy5diLzs77Lpp6lgLXCkro1RJYGDUFD6nDDsu0gFNBiDHqEUhWkoGWh14rbF3B7NqFCK6gct1Ep
TTS3v/3x465ST6vJE0H8GLak7uZwX5H4XE6JAgx75/LeRvdHPWG81qppZpysftj/7jXnrsEoueZ5
eUKhDuF6wUmYblrDIg3J8+QRNP6M6d5vMyI2CS9YuPNXXAFwIicV4fXYhlwnkdXWM4LIhK9MJgev
Pk7CGjJB5fW6jnTdI8uXRV+oXhvMVm99TA5CEuD5jihY5wprboiruLRn62fwrLwnVQtCvRcf8iqf
riKbqPHsiN/Sj2VbCLicy+zJfFGV48T+5dn791aeYKGJWMg7GlJgRDG+Yj7eO+qpgemZ0bVQUwl7
VuSBTH84vveSjPF3f7t8IubZbOQMBxAZbEesKjK4rvAZw3x7MGghk6AGGMZQ7f2gsXdR9Z4XCo3I
4dpDC1r1ob7dXokZa7kKB5kHFXnufFEJvEdiVO85Zw4RUT9wJAQWf1aR4ELJmsFSHquXhsNgzY2M
wOb/T8YKZN+8p3UNYhe6Dt/fwN/2MnXPEqQxtGRdOAu8MrEfLwmAt7yrAU/o4qK+L0DX7+hjwEsJ
OGtdv/6xXG+lEV2M6CudzzC6IFq8UIlY5000hbMohgt+PMxbrvWQULEhtBmgxHN6GWWliqY8bXdN
04Z7MB4j2/80mMNL04EOYWsymkl8fZk4kaf18jBGw2X5EEsDoeGZwHm16w1ZBUYRpS5ngJulbjjN
ByMSgEG6N2TGF0OJKyAmCFDbZzcHkeKrtGxYX3SwUlapxXlA8NOt4P+E74936DU8quiMCVxPaDBp
BGSoezhIvKj2Lcq7UXdvaYYvbEfMicgLOkeP+Fnn3uu5D2aZO7TpB+qGdvyVRLr/xJjr6LkMlfEi
viia0u6zM1aGtO3gbRq01p9hxGP6e1Zb989rEOYN760EEmldhj0U9Qx0XQrL+SU7+MtkqnUtzY2v
7uEODlioiYWJBRjMX1hwsWA38zm8gGfDB8Fvr3B8Uc51NIRdC9uDbkbiGlx20h+NaHA+Qzi141zr
5srwUHZG7j+G7NyYP8rEkxgDTJiASujaAY+tyFvtaBNICXmNe5UeUni5wgS2uC14v/eI545eQTbl
NMW67YOiL/x+MWK6sUujn3fEMxlAEVCoT7/gQYgDvU4rYpcRT7drcxHpT1excgDdZC+5CmHtbdZ8
DIj0xs9REJBisFOlm86WUdUbGLJhp2GQvViRGJexkItqkwPgfwtl363F5di0bk1s/YPiHRn8tQDe
wIh7x5e/b/HV4uUizo1Dv7yCbIj8cBspvJcud36B1L7mph/Vg59B7sjo4SXydYx/ZxxAx0EtpBCW
jIBEUZp6lnXtrZK0EseGBGX5171erl8w1a6lFmwF4aXBmocV6MC2t8e4TeIzUUc/J29qqPf2AyUW
2ni+dnjInkedIr/1QhT5trg/YkDj5bbIHnYdk5/3HPZTLRqSA/D33bNep+9AVWg7bt0OAd68zu7d
KB31gnV6/hOcsd+U3SI04Sk4/8VNSuUDQTraJUkeBjdW35QZnXkBfhsr/OMIs7POF7XwjLn3mZoR
59x1hX6EnfoM49Ghse7c7QIlb065tcVYe7Uuqnysvuf13cllMaM7oNTropwwdV1PG5Az9gzYLQ0z
iaf/0q5//V1c/m+mGOWNOg7b99oDIpPoPhB6oVBLrHT9bsmMGFrB+zWH7PNArjBIvFWGxC/PzQ8m
G1XDxKD4sDUuHsbtvz5cX0mFgA0fCc++5IiLqjTo+zhNpc9YPcVxrjnFpfXbnedmexyEblrg3Ydh
w+wK1wYbwUWZtWFMTGI2bHcXcvvnsFx3A2t/8pQfBQZBsC3jaZtEW8thDs8JiCClYbQnetkmR/tb
MimweD00TNevp7iaviyJ3r0duU/EUX23WS0BrMXHFH6SwjjGF42FDIuU+LMYLWynBaCf9EfMjCoh
qC7p1G8cRJmd75uJTYZqGVlyqg1/+iMnGFBhJcZFGEGg2w6DBezHRJxMSE7aj7smjo86H0cspjik
0yIiVoIK8RRj95/kwEZF23tt7/SIvBhYS1cbVhaFNt/0GTfHUVh69e26Sy8CBCcvWx7Xj89vcZ/D
Yc08DNNZfCdzVg0HzrvBYhdofkTpz9+pobAl6kgzfxkU8GJpMKCnBsrvOmfpt21zyw9mAi/i6vYE
WukNOur7AMDH04FAp62HFc2e9s7LOA/48ot/zJcELCVireHxXUz5sdtEb8H7QKDHphJVhKhjUDe+
sUv6Pa4f6RxhONwbXEULqjgtf8ujWGjlqXkoXeIW/kuAXbrfo2PoZenO+eleGpzL/xQJPDMRxqHV
YhNyZFdfcdFD2wZb7r0OoTBDJxZoPXrSpfHQVvwaP76ATBKL+o8QxjZljENn2UGL0OjU4SawTADJ
rLGzmq9cyVuf5mA9CWUr/znlxzU8vK+/LHtju6mIPTwMPFGFkjy3T7xr1OyO7yccECpG9kRRHeBU
fyiaS+EGWFlGAwGs5Y21RznTrrWWHJQvuxQQhRlL8wdxNfIimMbLAN8r8PXc96D3V1u8lrzGYLSH
uZAt75eR7qZwjjI8WpzZ2gEwDzydx/ZiUh36hiGPzqQlD76ZbbMd4VrokmlzkiV9nsOOsXrn+CP3
O7cRNZuzCLbhlrmjv2I+0o4cyYGrxf4ULxvLavjH1fcxhGL50WVVjQK1KGKUo2N2EM8QveepYGEj
FRN1AIiFPKPnN98DFO0f/euHJeP0DZuyPi7HqX3EYqzLTB2gygACM11feAvy5k7iemLJAtfYpulB
IPCZvDZZlCXUi/ANGuyKwyRZwXYlwllnqeVfe4Cq0InCOwD5VyQ8c7t+El275PBFDSrMRIwMLxgg
ya/mOHs1PqWg2TOex0wfpNMKDJvbzh21Y6SW6a2reNh7d5FPIZOW4q7q/ZnKNbgQRyIejjwwlw71
v14WpeNgTvm8dCX7wVQAQTBQgNqdJtN79Lz3XgCcH+XBxXYsHYydg9pOyeVazeWm7v3ag88+hPIw
so4yCvJsAxaWxMR34XEYUdpE7aTku49akWBUohQI1fsTuTzfGp+YZt+ub9tQZWfrTjWdXjVpjGad
nNkO469KUSu4CbS+GB65HW/XNuXPo1iULFESw6/HjNuKUO5dfr4WLKpt3pGxT1TY6JJJpnw/WbMc
xKFRduliodTP4VejAXLgHf+O2E6Ky5BkgoH6i14VmyGdFq7a7rmHdz/Lv4uZvwdzXCTsLHedGIR0
ovBv18713xeoYKZZzVK8A9LIsb1Wb0n9lA7PZliLq3+1SlTa9fBi8fTA8zrSlBfFSJoCcUXZCcXN
SccEkjOa5+DfjX7jJlddNaxL+DjoSYwRZoLVwdBAz+LFq0SaUSKjD+BS8GrIoaPPagHmFXkRBmZn
lq4PF2NtrHJBluVEJRiBT71qDxui4jYiZSDleROkMNU1/oGtiHcp5m5OAEgy+Gx4AntO+/nz3P9H
VUcx8qdXJY8KrsA7tJbXJazuYgBtjkxvyH/0I7qCzNMYzQIsk1ar22/kN61Oo+ElzwToAmMMteKc
T7JXsinVgqwWadE5pjK3zCHTRCYaxIkgrvLgCw7vnfpqtPvZ0UFc2lB9wA/c75hLLOmKE0uUSbr2
C+5leUkOlFkOoKqDQBycYkfGcddGU2Boq2pW7ixPeDd930v3DtXD+upLQcCb9wNnzF8pCifsQfnc
Q1HStpehmh+TVHPVtilZXFlAzb03eqo8OvLVQAqBpJdhsRsW0hfZbDBs2YenghT9Mp0Co5LTg/az
iEtEipDyieOL183ywHpZfi9xKpsgXlxaHJvc4pCJxo7gHy7Xp5Ydh14lFinBBv1Q/WbbkDXJX2+E
pyd8SDgwU1RIHEpLWO3cnXA3ZsbdFxviEASjG5ojOaLzG3MlCYT74FjyN/OLJaZowx+OI7pbWQPF
qA40vk1KSfpEijbZLfdeBq5Yp2tzp3rkE1f95RAm9rX4kDpkzj9KmMCftgn56e9kf8RvBMFc55YY
64Q5X1lkWRzdMWvhvi6xE4S/oIkOFeq/5uH8ibPmKoypFnu5bcaP4MyVqV6vEWmcrpOQ5CYKXyR9
oLzihHpJHJFU2SxmfTqLC3LuaV3xsrixoI2NkgbhNQl1sRFcQ/tQcUnMEpMbPI5CHb6WSJqKCndJ
+WxOATBXp8H7A4ZVhzIavNURgZDdkjsccc0moWyvTq+j9MmuK0O7crAFmcSGa9Z2KXyUWAZok2Hi
ZmUntRdBYysv4zxDr5AHSmbkGAT+PRHHGrS6T+VJ5mgbkt5gEhUEU5ldc2te9F4q9v6wBvtNlFM4
XKrnIbf7iPG4I8r/xraLpe6v978vFrYM8Fy39Md2lFUy6JVTQ0bWFwIhPolLHHys5LIR2+DLmkc2
QxdolVpbDcBKApY9XXq1H8YerTMt0NhMMPdF4WLJVfOBPjziIm9mC+8pg5WBZaJLawtGiA87ofJU
TXaYC6XANOqkn9R74KUlZTtGq9NFzkMBAo4ViVW7Li+JOr89KqzerY5XMWOe/YqiH8AZKVU/z5BI
D+0dWtF5fFNR9+o7Wucnzp1HsEr32ZYgIfvLHHiqyG4NlRXeDu0CQ7nK9wH/rZuzRUxdE6R9ZXzV
zq+qA2d8+FWpfQLXFpJKPLPkYPGqMgnydt3VzrBbLOiNIC4a8ZXzx1TBLJ3NK1zdG4xfs8E7NjhZ
KyNvoLUkfLbR5NroefHE+60B53w8pUZlcolHuMzko33r031puRdl3hpcCkiQSssOt77m73Svxlky
tnGQFSYBTDqU5ll4f0S09ZAJ4zM5/IY+gmWOXpmn0cWtiGor1FAH4rxRXYxp+Ns6sRRw2SRTxDgm
PIqPTrU16dOjUTbeY4R+gQcUNDwpSo2qe900KoLcYYxaKzi1V6c4RQiqJe0eNL09PBHTeN3qYlT9
ClCi7nZ4EuFTwglZqf5d1fRCzTYGrDYRZ5D8dUW+w4idwGjdRTb3ejwa3ZQU7c7DKHWarY6matgD
fnhgrQsJ4K9kgwMmR2t6CxgChw17FyE3p82zkkFaSDmYy6OwBqoS+Sb9juUD6btwqmAU/Jgd6+M0
TNl0Js2TiTufF7ron3Ie+urfLzdC3Fp5y7OhIQZ71sU6YfEGa3KOMc7ZUXo6y7ZXZNakD1HTnGJk
0PD2c4QyB5/CRXs+U9dZssIrtgYNduD5xVVl7v7TBIhGhM80H0nwa0eGQ8oRk1uWLqulGZ72pC33
favklGELFpJOd02S8HyKEVDv88poXfb5o3cXM4QBirCVXsrgzaRRnKClFSEHHllroTJoF0n9TZiE
x+OWQ5cmMvjW47vF61Hn/n2NAF+BZIbVQElee47+rnTmu/xXsXKzcUCKwisLLS87LfHl1MeH4KLP
hggMOwsXM9v4luhbXnKW384zHbwjEUMzjauYk4U9ITRjJkGcKncTFR7nlSOI+WCSsfefYoPGAoqf
+26YfKjO4u42qV1ptkStTkMOxfn/b90HzsypEM8cBHvVpUbikeGHGm1Zr3cPydtBCC9I6FPtr+sG
Z2xPaDLmVSwZFD076SVwIzNDHwT/x7y7pXuMUlwUIwV09EpkzIUFrbwVND2P1HCFemfWuMbx0HAi
oUO7h0aR6vxZ1cEnmutXe5vN299GWwzVusNEMgP4wZzG1Kj+crbjkm8hGVL3XOTL5PQk7BBkmlhK
ydC2oBA/GDtXhiZTqOdO4ifvKMbRyBE+F6HvN8F/caZSO8tVQ/RmRmjk/HnFZj2v6tixIBdmsd5a
t5PrukmET7o8kVjVG5LwQv8jke8t8319ocWf/NcKTVhFevc7Q+kc8WxuQ3H3kHvbuWuiG3QdqX5B
Cw0UlsPkBh9cAxtuRNxBdAgr7TDYOjgkv5EOQA/xB9DogJwIFvYgb0XFptGoAkWf51XuCnI1MYA/
8nLx8E4GbtDEdtYlQhSNQrlmepmfFAdLP6vDzLE8ykRT1Ge5AEuH8XeVm4MqkineYJzoQ1rXe/Wg
wSgwgMEGE/+C7v70oH9di+l9DZXErE44IVmlMK3CfkT7+PhxyX2A9nAdDcWiH6rJZbDkXDbJ4wVZ
eK2GbAL304MPvXxfDng+bMOmoROANKH+0bih79YBjjb3opOQU7lq5DyWO/37k2UIlAhdvGrK9pxM
2avBGh6/49CjG7luYH+kOnlDi7lxHmA+8xIadDxPJTeZXh0rrGUKG+GFArmPk6lc8izKQ9+bAjCO
lgfRJ9YJbg5F8s9Ri3z/j5fkZoeLrS7q9Za4HEefU6tKF+iDsXbFA1uBSZ8T7jbLSgX9rogtP/JB
s6/8UXThTeeq+f21MOXIYnlqXM+JQbxdl7QOrZh/0UlipCuHvtVPy/X0rVJgVelWEUiVlXWKCqoe
d5Rhr6YB3h6KZK8oKsNtE4HF7h195TeJl2VceBRux0i3MLImuhmpFkq0frBmeXH3p82oKm0fRF93
DL9ZDp3XL8B8RmOlKU29x8o0sOrSANL6j6MdwGMGF/apy6m3rLXbUSKvdnqyTSPaoubPyyYUJMHc
fElaN26Fv0FwvS4e2yN6k1JG7eTBTIJWBh2VED/g0PK3+tC18gw45q/lBT3KAtibKCnV3g2VTX7o
f0pQuRmJxoob3jPK18dT+j4bfV0EZAcK0T/axHlrOUTVoaAlpwen7s1RFKOZqVtQt7ieOsD2JwTi
J5ssTewrTdGc45E2k0WbeYvVH+OmW4ebfX2re06yC3kQEagpiBkVMqPqsyXdRIKNPOSl8c8SPpPN
+q3Hod7xVU/1dcVqqdKY/GARmaJCPifg2cI0bdFttqpBbnDlROk69tN8yJ1b64mtQMCrUdEvNLKT
hkxEh5p6dolaG2ebJItmXI6U/QmmNc/dVjNwz1AKsYWS70LeD+Hb7SGV9XcZ+irOZYfPc7RlXro5
fP+UWroDaCbpZxSeB3Ztky0PB4oJB4WqLXCOHJAjit3yv1g1laHGyMtrFMxbISlN0iKa8vcP9zrW
DI5AKxKX2OjsRjLJIvKSXGVnOpIQE6JRNmsGcuIBJiJK+zn1WfN7xk8Skq77ZF9AhSpWI/F3b9OT
H8n3rlUxlI+IRkApl2lYdEkNIDNfwYL/uEbbgtKEQspB6ns19ETiz9RHiM1FKzE15BGiwjGGim6P
mQ/Eqi4k+9O0ip+U544JWZw3u+zKjG4bABzVH5ggCNVkuDztOMB0+29GOMm2eBGn3ndGwQOaUHHE
ze+fF5XI5J5bZEh6xyBI2/Zn77MVvMmr3Pvuyl7fUicVIiQGvxQEkSL4BQwmqwbdPh+2EaKSCtas
rwgj+NRuKrEONNY+3+rf5puKY20PMu3mxKas890LVQBP5iK4ukgWNNoWD+ZtDuVzPX5TXZVG7cux
B9EPo2tY8z+XIa3uAmzKYCI/uppdvBY1ErAmfTCrDpNJlYiXnQYSDNhhaphKRBXvgj7kcGxgklCl
/vA7pXeYu6bMzx60gkiPziiVz9pep878ayAV8EHxBPRB83pZX9ICaM6uKUxPtU7A6gaayZIylCuX
So902az6kcwkCeof0Q03jZ6YSyiKG3w4iJ9MI4z3i/gF7bNxLG2JAuiwFcXo1RNYBcYFH9ntC4VU
H4av2AembnN63sQCqujcGnePtanzvw5NT0ex8X7ePqhxkGhMxApCybSW67n6S5IwcKLwbs378Tni
0el8lSgG3JwQzovSrDr44ElSrHlNQ0TMum0EU4HlPS5yRsQj8wm3MzUqz8whNWYr8O04s9oV390I
Hwn1H4+nTB+dBSNlQOcG3kCmGYPt/WIPDAkfTwjaC0AUcgleiQwnd5MyThOHLczuRZWpQTvrHwoD
s8D8/i6EUwAcQkcxKw3sZcxWskiesvdFRG3r9C2yQHRAg1r9eYslIatVBEseFXL6I+q9tgAOOrfi
kJvl2OLoxs3Hl2QnXAKFkBAOaJWfCXhwkhYb59vyqlt9V7mJ9NPbwq6Pm1T7F2Awk4v/0sm8qY2y
WiH9OtYcNG80zRf0sWQt+IwsKZNP17wW5WX4zoSqrgWVvasoUhHR+eMoSN6lJinxBStR/Lo0/o/3
41wyg5bF7sCLGzeN7xi39UP9FKWTCX9BmM4Ja09coLZv3/tKP4rYL4lDUPTGozDrYQWH4eMgNH/m
9fcSBfPHGumHHRYiJC739bvnRqjsXfSUF3XV7mBKN7IrgWP+b22hzstUozVhoQUmMCnFKzHwTbT+
AQ2uMcELgJXSrFKkJHDxRm8q8Hz5vreUxdMUQaBPeBSIMrzma0HuawN5zToEnkL3ghtGa5h7IIQj
W2MWLhoCS11mtRheY+nolFnkhm97NEIeU1UJzcgAXdSnhiOHUiziydonRmFBssss6Wghyw24xnke
RPoL5BA8Ibk245ilVh7vFQxj0YH9o8DFir67wM8sRFwxiQ6ivZVdwFpVMjwdoSfjMOmJUQSYF5Mw
T8Wcb3XAQqX1ZVUPxXtbTGwGM+2+NbkC8Rh/I0s5hPgtIFC+hwdW2n99nVvt10cK3YBZiqDXhI3N
X8LCaX3wG8IFc2Jjg2Fw6dKnmgNE6dkNqJohN/6oXsy8lqhrXfQ//0UNJGAnetCVv7z10a4FO9fj
BbQ2LYDHAEPurjrteQHHPmHbC0NxiTT8+YAD/L+t7DnPBsZ6hlAoLjpAjKDM1K16g4XXTuU8G74b
WPiz2W0ywZaWiMTG5h0Di11ESTKVyXb/Yoysgj4ajprnoYXHm2rP2+JOvTxEtZ/DQ9w3wKHT+anK
fTldDdNkZNwa+OGE2ocAv6DRg5pgk+JtqdALkA1wnPWCdT1ZOv3iIhQHCkBFpsDByeiBP75HiMwq
H0maFK++hOun1gnwJTX2OrGgBw6yoFA3n6aB/ndzBp2v2PUxuilNakgtGPJ+xJeHupg8Mi+SVO8T
bx4qTl3bd3M6aPp7V6o4nm7h04Bj4/et7QdAYS8bT66BKfD3e/JAByT1JZWtN5hLeGl6XcfDHjfr
mZmL2yfLjk2nSIvJQak8Z+HBPm55lJpgpl/hzdVdPCigDA0tOItskqn9EeFRfu2gM1484fDlPvVj
fMMjz591zUQ8cCr9wJQZuuIhUHrefZlSfE5lToH4QXyaAKJiwehLgf1zAoS8zt/VK/oVqRUccFIs
4cpoAAUVh7e/skqBIjkDBNiPJH7VBM3IPGOr3x3VwXNBfi+bFRHeRQJJcXVPYD0Rip/nPETTEINe
IE5CKQU/RRlBpHG/edPMmZC5i7xUGaPp1dCO+xGver21GsrNUw6NHYeHVD8m5MZR8ezZ/X601DNI
XvpeZU3m/gXFUymCBwuslFMa8NOvUr0M3+rz2C/tLw1WWhOeKVUxhHenCzZ2Wy0/I0Z9HNvCF9cY
b5pm7AZagGMhUDKXLPnNKoBeKAs4CAbuMfGnggiV2IH3NDFYqD0G+MzGWwy60/59xrfVBOO2+8IJ
sBR55H6Y4L9HiRqfKiQKukvLbKwhiEN5w5FMfKtp/KttIS+DjN0H1WK7GU5sydkHQDwVpAKWUv39
f/mJBYXvK0V/H44SwR274Buiy4HBbbgundlpmEgBcEO+ZsGoiZZZXlvRBNNZDOPWGAS20IQmo2zX
dQVMep2uzQrrS9/kBiaX7qaoTLts6poMjpy7k50eltiVaWf6YxJ1MNhV71xF+WLsizNKMSQxuhha
mi6Py/agvPLzoVcW29cXAsVssDTXMW1MlpphJmXcJqkaKXTfZPAUa8tkYZE5kv5IqlwrTWZ0hCnS
I9itH3lTkim9n9OIZD7DiDHnQk2kvaWiRC8JRJP2hWkCmyjR8msu6HuX7IQsiKfLWsxztwlh+d4c
yNCQvhmdSJAhn2ba6+xR9DcT02UgFH1/2xingckg4kyyBjj2W8tWve8vJyVLqjRTe6sj7BGCzpKp
bF119vfTNixAOLt7FFqgX57wC8jh6Bflyl1rVS6kOgezYUb3tfLGZ4dirZfvY/lmPz8MifAWaOs4
RMOJN9DzFVLKWlTTp3pmIuOFzmd2m/w2MnobDzFL2o3kxz0iNetl+0yAogQeI5fzfnbPn0g5dKSC
+KYUYcmQCk3U1FYJiX4pRM7d35PjvXAgzZSXLpxshkr97OLSv0WBMqBY+C4wLNirhGDP68WMzNHF
a5TOmiJQrwK6zkW5Dz55k+84LsDmPuB0J0KU56CkpIFKw6dm9uxhQwEt3YWtS2dOoBX4wDbxAPM3
4Vy/DWL1S5I0YnuwpW0u/oKLfF9fXmT8lWw84tzauLVzc5RavTgneBo2bcz12wf83TjI5Tk42KPC
1IievrZJZ4bRVD5Y3sf6Nh5MvjxzIro6Cqs6iEXHhCnpadzoqJSvxBbStkDToztMJKHjnw0Uvixe
G3C+WFxRant7rJMQLQLPz4/McaxzLcVn0DgqD0CZ+09H4mU74kC4d9d3t1pW/VzoHm15sW7hpU1y
+tKfXdZ8IK9QYcUiAbJRKcSFn3lrDdeO73GwxW+rcNULGAYZ1GAr0ZV9pWdmpvO55tFjK8vFMBp1
+NNblUJLudjPMSYvvTtS+UvYKSSF4gYpn7tZY7Q0M16sndgR3G5ZOzwCy5+UJdPMH2tc60v7P26l
CJoeG+ztt42lrxSSC8jFi9sFhR1oOzy2VI1n3vP/ZYjsW52hDUerdM/vHPQ6w8CPfm4ryuA1rE0D
K0yvg1agso2zXz44FjIW5FkZ7A3SGEXUGuQiidUOCEH4DpmIBYrWIFYZEzOQcpIWqDcRgEDNuKkS
ZWKA9hiIzOxcf1wlcfHLYCJB5saXaeHDWpc5ZAV4upJaThf2dXWBq5ha2gxibDq3v1oLVdQwzfO7
V6UoIRA6Q0ZFaThzZ1qDTj46CXk0974nQUNTdnjyK0Vf4SsKC8giR59ZpllbnWcN/b0Z+uHTuFFz
hKYEd/qW2I8+/EnRGPI6HBbCg5Lfwilh3w75szcCL1fECN3fBkGkSvFbyqMmBKwwWClcierz7mYw
QCafI3ZhVkuCudxm2+KutLJbxYOW3WrWOCzgxdz3z8CBd5vXIIQ4WSvEFC7/VonJ9km7Ie0+WQf6
OMd49VYcjn9s0Y/Td3HRRxBCDo9aqSUyL8MJbBKmQapQ72PmKyk+jraQpFZfZOuC5xHUlOO0pMNw
57xkFO4OYIBf1D33cHF5QmAk9EXZbGVjX//6mh1Lbo7GjHQ5YylX1yiIGdmm0OzALdu2C0Wvt08b
HJ9PsNtQEjXK85dKpIAXMcyBu3vr1KnRrvy5rJ02ERLwFlva3v6LuM7eC1jZ5No02KGnbhyslCa+
3mnZQD5XV8c4glerOfbIqXUCXbNRzKbTmcE6vBguSxLmDaEo2w2qaegev2ITeSduJykjRuO2rI54
4/yf3NR5kWvp2enNzJVKmVFNAbI627vlxQUyGmkQ2ujYjQoc6jUpkBNIJKx2czX22diJjcAWgTqF
d39VjBFuMN+mqtNszloetc6+C+LaBC9pSVBHqQ7hPFBufLjcYdT2bJVNyNAwnxTN9RmckhH53DUw
RcREl2DA5aXmNDb8/GuzTXG7eCGNJpRZxQm8sGeasgJSi4pFEotFCvSwfZ4M5Hrc55ZizOpljVF0
e+Ua2ZCo7133KDa4+zWOUwzIHJIfXwA/GGcXhxuz2D8bQY7oIcmLDevTwzFueklpu2NZYIUKpMsZ
+HHctzOfkqFfZIZab4dUYdSDfPwlRFar49DbcLOl5g8aT9RNPgBxIslKzjhhXSBh/N97GXdyfMEM
WRYuinSRVrvFWQsYcuUu/QE2NWO0YgOIGaELSHjQ3Fj26xbKJqmuMiT4njYSY+5UehqZCCsxkNNO
2y+y0dv2Pc+/B5sb6RwY6ErKJvHHRYNaTF29b0UKbLEfBhiWZtTge50OLfHOnD07DfX2svn+BDRK
5Upacm35Mg0+yG8IH6PiuS7HJablyOR0mcrTQgBdbzM4a/HeyLE8MVWJ8u/ZtDvlboFXzyNndq+w
vZWWsnrQfSK5b00qohXLSD+EpmFaNhQLfOOjxX2gIhiFPcbTlaNsqBi0IKN5vLwDUMlcrYnV9GZ1
5v4wqkfoEPNTXekHI2OGDZoVf8TMbnJf10gzogLUtIhXM4EFXt+Vu7YMXciWrO8P4602qVKyAmaB
M99nuNRILWpKemAu7Fjm19NkrlViOSWu+m5Be3WiEcVToivX6ZDdeeDyCOK/hPvjDaLRqo/GBEmU
W+7sUwYlkRmGDEXQcpF6RsdWNs9x+5J3ISr4fS9mvHgcSUu1E+rpvyUclNvTUGj6T2v9Hqk3HClP
dN/EmD0L8Jh2jsM93Z/6NTCxQv9Sp0uOVm3ZJX00okavgM9iRct+UxkzEsvAKR/Kppx0i2LXlsCm
pMm1SDwb3T5ai1o31DW4JLkJnHCECWjFXV1h62tGoTPCx5ZjTbdWWPoDHeJcj0aIri+ySjds0sDF
7WQRPlfBB8Su16GEwhj0lNIrR48eEJRMo3MUzxjK4qX6zK8KV+EyGqV6fPKq5Sh2n4INGGPwF0xG
Rv0M5AJeq9GkY3Oh2/jSdcnOL13CnHgUiCdla0CEvqUaCm0idKdaQ906rNY//YbLqNKOo56P6lu9
PjmLT0SEGBHRO8Po/JRAe4dYP2NxHtDEknw2dcNLewvk/fn5Yn+ZVPheTJxs8ShVe/PTPTfzZ+Q1
WlCDiY325VYSWY/x1KQyEpbGtMXYzc5417RqlxRr0sRdgHJBkzGbl4jLmo1nxmkT6RsRe0vuCdt3
vROqbq5AHhZxHay2LPhLVMKYJtmBn6UWd2fN9MgmUYoLjXsBv1DfJIgYOLCzOmhOBsSC2yt7oYJ0
X79WsuEp3/+7sO4IRp9r7bBoYv5wLs3KKQ2lgcsXXKyaQd5OiFmWmYHJ7t7fS9icehfHRDiK2zzd
o6ejwZFEw+UG0ffeIOYKam83hkJ8ZNTGGZyKvpDAPmn57ERRtVJYxgLTOANifggTqadbGjHvNfDu
1q/NcOCCTXUaU6JxrtQ6WSYEsAht7F+Y6zqOpvQvkNpmxzpupnwQ7p/JWDRmufx2OHXHymtG2+Fi
GpPoLXarFAXVLxmbmWcRKP1WCDy77I4z6KJcGubOv0uk6vcpaza9DbKEdCE/YVrXhI9Tnxu/oZUK
//3lB35/+zEb0CChwjHKUGVtfbhGlYbh7NO0kHqsapY7NqwQhQCgAgn4BSEJnpTYO8FO7E3GlPNR
DDAf1KclIk/uKMqv9KW3Y6jTy9ad1dmEmh3qVdlIKKDeW1sg00p3yXWjt5Ucj7Z93SW0Xdh+DVi7
cdZitweAV+7buezO8vBVIEE/IzW53/1FyQsvahRCyg7ssKD1IEQFSzTrO8oe9z44rOYPr7QkkoMZ
m5eDoXSqOrk3EcXdJqci+ggDdS1deAAEHpCkd/XEz4whXxHVjXIiqcy3TpOWbFaWNI64BLl2tzqq
mJYPe+2I6yXDrQjC6tEZhqL29susDvF3bHzq8lSTIwJA5h62RAH9At5ELp3MVv7ZWaKfpfUv1neN
8/UpaRDrMKcH6qCQPh3/MUWvzPBUULeqPJ7zEtoG9f5SgcuZ/r3/fpGlMfbWgsjaZd2+KbfyTGb/
csB29SbNN8PpTryKKqCvmnO4XDZagUgTMWjEItroHTWTqUsWrw7ZvtNXzgrP9RKRo2rHNqTU7Btw
u/hgOAJr5Awyz406UFssrmQkdVRvyT7hpSvm35zif0s3uRF5LJV9jUyu/TcwYYBLlMjeKFFvjjVS
2GcL+pmul8t9TPDrAWhy4RrVbflQ77Vq5TC1pyZo/sicO7QEMDPJPC1XI3uXEMrGIPadnwjEPOLE
xmmetKDhQ9X++AgBW5zsP5lVsFC3+AtqdEURfTb7ZBHGjeHdsfyTjqtXwy/tOjxNu+Q1cayi/NPV
ivac1RxgdaPH45pkP/hFuo1Yqw+i7jU2U+HGxWrl5z+bxku0dgnJIBEPzQDwx1YfsqTUAYvxYL3O
p8xMQFIsixCBL1fz4uAKzZU4j8UpGt0prKOzMXAtWBhpaLBfbeIh7Pf3fYe+5XyPtXomTvkkz4fl
n5WPmw/b0dB07O6gSTVwIZ5EHPXgXKiKy54qvzgpgIPhaDRxU3Y5zdjtWmg6C/Rj1mWcbT4ZDqZ9
ftH/N0O3KInIm9hSJRm2gB5vTYVjuTqkAg8Xfe998c+J6PjdgAQ6G8ojPw7nQquiPSsh79l25kza
1wyxSqgwsO4orzXr2SUhMyY2otjP2yHT9PCw0oWxlNS/81D2ptoSOe1HDsdZNtscPHzz5AgAvJ+F
ob9GIKXeYazz99yqM1PhD6YAV5G7TbhELpxKzYovzd4fMwV7Kkwc30ZBpS/LV4Qua+B1VvD6UYzx
4EVTrPQD2RaXqykMAEnKqtdEEWGAad+329FibWhaR38PUIrcQmO4ror1ZzE0ledV9aq/6DZsp9ke
22z9fg33SSTnGUVAZlvA/6T5uS+Ztoce6lZJ6k7onhC/slJlLTnn0LvKVZ1Hw0/r1gccty5/T+xi
xho1xk9va8Fe14ckx08G4L06QqMf6VqjvHuMzSgIJWdSJI2av9BMDKjX/z6XyALCWptq3nPiSAbJ
OYqrpzvUGaRSS8+0moq58PCIApXGky99/WH2dbKIzl+Lr0sdObWMLi8z1A1UBE2+vjoCK0jg7uRE
HkC9qLR0v6Vh6b5auzFbWsWV5rzp/hP5oql0UEiIn99nf2sjTH5QOesHlyAnXgT8jawPxPppanfA
vf9/Nt1+HXyfDaQjkOtzPT7KSq7dqaCg7Rj+2Ns3cGpVI8Q0G7Pe5Lw+zcn0cifv5lcThZeE8WJZ
XIf+/6UZpSHSwrd2SzLCv2sN/wgJNRJon9e6/Pd6OXDZQFidlxKF6NnesXDcWic5+8SGzHPYnwg0
8tJ6bYJD4Zc6nPcXUBFWbit6keCFLTXrxy/eh+Vvu+KCFGthCseOXC+4Oxha0c1iQwNUUDcWEylf
RyDh3xgyJ9+oCSdYaHACSXHeq2I6TSqMeKlofh598cjy+eCJS9lpJRobV9uhGTxV1D0Z5o3paqUv
KXzP9CxBQaijzxdKgK4ppk0gXMLaYlhbr9Wa3NtbdVezAv5yfxoavhrC52XujNBkEGza/MYHmEcF
e5dCGnR2NOW0B4NRWQnmZCMAZPsxYTgcYDZTxhSSEEUrPB1dGiDPtsk2K76oquSUgLPR8dKEBbNf
hmwUNOW8//Os6v+dWs5E13seqB9FuG6S6YqATyumgE2b86oowIV6Jgatix24/ytkLOJ0M48CUyja
rbi7xT8CjrYPQhocPYwt/SAon4k1As4GjxrvdfbtWt2Cf3yfvZJXlYL39HxCST4tA5E5grSkAg0m
oiKggZ6SpQO2/LjErOnyG4MRbnZaL/HYo0KtAxCTKa+T3KPWaDikkHU36SIjLNffV2DicSzCIfEj
IacTshLippFRWhmGuIsUQlawPhHg0Vve/BGWnAfVh0o/QOBgg0qxczSxgW0BzGMjO1DvC+b2RMWs
6Tu785Mqmz6MeT50RVyBRCIqZsFjfMGAAt8lvAV2/8Y1XuAUbaD6cBb7O/Xjlm1dnKRsbBG43Zyr
tlLb/QthQ7UeZhBj69+VeVXlrVp29GehQEsm+DF+VNaasdnVCZhNBDdie9qoxDsmLbjpRiN2tWQd
0ZovYZ/1+6B+OFesU8Pe3xL78o/GMIzAaAvpJhP8tYlAiSQRVhumDLPFGoO8jEa6JTdTEaoe2aNk
0yUP2JsLjTzj0Xqh9UtMR3brTB1lup0NlPsPA/NM0+kZk9WO4D/clWAtDGScvxEAFxUboH72nztQ
Z4BwdpzZ5GuQhqWYWZvrMev4jpU/vB301sq4kKzsqBmvQGwkHx/RTCL7TgegogXV6QbhpWMOP54o
7JvN16nXXoIhqLYmzpK5X+c9IGzOD2hotAas70T38CdzPfuPeyGklXlco5q5Sp57E99fWAOGq5S/
78OYEdiRmKax52Dsla+Gn/mSaSTFM4AjLB8RRMYcbdAioOlB/xXQ7sqH5C3s129oEWj1jmT8E8Lo
g2Y5b7kc+xzg86Zqqo+gBjK1dTtbDflJ/ZLtwL+Tw3ppF/ADs0cN0YExuF9XaEQ/DB1CSK67MrEZ
2h1bOeF8AZgJ2m7LRRskgGH5uM3tddaS4497OFfyUrjCgnotMfX1gXzYBtNAQ6Zuypf7Vubz61+Z
5rRKqsccve3Rwacfm48R2hi5uLtp4m4Y7R66qKd32zlav92P4ebS9uKTygIRKzo30OJxKgSRBuB2
kKIthkw9+lmXAexKF9+nasAjoLzs+9YCmZp9NO6jYVCaNPko/yyTpbJ/y9+r5Mr5WdDZoZJZXjqt
L6GhxmicKBvgDH9Qu13NRaxbV8A6C+0qCc/oBMrsORMY3xymXurzPdCOcH/f9JCd9WqRYkzLrbkz
xZvw4npZ8a9YTry3waBqL1dTtRw3rNcVyIdrzMnM5dGw77CmM+tUWBkMJryP11juCip0Lsl1Y5uh
r+TDEdsbbl1N10IqsjP3nSuAj/bfCzkw9tXJC5xcM7lHX0jbmg+8BD+ReXv/hVZopDC5HROcyhjZ
rGB2SPhtH5DEqcPe4Zfho0PZTwDYkFs5GDsQrBZvsPyYWfhUzkN0aKQr4Gyw1CcWD2kZqn+dMO/4
1SQPKZHjPwVLnFQvR9mRHvsb175+szKml8pKT3+raGayNbQyke7l0jWNqUVsqHiEl/iYFsq4H9i/
5ev5i8gYh/Qh2Y+esWN2JXndKX8vdLg+FJDWQYty/uJLHP7sjwSSvWXd3pdIp2XxPi4SKA6ia+FY
HEp1jxMPItpBlGUz3UnnN5p67N/X3+63Z17sn1ucarMJ4g7PJZuS0ME399C44w4lgI/M6boTtQE1
DTvRPtROLI/ivSOVecqz/UTAPsvDBLk1Af/LKoVqfNdGgLohZ7DUhM48P2tcrzmrmBsYpcNt/qNa
UsXOJxMsosHUkZdvzDR3MBsKVH2CLH0czHV1xxe1hev6gaV3RIrsK68TLZbySZwnfdOfBE4SVinJ
jkQVlIvPNT0Q9EFXPF6vrzcKmegxNkB3WTMxg5JJTRhJYw7/fRbkte0dhIt7GMpSGatOl2tdKVwZ
yxdQQ4ulOkBR+CeYj0o1OiC5mWn4yrPkWGvxq6X4ztEcjiLS8HNjpzeUnVWxiIbedOmA1qM7d8Nd
DYCvWKyD9XYKf/oBH+AijganSKKjpUL+aFPdxAuIKH7+Ds7dm63DiWmQfVyTJy3Jp4DNj4yUMOjD
wwSmXAhiYCYDKfLY/6y4Iht8njoWgTRxtLetcBFVCbHuxrz/oOtf6Dm6I/Ewx7NXJxHHvXlhzI7f
BoSwdh2OD/O0tbZXvpKvC7GQOM+rvIgRf1Yy2lrTx6LIzf1Av8e02mmyLavxD9vPqHdWXdK0UMCn
/nPuZMXC9utZEr1YdIA9wdkMbAZ4MfNo8RgkIXcME4EdtHmwsivXsettCpCWlznEE3uE2m8PMvqG
OIXaawHyiOKYQSogZtfFYqfDwhhLT88hV1U6YopJiF4xpZfDQ6m+8SYYF26ZMgQFYFpPq8Npo56h
FKcNWi2Qi7hViMEN9BiDZHHEV+Ux5eRYu3c6sylIPXvSFalarPRQCl6qUGYzKzKDCoUU5JeT+CAo
0xDa4v5pmw3NeaRenBXtEuXlcSTfXdV98xOup+oaeFdc8A+AqMPNkni01APef7ma24h9er2tyWt+
pqMMpsiarXIVHuWoGjk0qD4qQvDdyOWwh/EP9jjF0XbxeGXML0NtDvAKYdvjqy6LWMDsu6kw3/uY
rBLVGB5z0bNJjY2m+48Khb3AEl8XpXjn40Jk/kypsA64RE7buX/8BW7en/LNNrY8Q88LZlRq8iPf
GwPbc8DnsZGEOYNujklG7PbQDNmjRwY9TVwGd2a5WWsRscI+VG5I+B8Kd14r/ioOKJVtIrLCuz8t
P2bkQ1ZBmnwcnMkjUoCwwqMY8WmoJhb9/04zqszLyn1gXZwly0USDetARM9aXJE56WxI+PyyAp2M
8LBEXiy9OysNLYq9zYQLCGvdkNs09ZSTGaEYU3NeRhFCkVvAlxvfyvj6dPeQRO1VoHl/WmicqQTd
mCykMJw4EZqXnOjsWWxRmSXFhfUnfrnT5oiv5LdoSxb5m8Q4WtHqbLyDmN/PrYyP4G4c9Xpz4VDe
ZqGfvxN2EkzFxOXp89We/9/kb9PRH3An5Msq5CxYvcF+zBU5RD9NRfRX95mhFE4Ii6+eCoZ3Vcvt
TlP6HwZpdxfqofXtguhjcZq1Lkuk9XKVTmceATql8yyhdY9x3Icn7uXU8maKvpv/3jZBQ2UkQMrD
0WclqiHpcYZmu+czFEqG/B/yIgTSjbN1Lzwu4PY/DQF1cIGFO3BpB/OOune0ElonKrf8pcse7f+p
VCy4l888ZOCjnyuNwAOZWzPIqMPsrwsJw6RUltMPE6pVMEY8V8BihwQJLeQ2MhxI6ghuxJm2jBlg
So4l8jnG+UmpFKy+yyHNaYIB+t6STUISPF4Ya/E7oydrEUxfP/FiEz5sSlNrh5ubpiHkrEz66hOl
j56JFloH3MZNV0Nl4OPhNF7r1mnCHPe/yEbcquA3CIs2QIoIRMIQcSVPi6vDaeQ984oe7RdNqtp8
12AO7YIFjNwE4uWKFd/U7kd4vZ8snYcHbLgF1MkrmiZl+ul8JfjgaHj3UhTtziUX76EE7bXnv/VV
9GOizHtSobzI4EghKoPL0DYvFDDCbbOBylcN2Adc7mpib++L7Tj+wvY5n+P+8QhowOxc2BuI0xFl
5kee5/FH82tEH70+RAybMl7KaXo581WQGJ2OVjFYGQS26lud6X5c7Zz6ZtAfW1h615/vkRs0bKMk
q8Ihj+m55ocowActToCgc3yFPtl1uDO1hxDP8NCY2OQfhAqvvWOcfSNi0chsusN+37pUe/29a4Fb
Hsxqz6eF2EE6prA9KkOHBebGC4Xh6WxI7FO6pqJ+ViL+9ICTJsEQCxTGWnjgSQRHwMgRBDwyhu9/
uAM28txTwUkoRiqfERmF4uKIm3U/VkNcxdzXgEgYuphbgelNVmA/lICh7lCPqQDhgJP0UD2bp7jq
fJEhAQFsFmWVKgmr+kqQHb9ySfrrkyON4tUIudl7eXWQouHABqHso6aytE+o5LtJVpIHYSaEC26k
hsg7Q3+Zw3omwKlEcehnANX0tnTH9zvnPDgWDI7tOWFtAoT19n8ySuRn0V9jlF5jN6/OGEhb6cm8
uLdKxBSZUdsgdfYcPi2Y/IUfJXDMPwndYpLEcnwVPab7TnyfQUPFug16p6REZAkyB7ouqLBWzwGQ
2hcUMQReqSubfsKk4y2ektSW5wnh7prC+5mpgDhfepPYmGvkFYcgw/RSxm6G9UFl5tfqruNBvmfa
geFv20yIw2OrMliOvEd5KJM2SiH2hKWaa3O3P+9TX5J34+ylXRa8E5DlcxK9kZWaqJz8cPT/8zS3
0YczkeRu/F/IvVzW+6S9RDORTt0kuoQmY3n1vOgLSFVBpkp3DteMF/c329RK/ysRAQznPgrDG6mz
RqiyYAPMv9k5fO1kY8lzmOCyF5NJ/46bIosTzS0gfiaN0YX4R3i1BBXUyJe+XWBXPzfWrg+AM3e8
EIsCL9AbfUbANC9DXMiBt9GJDFgYj2etr9bY9VOGiESHPz6PGkT+dLv+fPg1/SPmNEHFqq0pJeoP
uoM5iFikFbrckQbS4qYKR4QBTUf2TJ1lZnrIfIAg+v48tt6W8sKxK8+jiKPC0UmnOIroabJ2UuU0
UuynVjFxsOKdxx3wz/pz5J3LVl1z3EG+UEym7qHJkZYj9WzrXseib1Q1hCq979AQylDw26AcfXId
gduM0h8YMOE99qqBKDDIcOi6nsoWr9kTuMfTiZKxh7fdMKfmMHGY4b99GqORIyFCW8e8C2JT2Y+c
ujG5Q4pU0s8fJ49u3q4Tflb5wspYM36ULandCQZF/xw+ZYkMZAhtdT6RxOypIjAeAYBM9P2WBdpV
ORt1GdYhx4BcKQgd1DpSNljXAfQdt35l13d2k15Gdka0LfeiVhLZQHR0rOS2IrIGAcK8RPxGZVh2
p1vYlBeYjGTZtLuk9Q8oURACSMYQ6NcXSB2znKQNmjXRklUPz2sr5A5zZG8kXkqmfCOynThlA7Ht
6okF1rRd43BagposZkIR4U70ZrcSkkrFI9tyaDEYLPiXBD8tu3HwFCs9QD65wDeA1QHwJxWvN27e
i7ffyLTcajwEOsYR9wNRBqmYDQ+t0vw45tW/GYh3ogclH/BxmkEgM6g/Uro97TsQLYiN3XHyi4wN
EeEaz+yzZMSZS8lKF+4JByxDTBg8u7eVXVAtjh15D1PUOL7E/eHskk6UV4pcBq3JBdw0ju/7S8Vx
AucdVf8AQs4CNdLgy/AkeuOwd7lyLr9FBDvlKmi2mdzu8raWReU+78bYAmnOfj390SJwebtcKAQL
SvTLmWwXsRPlq06YJjW2rxkZKcSlPgXR20MudbJIp7HDzf1mJnxbm3k4OQMtonityHSk0zEESbWd
3BSjtCtBKNPl7JfS2MU6+Ead2XrDM70UiFOkvZkD/1CL6xlNkqwWJmzBnam2DTVtDZiLX1Kk6kGg
Di772jdVq2svL1Dl8hW7U84gzWgmecBcvh7a0BoRtg+TRGL5WMRj8CE34yzSb7ahAo5QQZsA9R3Q
1p2eoC14tJ3PpGNB/5P164/vJWcKOkFlUVQxawJUIQCEv90eSFEjct62D6Td0TMwW/FFh5yqW/r3
oSYhGwSlXreI8WR/smudo2cjCiDCjfA3K8x+Ibb1h7enKd66fTs6TS8+VhCbfY2sLngKo+eNEm4R
umYMKshUyoZf7v6Q8KhiIfHQloBfnxsrtFPP/WqFZbDVegZQyfywkiYIpDJB706VMpS4pp9HojJe
7AjH6a7CoehqG+41s55bzQlVaqwhVqXo+zfLCKEHvwCz4oFoQCNjk0D+TBzHqJ0elJimndsJwA4l
FbAln/nTuZFQcZSIKap/FxbUJGon7jLciD7vGPTKYYkUUS1IC8XOkwrZ+8jexysQ2CVO30HTjZ8d
OttilkxI0CPJGCTmusWjrBWkWJdKGK7yriObNPdxTAhViup0kO4V3wzSU97qdRDUGpysifI2ovcf
o1nv66QDXmY1+gzk8CHPcyY+u8eDvgjyg4gM6THv+4d4CfaQeBoPrKl4W6qo8hM1M9Q3N80RUjwF
NJwllmDlq0a3jJYE8c8QfKpjGtJ1fElPqY4RTeap6S+Zu8oOo4EDzXY/SsndtdjVsay6zvyWP7+D
9CcQyq7i3rudPSh4ePeQJ+VmbaCD3GBtZc0O7AiSclzARhcC3+sSuA3xm/aT4RSJfyW03A8pw9Vw
k0Mlr20WKtmavTz09J6sNoo/BSEY/LFGtXGsa9WhDTn9Z7MIFWlB24eSyxqm57rjZDkYvclOEJId
Jrv2qmZCKaVuPjq4N9AH8zY5vvEDbG4gCVmfoXcp3A3hLeRZtAxoqSKH+VITZB5x3ttg5a7rLQn/
8yhho7xwHettjrH/3bSd/KfhbH8nXqFMEKU7qJdC50P3BsvxxQzfvTmBkcll4siIkr1kZDsJaFBg
uOANdE0J4FoEP6YWH/TZNX5wB+/La0xuKrZF7vpxhmTK44H85iuCYAkX46qy8VSv91udZzBrOshV
HUriMiB47K5myoDRWLyp9mY9DB0BEvkcw0Aepr0nzdiCzWIndzj9XqJ+cuSeKkjdVXRoSKMh5ddG
OIi421duYkXTq7u3q8zM4yWHoZb8WaD9H4ucD8XyPX561JG3mUg63MhLZRuYBHFtRQ0drhf3Aq0Z
De7zaVT/oHB3yxsDbCVKdkmKqtqMFxL8Z+ayG66/T3O47Hm8Q40TtuLF+58GjMyF0rb3lJtW11ku
hte6WScXiJZRtpYKJ9hB+JbRYfPSjOdS6wU+rR7kUDh8XkBqDoe8NO0p79Io+HBl6Nb/j11mG/Qa
QAA7hMaKK2Ei1eRgSom6j6INx1aGUnMMYZTG/j83QZadRJ/5tphBs9FhSY3Cs064VYHv5nUN49z1
hijvGJMPezdN/cZYn1Br46svyZW1OTfbfSN61Z2EgAqNxem22WrJOM0ZHAiJGjlmHsyXBLffnoH2
XHvdF9vvrGb9py8YhcHxrizJnlrZ+RM5a45D2HSAJ0aB0eiwNY4cSsqdTK2O7EP8PrCZzX1QpSdV
Kr9ePqW810ZFLPGpKhtWvH+wWt4ycRIEgLtofda3MvBTuci9HLtoUzbLiok8ZJtxbTHfYwPovlp/
obl+Un+u0KiOi2L6andcDRWqyXhv4VNsAF13CMQ+CcvyJc3ppjxvQ4d2G3jjoyaRcK7SxFtx5zPS
2xVsD1h57fiKWuLeVnpnI1UcDLiQxcEzJ6c9jQgJn8Q9vGbQzGDnR5zmyEjTIuhwtkSPDE0Mx9Zc
4hiaN7L1lC2prPW3knVmEVPaF1R8RrKsow4bQL0vvdySMUo+C92s9TIqchdUY+oYkNObO7ytAVNx
Jxay1rEY6d7qtc4SnQl2Fh2kZAXea0ESFZriRExV6eWOh2Se2joDOw6SlExBlQHMnIFqiSJhki3y
UHBprytUf5MciHpm/jwK44jDnLhZRKru1QI9HB8wCppqiSb4AP9Me3ZR0Ni7XsAfFs1LqDnZ7HIh
zAp03haQjUeGrsahB3QTJJNMucNg8KrRVV2a2Y/kCKHH6jffO7Vm4t6gOzQyQoP7E0mbrEax13FM
NgGdSw0nuALOyW+nnI7l6x7c0jDGzpIq9sXn9swBHPFxAHz6lDt+6FlpMH3wDrODtFAUJAavTzGB
Nun2RB8A2OQlbw72+3sqrD4PQISWHTRkpUrqPObiCnAH1bDeeBeh8vXP9G3ST1kKNdhNz/DcYza/
QdGfXgzwTlaJb2t5LRW6rd46cP1ncPxRl0MwhzRw2yPyu40cL2SwzRp4s6sw0P4GIQOQ1nWBxDET
hdWz4vOjhIsOYvbfXgZQo1/+p6FCdXlTDQcniJnzJyOctO8FDeQT6RPOXrC658+SNHoD+AuCcIJo
khH4b9/DG5aQn4JQJx19r4JRzrSEDDw0AE8QrTOx52v1HGZ8YFv1qsfYORbC+1NLBTIBvwSAhyvc
KOdjc3D5TaBn7rFOYbTMjv53x3LvqFbnkltfY8X8WNKuZR1qah3V2yPyNwKZ1DZbBGJI+MQUKL32
qk3gcQNnSf01bkXvDyC6PuQHv1WMXYyC/S2x5iQomdb5B84ilzDmtInKBHtco0ud2wJ7lMHuuKdH
ywF1JjyxnKuwrLqGtagr2W7XTGnb1yKQ2mhLqQXSYC8rdjLOQ4FlmnLu/FVvkcSLXigpvNWAy6nf
iGz7ni4H4tenq1ALPCQqznlCsMGfFwicreOy8hHxAY/P3fo5ytNaRrof5GyWr/071A95TUnrjZJl
A974e30TlpiA2XHXdls9lMa2HnQlK/fUGbJazBOu6lgO/GZ8dmTAX76zulyTTfECb84R9KVkpNUp
8aIRA46CRSfI/L9oj0fkdTeI8710w1l1NH/BHysyS/Jv+nEn7BqqevLdD56z7vtrV2yN2mTZoEuk
T1Ik6AZoiaL8j7qEoUYbyDCOenOLxC3hvhPVmBX7KmZMDHQfKHAeDiaEzNNAliEufp25GqwwUFrY
of+7MAxZreWCAHLpZLDKOD4xJNRwo5xiRdZEiohs2wVtlJwu65VnSslG1+yD2fKgu8+RroiZRKdH
4g+eJYMbHIJ25zj2UDYSIQC8HUwKGg2tC4O6dnSPhfGR3Twnom0FBOenKZUU2KtrsvMXh97S6rXY
3AyVZ3q/GFe5dcIOFNYRQ1ALyTEO5eOEeeZAboULcgqMdhwNGfs0RIYVAENG44ag1V2kpXXU5HDv
rnfDdmqEKhwVVAjEQ6ZxlFWEP+480aeSzEAdY1BNYAvS9NtAGcGy9mQgldzD8/70dIYE2tcR5VBx
og00G2yjZk15mYdMkn3s4kgOO4a2OsNZiVkiz5w9j1GT2yZW6t0bbfMcDw18zHA+TagQduKRkDRe
GCo0QDAUjkmA1wRWwFy8bmRONgw3U5C8oSWt64ehvfkknazCTF6CVLA91+j56JbCZDUJ0g+islem
2NHIFDR7HPONyUZmGZrOWA02fNyTdbsbhCg2oVJ1bKMSoNxwzOQObzztTV5ZaL9+Gv2P7bwWKIb+
C4Yrug13Ez3MOzdHo+uQAwOkmIasleDJSdD8XzLqDQL8de39yaR9nRQV/Id0ao4XFyJ6Cj0jACKE
5uuWluMhEWbLn84A5jSga4Avg3QUEMg3yJwGRvNhQWeXnEmbiXcx30sXOjEC9AJuTKGxrO28VXoA
D3cctshSg2nJBJPftXwItbnEEVGFV1D59qR43FAEgUkZGjs2Z7pfD0Y4YtSi9FIphOXAIJqtbBCh
e2V+gNOX1WRRaWHvPHeBD+7+/CRkB4rCfuglVX1kXLU7BbL2wfjLn+o4Dl/hVRAHoBOq1lP5WsjD
w/cYt5nwbcBmLHM9nYhGYR4B8wd7mIr/HOA2T9RosmUrx28dRq2YQiW7pQSHFoyDzq1QWmFFhc8y
GrLUOnWamdZ4f9Js6e2s3uICjm3bHTa5jdVSQt3M16leYNw2CPnLBIaKb0a3DzEQNlKkIr3/Jt1g
uXpX+rmKwRdLTsNNK/fgqWsdDv88HgNr71f5NimRKbfq/Bs+j6tWjOfTODbY3evZmSI/pVwSm/w8
B+dSWQYMfx/HwqCAzfAbIlw0oK/fbWCfmsl8wbU772U/KM8iftgEoGh57WDZz/Do3JXXb/4kQfGJ
WIzyTvbUBHbY+1MSO1V4uAPHlOJGslwPNt7d+V5DF3VRtRbBpidhUGUon2FvB+9xdSEvR50BZQ/4
ZLFEV9KU8IuivozbVbjdVfzhVMrkfGnYv2ONPLJpwe00LMv0ylVZ5g1Q3Jh7XVIztALtvJr71t1W
c4V1YTU51cIMOxtWeHXECgwEbZUxG+zn4hpdqbnNwWumK63xg7SrQgU00gW1Wl2EyzmYmd8VKETg
Sbe1u7arfrcDlQQwWRb0Stc27VbLhM6YfdYHjQJyzxte7F7eZ9ws4UOD1R5gwoia1lPGiUnfI6ND
NRzhAVFnd8uDnh6O1S7U6kBE89zGizU7zSzSu++QZi1mfWsc2uEzFzjAY2g08K+9fbPAnv4b54K8
67qw4Ftlt+LPqW6NWGsRv+BDBPW94cZrDhdY3TYlb22lFl3uuq4GPG3J8Dqc4w9/xtbv08y8uBr9
CctcLfEHrPHuAO1YafBDX86CqWIw8XiDyqk3+a0NnrMv2RHYqTYQs+W5nnJGGSuWQdz3nUMywfR3
/hPWBUfQLzQfsidmAge3TUfWFo1nKWGIg3I4RfgQGTKvqOMNtIhCHYrLPLbe2qUjBx0FAMXkZJBb
d4+1ON8ftJsVV0ujgs0dmc666WrYv8XKOrqonilREjMCdgBzYDsJWeadqqyu4q2ybvE/OwTx7aIB
z8jiNVEzn6Hx51h2HQX15FuUkWi6GHqQ18OIkkjc2SPRNmmFryM0gagUbj43u5Twp0sIIQHsbuoo
fRzvkkdEgo0zQB9tfHHcAV8SIoj5PKD+hN4l3cFCYuWhWXtqEpyOO5f3GluMUIWZ2QFnmqTVwgXz
yitPwkNSZG0GVuDqX4SAMy2v8OyAvVc5i8Z5Qleg3g/03LGZBVUQLUnEt7YUu9g+dPSX6f67rwvc
8RnfseTMZtERGBbKvo1ikEn2T9OpyS7dmMId5XBisJOq1mUx0ZUgLQ1ECPjtwECA6kaf4BrKrASE
e3389fcdI2j0+AvDCeogjd5vYm08q1UkNsbWmj9R3DY+lYEZGmrLyjxzdbPET4ksFKaqnz+gBQa6
mwDuDVeEUKOtAwpW2mS1jGu/V34qAebhIMiamXucjQqgMkCt38+ZdmaadzF8rcvJQRxNDWaHSx6L
KLn12DV/mHGIQ1BAOvssJiFPZmx5tYkLVOqgRKnuppofOptnyGynkhMZ7Sbs2WZNcb9Ag0elkpcI
YSaYfLiqsHs9VjUwcTbVNIHjLrCYKxAYfkAaiIn7plpCdRYjEjnI416M1fv1ccNe5cMXdRLI8ONB
xvgNPRrsn9zNkcJNscpFWKUlPbmnE46J0enbOt80mxvbo+23cZA7POloEZCAyMPtBquei69LrOYU
2/o3T3YNPevBIDXkeMtIZnlASfOthH17j73VtU7az+qIofHKG28IUKs4tisLgMG8/haTiIo2mRVX
6vVWWrq6hFR0J4ox6ht2APx+A5OYfosak0C1MRaL7L5K4qM496nYKvYOgmQF+ErI1JCdtVZ+YMhD
falbs9AhDtxBspLxAjBHcai8hz00+bPXdYm3PKYcD3BPqOPM2C4jFyfgi/6nWqsuGzMv4i7CkwQa
HahybJWO/ONHnwqB0WXwGsqMi79feh09BwNdwu/YnQ61xX5T7a5Sdgare159jZoXk3cqQO1MFX9Y
rYUx8yeRik3G9dcHA3MoDfbHPT8SqiAX5MW2JtvNKlRDMx9Aov38GgW3OIl6FTYOlMTbogS0WQx3
/cjG/J5rclfrLepUYDO7pZFAn3xevlXuPXE9w6jyFJ+rcbfQOdbyldISZbguZyyoD7qu4aC7MDeM
jQs0GxdF69HspO4umYa7JMoSZMmDoyf3+ODjtKqxfhUOwMWIzMLyqI7794UvL12pT0EnL7p7NcM1
AV6HYCPk+NvfRcDhJsd6vEGxGgmrTnSrwy5VFgvgmytDy90JCJif8RD9uqNqF988rnDqcucz/G/2
qXK4JSYe6x7aMd53f4j8m0psiEtvwPL6CRxKorroYWW1NLqctpfQE4FEpm+6geooBnW3s0VMC5hJ
H/8uLZRBPX7hwH1dSGnhhp3xULJBvJHS2X7uVzGTk1FYKyGKbtpLUmq6HE5HTrYxkAf6bvaQPYE4
52bZKf6GkxijgwHLgvhHm7pPFXsK20KKOkxsJSNPIB99/IxCO0r64spVfSuMWHe5AW8uLvBuNczO
kPoCBUcjZqc3LD/2I5Usuz6TtqV6GwStF0qBDEXeAuWN8uwyahWXF+xEtOzrONPZPbw9cUK/qWEV
gl7v+vU+Vf1LQ2JAXmWmcA5+FyEyknYtKqMBb7MVLPxk9NBv0tzTS92oQ3g30nVDvYK/OxwL2fV5
BzYr9aU5OCsmX4yuOl/3bda4k/mDnD+5sAmZp4umlCzvNg/L5DVpXUfoR6QXiGAsHAtD3iEKGqv9
hH5pcFbUm18uUufMUsrFf3FSMIjPTnnxMtVnHJJoJKdxfALIFQ1yBmRPzUYEDsLFLR3/B5m3DjFh
QgsucMmNJhH44WPZ8z231YkIpRzmvS1QO5VCS618jFCUaSfmgJjFB+NlPQhwNcJiuO49LDHfEsHH
cfVZzjIbBSufyewbC7gusjs8vhoEV+4180p+2lCfBWGxLoiif6mDTUgigNCxtF3qrVpw3rFTksYL
J2HZimP3Vuw4QF8lsRtqljzfk1YaYOs+bF/U+BdYo8sHaX6nnBgiTBLf54SbQpYAK3QaC2saKreL
S2ZbnR8t3PQimedrmGIxZUhyHuTH+5rzwT+nwA0F/UG4gYWCBg8gMq6v+9p4/rCCHXR5SRNetOTU
Xrv+OQicE7fbAe4SnNf/biLmM+D1obaerHAMN7XM2dI3ZodSvh2rCg78WDN6khLr0S/EjhD0F1lS
UxRLe0TfO67I9IAkveurhXx9C7HN5fDelZ11FLgVGrutGtChXlA24pjZZHGHldZ30Auh7THQQzVk
p3bWdCLZ28gHV4XulOWq6dQHoupr9INdaWIk56kj6ult2rvDUWKnZCXp+F0WQkQORcn4p9fRTbWF
lPObsS2YRL4yGCumdCd0tcw1KrPJTKtMXvxfY6tyLeZ2EgeqXK3oTQrzMHVqeVwnC5Qx6AOd2COt
R3/z9pLhzpOxEG3TfUHgiucnM1GK3xtOkxfLR/Ajl0LwvKHfKIgcp3VnUKrV3VomB93EgpGnZUgH
dF79VsY3BtkhnFw1iTDQuwngkBrmhyABn79b/OoY+wjjFKCeP/2Af0ciXw1u47xELJxTgF56lbgX
wUt8anyqzo3+YgUWer8+isqglfzpBpZ6/BCCeoEY/iURsQ8sDJT8c02vxp8T7X2FIdxSpq1CGONT
fxbESliRcZ84lpfDwrNaK0IvC0UMGQZ6SJ1NihrL9XHw2shlFUjkDZSi+hxN4TR9rELnTB+wHYvT
18M66jDJjytZIgszi/LxVavc2fJjbxD91wyhjEm4Mdffo2Qk9sLfko2FzaeCgd1hIAWYqun0ve4q
IQJ1u7WqMhx9EpNRh8nX2wXnPCr1kybrYXYx14vAZwzLJwByFm1YIIihZNNoU8R98xNIpDrbjhH9
Goex35m+O0b6su/r9YYM0SXSNXYsTXlhQg6BdeO6UY4oHUSke0/cZ+V1fpT1mYfS/UqKF/IJbtlo
iMPJVLXIdmvaU+wd2p/jtji5CArAaWIOnI4TbuldTciezVrcYC0EEBKKDIoL1yLyhw05F2nxy4va
cRNQtLOzpwS3znBSJsreb0yVVc7wnk+mULZs0U2PgtglI+NIe1tz1y9KMjJ9++l1KBfn9QhELCL0
SVG4JdIco693qhS+7V8POfgWsUF0O+dnEoZdr1cAF+RoawApeWl/WedHN94j/4R1Q0W7FjbhP1WQ
v1v8v9SKMB1NzYr9cvK53Wr5raEGDLS/6zyLWeU4wqYpCEMxyGPvAho1UJf55vVrX/MOOoYSwW4s
cEWoMJ8PETH/IRAI0R1hIN/D8B86/dFydD/0zu2s2iM3tRZxaN6Yk9fKH2IMzN9scEvfv9OMFze0
1T/Sl4bG8kEMaYOdrPV2/7wP6ysXirUui1BWvSUktdeDkU1W7Ooo0lz8kkyIFaepoBb4nqjDP9+N
e5Mi4Cg8Kb1aIjUN6jOuWauTt8EqITfHwt7Y/UoBehFzEFYO5vFLencZTCfaxsgki7K67quloSDz
0wGZe/cIXRUp2DnIWh+im8gUx1kWwxPVhtVFS+xQ0Y/fhiEB+V5iS0pcX1FvQLtasFdhPpjnUrcV
3MCZ/jRT6Ijymiu1aUTRrQSsDjeW25B88JYnyAnOMFbNGpz9sB/iJVMY0sZWB3xOYGlEodj63g9k
hwTUdSeKGLEl6X6mvOFDcNr+/j/x39/PH0LGmDvbJj2j7Q5vkV4dGc/v3lfL80No8sDFUQpi1pWV
lBixcy5RgFU6+0P6lzFSgUQz13CFwHDZ02bX8VF10IBleXAc/crwFvXh4f5kZO2Q16o25FSe6hjh
FsrSTNUTiO5NAMW43/uUSf/2hKel980nHclHt06gcVBM/qf2W8QvyRYy1aOEBRXZZAsBbp+QeFG0
4nLHdGZsD4zcoterN+v8m2UBn67mm6OofhGtC0TJWmK96d+s0Ockf9ZhWe7LJBA3ZBQ17z5hgTnk
a7y3sEWa9j0w8aa0jXbnTPTiCauSWMGzm6P2WOS0Q4MwHaMdofi9NIF76B1y48zcKkgdIHCexE43
jzSSXYA+lw25gCmS08ar+Ich5cvqsyjvD/fu3ENaMfm0rmdscfO5ST6/gRR6LEm5mPLtinNVfdiE
1VT1t/p4LdWwoCBULBjOOFimO72ikcjxDNE0/0/xDCv+g6BIybRUr10S5g3902LJZimgGecf8bm9
zLJobsow8jrcPZliyyVdAO4p6Q8TQWcf+Dm3DLzxwZKqu5Rjo5f/f2C6YIhb1N542/7/fdGFVyEj
jm0RQcgiPBImLpexGHmfZGKjXXidzPv4dqbLbuc98l5W0BYLm4Ym6TI7OeYhh1pdf8oPIxhZFHV3
xKwtL1qrpAX+lATU6kWBJphiOkC1CGllupbsxAG3It5ZajHpVoJEwwVmdcx5uEyi3mePkosPfHLR
E34gDY3tlO0niVaqTVKSVd8SyvSEXYbW8KnacxyByHlFD0pLgfquQ5jG7ffqqErBgc5Cr9etlHZF
90BFP74rnDA9PM5ZOjVhhSJN4KsdFCVNvxfcv8MW/5q70NO5cPjeo114CUnd6ttfbSp62zVQVpQ0
74xSlTTMPaI/+OMswfJLftGIGEaQHJ+7EO4cOEG+eP+Aq8uK181qW1glDGCET8YGMTdh8rpdb0GU
OzgqA9zk6YHoL+3dmzV62wrpf0j4c/grZNr1UhiivZ4kx+SdVVu0jF87yrueHMk4vN8Ch1ohRXxs
wz0DkAvo845jtTWS3XjByCoIZ6j7DU9z7SLGwLCvp+3tVf6DZwQlrjF83Pi0p+NxpaRsYb1JRBbY
/gyps/PIZZjY7e1n9IiToEYjNrxNQSkM0GWLBzGlWUJOnhlOwcQiYLUEC3TPwUpojXBbGIc0TjQp
d1SLQPyd2+/VQMmfvtJ8pH1QJc3/K0rHkH/SxXF9leDcVjX3tAe9j+x24aebcgk4auS2A/w2Ma9f
jj+5qpOcd6PIk8paGCaAuAtE5rjYgmwV/xeToOG9WDQ2Gc3mev51zrfDNTLAUI1W4AuqwU+PNruV
G850By1iJHpSM3OgMjFa5+SL64xkhZJQWiRbsnAAoVmDaXhjLvOihNlPvVYDXadWMqTN51FK8WR8
cuSiP5kxD78AB21dLYA0x2zDDGqqIUxi83nEP6HFEWWCQ+1gyTStGrAZEIf6AIvJyEnwCbtIJQmn
/NE6p3XHlnsByGxg4MNcUXaEmOQfe7BS1IYbsS/YJyL+b6jMfygXh65uKcIyBz04YTBJtb3mKSTd
1rTfwM5aBLoNTsngT8MXgRhoLckkQCFLZrOq/ZPSRqAjJkYg+eqh3mTzkTGUJorkwpl9XEOMsAaU
7zWbfJ3LOxmuq6wMmiGjR5E9RXz1m+FG4pSa2sGgGd290nCEwS5h4H7qdf+fJeWnPxU07TQg0oqP
b9h5MmGgVrAizIZkdXKh6EyYiqukfpb1atAxlbcKA/fsEVYpV+tQvburBKq+C6rArQyBrr2CuV7q
NP/4pxo9ZrMJtpt4G9G5fQTqjlmnJtGxhRSW3RwH5M0vqiAKJOyuIV3JTTp7JIfpNMLEVnYRhD4V
63c1CKni1nkgF8sfnNotzE9QMxN12ZgvNtqij8zA1jFPZgsRqrbLcTRzWiG5i1b4hZGKGKOZ8GcK
sF7pp7c0M4yMLSp1EvtSDhUfvsDY/HtlAySpxWW8b7sbRecTpxSf8JUYsoChZx6Y38o5AEqLnbTI
6kPeYfoEQ5t4JyVmEAsSb7fUO0pvFpiMNhThgrAcSb3Tq2r52OxCy7LisRhIhVhqCOI+bfs2taat
mY3uJRpUBX2dR33WnkCBMvU/eYVttqBV0QFWtN0qss893r1VTg8qqtlDYgbL0WiJNp3thptadkJQ
oKXOjjgiuhp6NK/WFHIm8DJ+TxoWWGKGA6hCD+OKqCVveLRUXqrUx9GxV/7hC/KObbeaaA8nVwBR
WwCyPR6h6QeBEo1frkIpER6IyIMKDiHbZY/DpNr/hdiIkj/cXc+4VxtgjRf2fkRlhngoEZ+Qazc1
kl5yWNdrtHgXo5lmoDFpDtloTSdbrGVfQY6ZUGruivdw9cIVcDE/+/pL9DRgLqG2Si5JzZnlQX/G
SZWVX5KLVHwoFFuWIirEwOsDidVmN37ozezEC7QKzoyFxYw5ylGy/ogtsv4D5IpdSxgOOQcfr+n7
b06UB6Vg46bVEUV7ogUcutuQBKAMVgaTWfl75dgRBurGDP2fDstIwkuXllX+2IF/SFrfyY9PnrjO
QUqxyx23JycIlyxY4w8bDqF7NrcGPs8YPfDJGIz0GUNRcxravaQ3ID9gtwKLyRJKqolxd0qT/QM1
w6C0BNTSFQjrmQKL8Ex0zkP8lxAFc5E8hAxHJRrps0lNVVzXloHPzoNGmjnzMZmJm5UjNtm+HFtm
6P2g/b9qu0jv+PzjMGRAUCHS551MAl8bHnSCNpNBSwlUW4CJnuyGaQ7k6pTx+HB6KKkVuTjrNdkH
1fdaNVhaBVA+Rnvo7dxHUqcrq0TJZt1v8my2c58PK8Kk1Ylb0eL/BtZvtXGn2RW6AKxSh0RLN2f0
vvIwLh4vYZnHqm6A6EONxDqOArzv6f2QJB70cGx+8eLWBv96CdWvacDsY571tMnVgTtjZC+hLM9S
Fy6stB1uEiB0Z1t43ukaaqAY3P6V22b1v6PgejxrTXnShYXVsQ9NKa54FK8ub0UFuqnTAaK2TJy4
uhQPa+MgLWysHtnjo331yoa2zwWOyZsL/MoQQX00yNP77zE0Jcgl4zJzRxGLgr/luDMSqr2XqcXp
FICONC18dbygNhg1aluUXc6T0w/6vMz1pRQX03LvVvZ+ow/IJlPfV/Qi4vewUQ5oyrS55+MS3PuI
0WvUNiLGcRoiaDdczUpML9bCayNI/nVDKhykLvtd8vzbvcRxqIvngFB+Cx3H8cw1UyV5wQIG0yPc
ZYn3Usfecm7a/cDS/JgOuiGMM+Zp/Gklb9PREva3ndbXTlxfVWJzjcnCKDn0EXPDdO4u4PGwMLGf
N9QLe7FMM0inamTtojRl17VKN+aFbM2V+9hzWKm4rhxik382IzP65qOTEMX9i6ISLe4G9ySLDGZM
Ohfnbb2V86SMNHtE1iAdTiH+AYsTgLRDp9fDTHAACFPih8qf8Y3vmbCrM0M4Sh27t/jdyRjIsZ4+
XNOQUCsN/R2/o9zZCPTc3NHYVL5X4StIMm3GQlhN1xXtctz38Ih0b7ygAG3CWG80QP/Bg6UWCJlh
+yDoR8yus5ngWqDAWuqPM/voMtMiKlETQ0mEqPnYYRM9MJlzndbRm+ri98nllsaef9slA1nNixSQ
HVy40wzgd2s1hp5Vo3sj0PBcDQqBXNb9FoKEXJ8vnArrmmwfnygG6yNdNfjWlfBTJE9oYbZSq8E9
lprVpXLpXh/kcH3K6MPkJUFLzkh9lca/0oAifou+ZyeJLJuqlno78aKaHhiCRar43ENCPAkn77p9
089/56LucA899n7wtkzEaSHdwlsnmqXHZbuane8x/IJrr6+r5GX6UZUZXBhcL+gNevFKcujKihK0
N1m26/wAf2hECoTqi5A9VH+r0VTVRgH9ynQViOSUG2FeSl7+7GGRWu2nNma56IaWXLO7TQmWtXUR
BIK3ukoSG+bId5wbBxb1pe3jRLjxdNrSv044Dp16j7wrWyTc+Ef6Msvqq1qb4SupESkIeDvasECA
Sigdm7e8ISlUSAyZw8Y3Xd33ZzyQiOxPxFVpuu5tLuCl5iSTnN67gz3Om2P+xLTJ5TpE2+QP/WYn
ZIStO6PW1lyxgeUeXEcZxO0Cg/DAjOBXoZwZHZk+fZE6g0Ob0WrgF6v6LWfX9N2GAy7+oiEGP5It
WSepa0YSzu3wAuTmW/mOCT1ESIZPYd7WSMvyvQqZ/Ey25IL+I18lhAe48Cw7Fsx3Musi2nHk1QGn
uOdrBWsbfWD507ERyas5bml+2TwpdEKT2p2tPcVD56o8K/0BZlnWvYN2ADTINoRYa2wQqa37yKQV
5NcXBMvdfG0QP9iMFGPbxayVO/zo4QTfpM+rigivrYAY/vgrz2VZdW49EhZNdOhi48KMlCAUYix3
xvcFaziRQSPBpz2wU7HUDgTileo81zcEaWwIucWorwOgOte9peADJZTKH5bVgFdtglaLStNF9QRX
+FtBKDOSlHciuvEtAkFAvPBHBci9nEV71glL07/3szjW7Qzrw4aRVtwjDuSChZAi/keJBczXrDO7
jvtZWb4PIiWj7n+zlAztdG4OPC9P9yZqlE6RwCe06lJfazEHZSKgZBl3ZGHVTnIa9u/iWpElv7nx
ppANDnX0jytwUVkfiNEE6jLY3u5mULLFip9Mi3EOigvkCiIrhBReEHzldfx9/1MDzSn9Iis2Lo4D
A51uoNmENvT+3OzsF4ryo/8ql6m4cJKbaeAca80vJrwIUrDtSlrC8n/GI/Ng16Jk89gSwJi3b2tH
0Vup95JybfBWAH/ZffaqFIj8SBK4XI0qQ1bF6bR2qrmG9xe/9k+G1KIutufpOf4OS4STV+XiMKQ/
Z4TBoMsSQGLVcGyj9xMoyhfh4wniejaLMeeqxRwi9QrX4H8kTBFVufwITyOjykxh/D8NL5YXYtWO
r1aAq8wYeP+B7NbCqfjPBpsBRm2fASKSDIq/1odB86sLRF7hlCQkE0DnIImuL6qretxtwHdYu+mt
m1H4ulmA59Ynf3WXI9w5M8LQN1zEcf6ponouXsefSoxxE26BRKSkoafu2KKbtFVfvsSr0zLeYiDk
FGRLbtR75Rca0bTtfooStUgNOL8381cxSqeFyjA0Az2Qs9r7d70Q+yEP5cArJdZKE51QRiAkMDQw
lltX5XeZZd7ToZWnK0UGIg+NCjep8Vochv41ONuH4q4KlE/Zt2uc70ednJNmoxaIidfXXnhr5HsF
Z8NkN/H4TSnJmBGl7KMSxce0iNWIa6cV7FgDyu4sueU9IzZzYZ0GNQoOd/TzBsWKGZLcSmFfaOfX
bPTV/9AmU8dV+ge5ttzbjHzTh1OnlenG5x8Cy+4FoNnXA36TgIHHR/dFiOB1UxHLVc4oAbOY/ezo
04KZv1P+1L4wnH8Fism0mZLTDFDvpIOB0hIh+kY8p5lE7M7d8EEVwZ0nW98ohKsQt47skI5gi1U1
Q1onfN3Fltb5PEnQALlqFkeJfDKY7dn+WdO0oYBF2F7ZJhuxM2odnoPsuHDyD9SWRu82PvApfvXs
WiQvUvQ1w6MSUNXhDExoeCB/xeupHRKmd/lodzpKq4jNcXm+GYkwDOkmAGiDSqJjnbl2yFuVTDEj
nIGJlGKg9VHbKqhneCzaXdvdObHw9tb0EUnQfz0e38MDpxfZpUpzsn1ydYc3fHPde1+JScXgFlUZ
XVFwNVaLRgEjYvxpsecUWVie7/7cNkNrvvd/xerWi9Urg1UPAkOLPkFGQcmgvatXLoszsqZxMSGP
SGF90FE1eudmOcK58lr4pmdEuWVGg++Bg2Fas82N3hqio6Kg+l7/eliIAWwit0Gf08hAURsrhe0P
xBpWRT6E8ma+sl0Cqt6+eccZKRNpZj4rkoOZs8rLnahbRaH40fmF5+9Uhlt0He7xKjI5aXbTBqm4
+umpVAWJxCuYJS+K+wxfoK1UetbhjB3W2wdaVGbXsAYT923k5yD58wxbeF+ZedXkTQ1hXFCGDIUn
cEodeW0EwGkJ1fx8efjBvIYasPA2QepX5q1VOlNVXGnsEMYZ/n3jrdN0CZ8dtW3EfHbmM5mJv7X6
cRHlAkcOge/tYgR8RNGQOR4D6t+OdCeDYEwOy9t2xD/4rDc6kWFxnXJp8q50FmRmPtIUcKLA2c2t
dm0zXahtIuF4QPCNxoDVuvKWrPC8Eslh4dQgXeTjSXb48hnwDDSfqWh4S3HsAHkg5ZwMQv6p5vx9
LKJqtYGPiGCDKySs+fGgZ2uINaWvvPRXPwxXzJNSKjuOuri5g0OfxuHlUTzr8D6+U6sM+sIFXVAh
yNUip59X0cY+JiaADsOVJnDDwX/hNMiYPpAm9e/OQ7KuG3qWxYajiJx/e//Q9WMUIwLRxsuJO1Cz
pAQMlefLbHX3eSHpj6hkPk2BzhX5UwErLYdTjZ/z0CoGzcShBmByDcxLZajD8MHlLn72sj1GSAyn
5n0BgVquaXSm4mHP1QESMhPR9oO/aVuI+bQ6vTutJxH/HxflyTryrxaKyrJzrqSO1JHC+eCTI48i
BPAsXeAp2/FPEVzPm7LyJpX49baHsKgie565MNzZADMNOOdDCHq+bfdl/tm0LRjVqp+haU3Ctjcl
L8GBBm4OR0HnUWB2AbQ3HgC3kTNk3eRf7uGWTZOj0j49B6WgII7GHji0NgMq7OpXiJ5t3sfGL/5X
9yCKMB7xtQ9cj7Kd7HMPNZWQ6RIoeN8Bp1TTJNZ6oWq4Z7phMjo2DlNTnu2pSuIie2pmqWAb+jpR
D+k9uS5oVtzNzWy+9rAZLTKDQ03+Yu/OJkq6kjt1hQwQ3/xj+YqVmQNfx7vzM9ind9ILZP1h+/IU
ct1S3S9zgHZHjSxu8njcmkn7am7jJOBtfvP0pOu/IYEBP0oNLxGTdQs8VKczL8MLxz8MG4+x3HnV
dtDQY4FmwY8I9JPhohi2TzgI3lljS/9CCe5TFH2nPzUXpR0IfGEoURv1CjXrNZr8aTQUr/8kS4fs
WOTZRHatTXQl+BJ9SIu3SwgkW1tafGtKUg42rxKeQ2G1DoJZCHdEaWiLtHlQ45pK7KMAymEzN7pl
Ym+x9JvTASO+FVnxhIQMBQltl/ghTfSumusZKHBUKlIriyI3BSRlDT7O3LVO44OZkUDI8C++gaib
3cNvUeqMzosxn3ENo/7z9d+HvIGS8yyHF8WXoqejszynxdwCbxbzM5vT+I5VRHYCNh7C8zNWV4a2
4wc+QJftWxa0yxMa8BMgImklb2Kb9h+EfmJALK3dNsPsWXsnvIyez1jDVWApGQn2x3E9RDBEnGLP
epiDclj6hx0JZ53PSxvhCd/peEgJuI8kFSBho2FbWJXZcYqPHnzUqZHaCieVjiLuqsvpnLT6auJQ
y5uiKrCnw5JaW6fnTj7z7WQBR9MLg6krJrqvVJST/xRA/XUsRL/+OH8PU/hRts4aLoqVGlJQH2nn
Q46AuovbJtx/qCQsDJv9Ot1FlzjO35KXnZW4z4qMs5XWqZ0yGozI81UabAk/c+WZ0wCyzGytqqq1
CrGhwmMbDWsM1YQCvL4Buv+UL+EhJun9xdAoQ4rwaAqyugrSzLJCnDRVjsGhb3i12GUC1G2TjDKU
aljjIBvwQ7ZuBIKxHs3VSe7bvWIt9IoRTpAx34QX99kgKo9Eabovi4+qw4FHeQvO8DKE7U9/XLsx
mmeWdRA6Y0y0THMAoe0lwuaj0lhtOUPOTQ9DrvEW9h+O3mUC8v8QGfR+44YxeEhJ37TvLTNofpq3
OlLGvSE3PEhO7/mQHgAqA3NTkznb70ECDxL9Qz78bZ29cDBl8oX2uSjpiJpEhbdsymgSo+G9xbCf
AXdGHLdJHBbtt/pWGf7wnZ17DRcJgqznVTZvrz1kml0AwZEDAs3dbnzlUM2g2ppO6+SvDkuqeDvF
aeRrg1ff8CNP4xAjOeggEff9KVqQZ4tYtC+u7OOs5qTwEs4oxtHYXSY1ePzxP0pB8hO90/G3xJ8+
DeEyFdbQ+KFcwlOMwMROx67vCbq59PXVYUxm2I/uTeeGO6v4o8Ef+Zwiw+iADmHa3suaXlm3e4ez
nhLUYU1RJ/51Flu22eJqlqKt477702T66CJ/M/vNr2fp10OnEZRBV378VXSC7i280Jt3uJbKOTRj
NA+Dw3zuhnBs3T597gxqXryXxw8jICujjk79tydQwsR7A/5M6lKeNdiu+uzGyoPS8OvKUf4dPgzA
IXYDGAyZwjpAMxSWzLh1uK8tWVgtc5s3epWhpKUE0Q4mn4Uj6FDVCJOMWwtrHpjblk7EV4o5YoXD
T74giBfssSLN8AjSWR16SfI4b1kf54uTvzfNLRArKwgQBl+y0q8/Z2HiQkTbEypn8hxN3xDCsFBB
5HJGw4P9OpubtwoEus7l6XKcZfvgohH8oCIr7ocyuKjt/9rT3o2GJearqnXD5VUuQmY3DNUEkU6F
Xe23knVGflgwIYLCe4cPqEktojpCxXYvCHaZeqvZk2X+KRh4YiTJ4s56WVKQEj3EnozRkCTLz/Am
JMivVuJeDse03lQiK740Te+nMz3jH3sr86F/KLe6x6qzZspuOjq4OKUqKBh5ItU68qayw3DmdhEl
z0p+Pn92YkyttJss855Qe3mbhsk1tu+ZTObCJr+7ZASeOMFkbJsDjBC1kA0fLsSg5ew+D7bKaROY
LcNqwm1CW7StCvLwL11HfpH83oMDOEZUJEIlTwyGy42ivhIq0K1bMjPoy8OgtUTsNi3jMsX8TPKw
7HEjWOvg44dqhp318DRCzPZY9QMW7m6u9jCj+d2gnnlOe3RZwsxC8DlxNoaJloTVDhuc1E4QeKp7
iO9NOielO4xa5/XUFO7YgRwmkP5Z3fdNawg5jLNBhjMqcjqgJWmmcodsI+fUh6LcqRqRtivOk9gg
12e6WCP4jprXtSjGboBOa62RAHeJeebQ5yKiX+kWTV0iDCGUzFJ8OiFTxFXa3VHeefYnrDC7ueux
AF0YEgLHqG5dM5iXXx4i0giEDr8k7dF3q+fQSuIujiJol+rO3x6kJyZGgBYtleZyBHwBnZY0GKbE
QKrRHsngshRAAyYN+eXBvs/Uv7rxt4GoUHwkSfcXqjtgSncrvhEYlzvwrTvQNsBYWaMOyaBTwpM1
5BMyCWP/Jkb8LdYWBTbZQN86fKr09MvbcRJ6bfRYnI76/P24X7LSjX7baoVam5s3U6fhn1FHEcIP
QUZN3BFd4SjgIbUGWrH0gc4QE2VqWcxJeagy5Vp+RZcalUCKxj0NDtPnCOEel2n+LWC8nvCxSTKB
3Pnc/q84cMHJWIaGF+OXdyujY5X7/DZ9lG6CYbL6dtUxIXjjbPf/i0BC98T5OzzNs0Fn535t/P9I
FNC6bKG/2dZQswHqDd0+iXnZkHPmsng4sUcFDunn5uUzel8RFUpUSW+7bptIhPVPWnbml7jQ1XVL
vRjPQYPpuOKabvhfUr3gjENNhd/aOV081A2dbZ9Ip+pJzXK3Etj8XN03DJehUKsK5APH32GVif5O
EqxO/qZINxPdMKDS6HzPA2Loo8wnYfZ3HTLblI2EUfYpY3YCjmuZnlCD0pwPzV61076kVwkdYlqR
wEM6Yfq/hsbA8s7mL7eQvAcBo33DlC6jD/KEewnC7T7YZWyElCdEoQE4aFaDj7ZLgMZ+PKLuiAeJ
hxoILHF0MfJ/ldv96GYrF9jjctmgfXiTYQgkqZRDd7F9NlmvenoTEpBGUBEx7g68inPjwi1wDzRm
/PqlRMqFJw2H/RTeKG7r02xzzoCm3XgrbTC8cnbpLIbXycRoskwgW5cLRAPSTMQ/JVx5+93xyiIZ
334LKYXk5pjMYfzfwxRBnk7FRcOrmtS3wbPayDdcrHzubN1xTiC9lu4H+Kz2XM5OGMBacHZL89mQ
oUJ2q49iUXIINtTVMPU9hXlFg3ImAkWc5a1Jc6LTPnW2Hycw6NLli2E+9iO+aOsiRudnzvdiGh5w
ZhxaXqpSxp2aKx2Ut5CXMdk+NjZ/ANdkYf9//0KPulcueFrwpyvdwCjW++j3QW2pbAp9hI9MNKMg
Zyu/JHfWbIHIZQGnnW90PAqAO2uytICLt0JP0hvEopm60/PwYL6d6x7FwFwDbdjtsNv3w6bjsxWJ
DxkDhNsXnLTWxtt+g9DO84xQ9IIM0NXCmPPYPvyf5NTItlflXNCmxehShKPO+nuAnBv8UOtRyR27
w5xz1nuPYeWBAKpAizxbsrKgJeVHg02I4ojcyFDSGS/OwzeX+Y8vhCr+rwAMCgPkaif12L0gwxP6
Yx+PCetvfSGXN8M9k6gkDWArCuc6IsOMbKHEt97R+aYXjbDxrCU9wfWZSAJe/J6ftDp1El3qH4RG
eco7AGEXr2bqrtXK2+XwztU4Subh+4118r8xvtw3Vn188FF6Yx4IpfEplQWC0vuMdsj4oP1SUrLL
tVOUzq/dkveYSTuQ/veZ8GtLb3Otws6JUg+qMemCy1Uv+N3zfT8sIa4fAGW471oZ9bcfFVWler1f
HXfc5PUVQ9wWmqf6uv/VLk5Vmtynae4KXf8GAQ0L7dNHk3V7tcqhUkO1oOS5PTGcXIl/MDDEDRcz
efaepbJJlmQkJXiUt0JkiIHu63Rwm0voV+fVXbiLbR3Sgsg8pWh2GXxjftDFtvzkhocm9kHSUSOy
/kPfyHVkHYxbTxxryy145sr4G3x+siXA0EVZ8eVLN0ux6POe/ppkr/akWa4MOBKobRCClFSY73t3
kDkeJnIj4cUx9zTpUyqV8zD/3tlijtvPfQvYswkljpZz2MzeNwhyyiJmaX2kKdDqvQshBBK0tmiD
zbPgH1TDoSk9p4Yv7EfjDkf2rfTaYm+v/44K736zYP9UocafnABAj0fRaqIL71xKojG8bPFdUd8v
pvMz5Dg44XzJ5WKQtz8VjIaikbNjuDB++1FdJBBm6yt/zG7TJ2jdSGdugCjfz9WWlrMaRCYpNi/g
+sbpCFZvpSBjXz3tw1YUgWRBLsZqnNxglAoA5P36bCoNOco722DM5TOOdq23Lrq7LzjAabtgAp2y
2dTF+aqUfWkF/aXYcZGVcNkmTeoq4jyLQ2OmHx0+knp1VyEzhI7VcPX0rlU4AK1U82XL/mDl1k8/
lpep+WXCM4Oof1RG3G7z65uVkM4nJAVv1fi3hc2CPNkbXLuMDTbnplZ2NOlQ6nlTxqiDcH+c/+16
Jbo8S5rsHi8rXDqPVQCtKJ/hbETa8UXej95dOy5Q3VxAmTXxdcNQjkct3nvcmjJcpFqzQW4JlBC6
im7wSFh4FzvEV0LiIgNojNIj/5SdHlgBNwKa0zCCn2cZdV+w80wL6PdRuop1xkdCsrD983COIJMp
bVBSb8FcXlex6kBEI9cewL8FB5QwsRcnLu3z3AWAEiB6TQArl/Vp/g1luGon2PyZJhsojbjUkyrx
0ird28187YTt5yBw39G+q/fxbEA30LsqXmPS0YT47UoBlm4Y/3m27MyCzCGPH8shnZCGbjWr7Xsp
bt8YME50r+Qr5U9YtkG04eaLPgKf/VIoiUcMBrdfyrVVz+mJA1N55aq0S4I+nncUrjeVkrWSzF4W
qMqDUq25qdPgkayxIJHipIvZddfhaqfDx3pnhpdqj2Ty+L94C/IfsSTegtHr+fPgC94ndzgCxCbh
dcBZukjfSZhSwr788RR7w7K8ZRx5f6dWyHfGCuwn1SaYGYvmaXmKg03HHS3ydZEAwSf19TErIGLu
NgYObYGcdVQpJmYROjo/DOermkYwkUcT6OTNCkpXq8yv4uFXSz/7yIAew1Mkk0b0MlzpoUNO58kI
10qqmfqkH2WDNAVUxTakiYeBGS+dMc5vbJKup8e90XiHF7l2pr1JmLtLmhBL5m0Ai+kouDKK1CPd
mnkVFAO6A+oqZvjy3fqtd2lqt4fvpvnMkO8wnWQwL//QuqdTtQmQT4n3LSQOTSYlYzl4/3r9PBUK
Wp5xzwwCeCtwmrTuD6k0Ju+BL345Eh33FrF7ORie9aLMrIGOFpnfDcTPsgup91YkfgG8G2S/dEPk
3VzNfgAm3uj76rSvG9pR35JCVE7HrKBELFDn2CTBKsqzuNusyYwEpPO2aWkGo4UsU/bHu6ZoY5vd
iiW2Bk3ZQlCSlTcUEvCGXk3I9RhjUu+SZOwTcpxGBWJhNBciCOe3SB+Kmm7Z9z5ROsWwwogkVMIu
LgLBD1HuG/sACSemKhXF7W0S4qq+7r/uymf110SmGNYLcxdP2fWerllEHnGdT2bKOozrmuwCP0tH
44etuDlN0BL2FMELUAv9I5V6VtOEvcjczjszJDMrTL0+YKzz1AqzBaI0nMcjDnH3IHB6lQBS+FzA
hrNYXNvSrc5vb9wVSH4O82EG7Y1OhAIfvphphgPUEohGJBCGOJPX0pr7FeTCzBlk2RX13eWzm7dH
uAkHs7V+q5PnMqesUuxvJ4dA30ktyeu51n4F1Q3lEmPBZXMiOK3/H/znsk3vBxV3sKvUMT/++ZNY
QJHqOSLUyUS7IgR/sTXBGGDHzU6F5VE0vIsxzYyHbv1xM6/ToMX9sDwE81E8t1SVAIDDQ8wwTh6T
8idnIxhqxvVeWtzDiBWgs2hSdcDQaGZIYAvkMraChPXhJ2Vpjm2vqddeNtVUylODPZ9B/anB6GRs
OGd1KUheLuVYTMBh92qvAkYAEO0ox09APuoOCVUDLAsL9iKhgle01yleAPOuzmSQnqHHc2CTPnsr
ThsPd6H5YcKF8m+w4dZhavjUdvWjLEW1yeG+HPuWp9T0+T/feDBJxcNeRWal32UC+QeLvvFUXDIE
RV9zI7zCPXwblseFSR/9ojRWz/r8NyLYYpIeqWRG3x2jC3kfe58rOgyEMrgfUZbkFSp5jm5YBbTz
ho98DhSlRzaVWlCzE6lBGwc80mOOFK53HWQRgbR3+xMMKEfZClwY/zLYURFiruDPhe/FwOEXGcBb
0rs25EKBHyU1loNP5LZmSuGPB8i2n47T8CPzzOxkNiEps0eFCN+XuRBELzt29ocpp+ss/tvLmDF6
UCr0tnGcG8S6vqjOL71iOMaUA20sr9vUTX6Sbtz7fRtlL6LFNKHQ1l+RQFPgR8YgNQJgLNXyfphq
dMxE3yLOAzw/LQMS+QGs1vhDABBvCBAsSZ0AdsEOZBJ3Pn8he3wsn8V/uXn5mHvPVoavqdBeXY2H
YfOEuPzKBVbGpznAoeCL2zJNTgncNwB6d98AxsLHHUixJXxa/geLyWsvWqNjgyRJ6k2gjrIHdVkn
nI8LVi/NI8xxvjmYMijybC3UAo/0zMeuENy6lbXLKc1Jif8VGdOpseYOVRPK00/+mzcjJ2HZ7fuq
vBt2RjPVf8je1KOsqWIEeseqBOGa7NcsE5rKffHgG+YRKa8v17BcKc4JtfDCGnCPvZTw3mltJmwT
phSMST8STGVvi3lvR5kU/fwOEAGMHyGw4NnqK4blQivcL74gumBTR8GQc2CT0nJB+9UXzKcSmz4d
S4cGVigVADXGoVMB2LD3uh0I0Eo5ll84R71OhjDC9sw3Yk2v9tEmGBZApw98x4ayoCZzdw8Xr7O+
Jj3X1rUJu7Yu4I7WyJz/RPAPtifFnTzblo0pq3tHzRDDTpdimm9dbbd7wwovzGzsrDa8So1ha6Dj
mVZKhGcFyXdg7nwzh1vNaQ90AnDn+Vn+1tVhr+JxwqUm8WpHN/3Lgax0/jA1E5exD1fizAV/SOE6
ajb1h62TqrlK3lVD19mECHAWHcZngwVNbASwav3wC/MUOU0q9i/Nqd/iH9xxJNbSstVeBR3lQD2O
GtP5TOgB9Hs7C2ymp1FGCi/q6g6abRaeyKWJm6szxTZkqopPK/w4qRu80y0H7fhLU5xV1GNrupRh
iK5qB9ewwLlc4BHsqhdYKGAS0smwRz6PO6WGpnZoX2KcDUEfUh64CJGw9CttL3bAZ768i6ok1IyD
NYLtdzF0HTnGHu0TY4kkfOEB9ks8fPVLya1ZZCEDGCrcW0Ov5I/rPF08kKgxYmyfPwGMdjCWEKTC
nJKGBA9vIg3OwLi6oSKfS3qyWn2VAi/8uu6kWlPTblBLOJV3knvaljFEKVA3pId0Mc1XI50oWle1
aHw8WWsI5iLqKd1hZaDjY+Bioie6XH3x1OTyVKZee+IRejMvo9+DynFiTJ0a19r556+80PUIsC/m
9sHC2nWggcO/6rUG1XJ2oK6w26QiQZkjfywnU/HXxmezt6kKkNUvz1bE3jFA+fARzysmNUD0E5hd
2q9Z++VlmSGmo+VRFQI1yZ+sPGFDwW3NudjassDx6s4MukMDa+6mlnMBcqWzgRPr5p/2Gvp8VHFl
VznW+qnTA0H9qlckB0PoWawfnaqwTqWYiOGdRhoEw+XtLOfclBP/nnFMM1Sc7MqOG/Dx1peJrsdw
k5WU5eLTVfr4lLQDAuFUMfZOrpaHCaZ5Ddk9VbiSNl0jiW7iW20Rxqo5FFoizgKBDzKOAC9JNwYb
ZIPg6KqB0xOCIvPuTTl0h1oM/LR+7NPPKuk+lIbY9n+BjmPKE2F+1G38G+VYxo9nprPTx7CoEIUS
V6+nq1JnOriJ8i88tbXge3eHNgERuvlg8f7FUqObwG3hC8ZwCyVgQrCy4EyHOhcHaMhWmnP/v+aX
wkGIuz1YrQQs8RGIOImtri5FoKHbQRqQ+JtBlwC7TaD9Aaq2AOpEpfuYQCgadJxxPe1QKgwfRJfP
cFhQx7buXho6v/yfCXbHVtVUXNrSlSnMIa9HZynv+28VQ4sKJODK47pb2XdUv6cm/PwD38VHpXGv
4yb6I5ZLOBDQID2ZsL1VVTbv/jqb/UtU/Vubh4UziiW72l00sDNvhs4leVLZocsJfqnbThlaiRwo
zc5p7tUPKHW0xESs6bwOkzcw5ppMKg44/ABrxeSVmJhesLejhGJb7Y6VXYepXwmzk61CqQAa71cq
SVerKRVXBXGuNHZnBnZBchj/xQfZ2pRV7fc6JKvoI2eIDAPD5lrWJeh6yXBJQlV2qxN6rpN/7obj
OD76evJ3TVAVd9JcLGwIGA6Jpa3iNX+ao+fWpbxDAgvqbpeKhsjJtRyR20A48iJ3Mvrnk3f2QxyZ
GS1uPgil1lXfYIGCbDXFqCTO7B7Nfllncv3j/Gvk8rNEWUTWCTyf1M3zO0uYdHiwg1VPvJMP48gH
nAtrB1k7QhYgUizAmXJ+RAfKEJXIRZjfSGwcarX90yrvg3y8ivZ8wltr46fzkVWpj+ZjC71iLO+t
Fl9bFG4auLHVd28WJSb8wJVbYQJe+bInwr/TEEca9YtBY0rLKuHMP1gDQrVvhqho4ADxFJ/Yo2AU
shZLv5Cp7xNgf4AZpimQC7thmd7+kgzgYFmWS8TQ2bcHDhVk8+bwzwafvG9vcGXwXjJDFhbM4YhR
fYt2xTzmDWNcXqyJ7GLT6klHZd4igj+rGkrX+WY0U1U3Dkv0z3XteghDHgT1GDcITBOAMEyJGIpD
uTowblkiefP2AidgTFqcvQLDGHZxBbvN1azp08+HViCaiFIJIpP07/SigZsbNSkjBgNHJynBXV9o
jPPWlHn0Mq7r4FhNMXE5RGQQs1n2ZCJTDD1PnJmuleQbSLFpFAOexADBqkrjLw5FlqReECg150CZ
wAbBoGZwtk/DeLWYlJDO+bp1ax27h3CmY+68Z0QQi+fnvwGSGcBfRhtDYZ0FDW8aN70vflCaK13F
9N8pMKldsKU8coVY8m9x4m7SQl4vJqwOj0RMOF2Cm1MRwP9QczM4uXGqdOHf8zhpT4qup+Wkm3Vn
or46pHE8z5mrAGlA49sHe8jCc7WtQStfGUooH2IFPS8CNIbAssZu0sUbjNVjy6RbxsVGkAHu0s1Y
L7o6SvPm3MCfAYs8RSRrq8hyAv6i/49r+DzEKO4JwkMNxdtbytzyzfqtYmbtDrla+7UFqgEP06xa
qFTgegWcvMARjk5CqVnHWK5LSg0pmKnTleD7kpw0CS8/ZZxRuCPZwXz8/zUtx951G4PBNrXJNWNi
ow948HOeEZ+5LtL2KI2d5vgkrradZPtp9n6WyEy6bv2dCJjp0dQ9x4PuFiVbPFBdC8X2U4sL62kp
W06z6sMTN196liL4reXlY2oRIU31i+s5gKt45MRuqDDXfd94m+jRfJNz5+8izTG09coiZvEFxXxM
VKkFRWJE+2grl12flgs+MqbTJ2WU/FasOwlGfOND6bqaL978ddaJ8fTgotWKLK+50J5Sd8Irep1Y
ka2sRNoBdRN2Jx4RHw4oWKffrEJHxGOKFoX+oe5t9K9DwtfH74x8VaDXfxxSCr5yihgTAriMr6j0
FpbanO1reoXwsJFWrzBqhvSxIxOrJScVyxG2KXLb0iBMr7HL7u/fN2Iqv1ELewE2RP7uukk4FhQd
FolKoBCYiidMjo5b1esLI+OYiYX4wuvu4onAKImqhrVlDEXUAC0Ke3ZPfY8fhnDcWOwvzGIYHA4c
OUxbPakjncUEInNltowSzhBIIYKZtDOHhDv5mZ+zGCUuSiSjOYfkGauN45pKMCrIyQ0aRi5IYit9
UOp6hsmN7/56AQMBPf1X9dC2j6z1DEUQUSvcL7fqC5l7xTiv/V+ljKREKz2Os1rUmRzkT10By0BA
smdM4K76QeN+C9NL7JFuquNt2H1gSdsHJA405m3yRk5rAYmD0Yme6ihY388cGsXJt7jaWjiRajGu
rDJiEsNQZIjz9ErhzS8GRbYmYB9/0ZptNmpmXaDkb6DYSLRr1/05O4hbXetQyDJ3Bjbcue8p+jhe
2nqMYM7a2H2oiB91VrUEx6Mv1eRa6vSta0uoAqwdyY3CMqEhr75D+qVev3ZlYodRiTYyQN/R88r8
qdDT5l/6+CSgE5tiNYZZtQfYOFpzZdIRXQ7OWzOUxSoMNHNYMwdzUmcDJSFztFkMz8FdMEyBkD9L
GNeMA6fG56kMK5xwXWx6Odp6Cq8t3gaLs3XRzBRrxD4rhBm7BcjMbQ31jUfc8k8TQEnIxwRzqWpH
RYMvExQsUQ6su4DzVBIJkUppk/1WpiYOXyQRil+tcN0FK5p/ut9xfaYPL85oFlwVEy0DqE5PEF7d
a8mmDb8QmCZXZtPAClB8hhyOEtRCu0sJZ/nPzYQuAEfC7iP4yaMtinZpyPWBomI8DHlERAEO/A0Y
7j1z6Q3R1jXsG7roiYGsiDrW54+y7bsOepnUrnW294fO6jhxBcjaMEDTV8N+ywXuPSbf/OMF2xHs
OopI5unJ59ZLDH0wR2IjTjvz8OoNfHs+vbCVGixBk9OWh7Jiv/gkiF16B9144CFD1Y4BRT+zXpCT
igQj0dv6eZYfPw1ZNJHn1hNxsjcPQhNsXYCrob8z6haY6iJH2XlpElNtldvfQNw6QWy5XXyQBsBO
vDGAPHqoWOaZ4klbMt3rZjwM6vFeoCBHk5fxiWmK3MJAHoo9qRJGLnQqbKkfwRWoHy5W3xCP/IUt
pO7dn/2mige3hAhixpCaztVoaPoKWmnsgxMWsUBc67wXSH9K2qAzLd5MOhLcCJ88m9I3erFdb/OC
zu16TboK9o10ft8M5CXaKLdKgHXAtyi79x8Mw9jWBKokAKoo2d88uvXzcvMBYHH0xNMtMaGjOowW
+1IZTAr02F0ZTaBOoaFW3V9Q+4X99yRnLCb20psLL9bGr/Wy7td/pmZlT+/6dMLo3ynl9Ita7opw
U+iCJLzqZ6BuOQfJGvhaC8jBR402GZyL8g4iX6KnVr2+xh9WG3kEoRsgV4d1wueZ8oJpq27HhOzt
QGoRPWD6e9aCsrSIjQ8D1+Kz0251whfs6DdSlKJGjjqxko+RRpnpeKEhZLxySzCYnokQTE2abz+T
NdDvhv1ZlNnZZGeoG7UMR1x22iJrvBUJIaCJF4OJqi5SXimVRZev69aZXgKBjdyLCpAASC7h0Tj6
6JlCfs1VGx5pUU0ToJl0Ck7QirzcdktXEhHY8RUYGZmpOqdmYiGcazX14/Xhn6RWOpp0puNCoiqg
/C372wX4hWhFcZRGJCeuIX02BzOcXE7nrElob3+GlBgYsn4qcNIc9TaQfIG4ISkPcDB6m8r0KCN2
OHhS0LfgTwp1mXB2sjeJHpnGdLhf4XeRPXGlX+r2VsK/uLdpo8hCpI+A8fql6wW0KqICk4NogPfl
2SJnekf+EJt7Eql4jVvaJNofGASWel6odXs52Op4kestspqfABsecgN0yv5n+CIlJPFSwGC65f5X
uIK7bdomP0eMqzWy3i3GStVXm/17aqNwwMLvRV2THW3d4RRxdRD52RS5Dd7ljWLfII2sI94H3uL9
jCPiKSj0dzmVLQFxmCY35qyzZAGgmPvQgoUe09zPG4AaTDBXzQyjAGeWvnw4l5jj1oXqa7PkosxS
yz4OSe9ToE1ZjRuFX/Y/Gh/1L4+WRcZ/4giGmWZ7BVag1hQRSM1kspIest+1ujRBtOfJJE/tfdYu
42NwpG7m1vG5EFuHd1NE4zzM/O/ggkMflwQrzimURRxXV5yTvD2ZrjyRIZa06cVPIN93uP7F8ycl
ZvMMhHoZTKxcpI6MOz1Y1l2r0weHTxH2DkHf4DMafC6Bg1eaUgi8wI25n62hFsvX2x6339tFliqt
hJO+jKKWyaI4zydMKAKhOOvX0zSibvRVIxfW3mL2JmRAK6MGoxWOP3bTofliSFDYlE9owTsIlq8E
IeWCAwMYz0fGtRMgv1OMCZdeDVwYkhceOb/Cz79elc8+gRjIj/xAJp2fRMYKZNx9bBexLtTxjktl
L/EfO39KB15Od4WFDTaqx3Bvbkzr8/b1/bT/X2h/DYfjOLo5WuPADtD4kVsu0+8CVYXA/7zSnuPL
x/e9Vz6c+nm+9QrHrCHuc3/HyL0bE8YWZAG4d1E3NF6X1GXoxGNSt3YI6MmMaLKo7qiVfy+N1nD7
smQuTh5KK/WZGofQCkc2SJ0ivh0AirNMyi9opPefj2t5CHrbqhlFntaCMaNashVEkaDPrJh40ZAr
wHP1cUKjVvlanv36dngFzOs/XHzX28cHuNKvHNfTrAHSt0RdCEw67xufK+MoOkVOYJrKMYGXng7X
dsiY9lyjLK2ruBP7bNcjFuRh7jVgAHN4NI13TDsvAh3PdX8Q4SzmSHnNcztf5h2rKFY7b6SF6zGM
teWanj/h2yOF4nv9Lz+oaujC3jmBf1g5WtiDCKVWX+Rd2QA/YXReSRlvoNbEZGk0cWsT0BEidlCl
W4cwM1xl4NdihbDLwi4BZKXQcWjI8I72CCk0BnEpYJ7BXhKtwddfBrxav6nOq51+sQEVuPM/Fubf
CxHBtfo3bLgmprBwDh63A8pk+rtMe4SOdxvtHyKI/ENvlNBm9IfAO7XRg++2ALsDl4XwIRk3ccbp
QZoINxNggkBCC99fSRux406g/p1ZkpQZ49h2az4lsLbyqKTu2M7rxLRZIbwMXyqxIbJtwWmn2A0f
gN/6+erTeERq27LPimhcO1IjKuhIunCuEmMEOgEM/i9HmA4YVqDYmN7B/dCEWD07oB+nnQxOkIGX
Kld7D41kt0JZ7fGzblAvnIg7cyvM/6rha6ZIv/e3R1VuXlBHBGqcpQ3em4bXnFHnGxl52hdoaGQg
vCC9ntLIlPZ6tXxEkCE6lmzEMXV7XBoRL1feumu8CYfktGlFbGWgE/3IihoPmSP8xwbZzzbmQEJO
xVnVHX8UF/OWvXibtRV9sSCrdOmSBvbl3VIZHLwju5BHQXh6/K2CSyqt9hZi+EDZaKO51KuH2JNB
ubvU5pAUXKqqiMi2O50n99xjeD8jkdw0cuXIYxWXoknZehYP33ESqQ5YbOVmYr+M65NaPs5sAgjU
3Lqs+ykfy/cKxWvunelQbWcxvIfVJwKVn3lFOtbjUCm2chmkFN4fNtLLlNCJAWxEMrq6FzHxNaS0
MN7MZmagBXwxVHXwtx2Cmrpoe18fmZDwOzqNvcPnTXvACcBN5GnZtYmm9GzZGVm+ZYQVBJ5JQyF/
5/FvshsdXvHG6Wx6hh6sAzTDp/NC+xxLqF7rZEoMSPHWAKU8T96VB8QLdAdQd8VRPFgTwcI4nCkw
f70i8YJlNPf/D2ARDM5BkLLm7sFfEny7TnIJhMCwlrHmTxOxucFC0qqlfLeJxmypnddEirElBtfB
oYsM90401XOpU9AmB2lzebsX8RRcuoM+3i24IqR9yzxQGsn/CRf8CRV0/mgglU/29VbmIUtE1XWc
2WveOdgediV3BEfFh7skplnHNL1UDbJ942ycOpVA+LrrQYZ0RY+5AKG8ehQZPtK14HmzG/QPdFQe
yvMVEBHpDDr+dV3GVjpVrbrKeWR74/s0RZ0kx7pL6Dn9FNo4Wx5WXO1UzB+g4tMuLBoW/acFQwJu
4WXixpjwk/6fXDlL0EBsu7zXShv15ML75aULfes7+uNMMVawY1gRj55FJ0rtocExapDEJaDyXsEa
Dwscq7mq4XR5WLW1uJ35JDcKI/9HnJ6F/XateavQmzZj0MDo7kCLmsveaBEwzrq5RUPPEOlBBiyv
1yoK91yGAJFiyRHGNz0tRDEubaIIL83T7xcfjFn+NUZLRVz6pP6UMK74KO5qv/0bOZ5USF2KhNDO
CGvDNb9RMIpf0+KDVmoTD3NX2aguXlbGQzTS/3MGqng+fjBp4TKRl+wRtUdTOqx3FIBN9Hl+Ee93
Wgb9gsGLAmIQIE4eOsDZta18xJs+cys4HmmRbD2RpCRs/s3McAbBzxLYcofhuEyhgTeNLEcegAJJ
2/YtxdMSolBlf2T2b30R0vN6Ofrng8Fcs2rztFTKdB6FZVDa8SqopIFbEEMyIAmaY+xQ8Le5DbU+
l7sZH+By0mTn+1EQBagp2bRoZ0OOVXd6oiVrz/Ji4GEk8dKF/HHjZ8DZoAR9vrjo//s+DcQ7mQYF
CjeHgJA1mURBPTOO2y9C0piXdbsW8zQjCAkYlu0oOq7Lhtth++/RQZOnqG1TKB1KM+PvN4t5L6KH
q8QWZb/Fi3mS7C5ebhRyooKjGWB2VsIH8FSPCl0C1g/571cOWMlPzdjaW+GSaLI3P7+G55huIL1G
81PtW+8hYjFmVyL79eirwUHPfkMzAScz91bLLh/ARNDFtag3MW39hiiyuvyon9FuyNv7gokO6uhs
Q7fqR8i3jHpHzsgBXgebY/9edLqkR6aOkiRCeS/JhNaF+FSeA8BJiYaZAcW5Rh4HiVCWdMI03bGV
FG/X+ST5fHRiKcn7PLKqphe5pk3oYXK0eA+v6TGAVOenFBnMxFcftRssrpojyXG9sQMrymaf+f5i
92UoIXAFxcHokmyezzkNcnGqsQP4lzY6JATQvlmv+KOixHOBDFw1cdhSxhuki/LbdLgoo3ClB+3A
gBGijLQqNlsNIwa1l9WupsfCEKMpmW/27YA/ffDQRcYeFkdsY07WZt00pWXXOmL5EYXeZ1oFmDRI
Ckjqr0A/CwGIWYOLAzz7/N4tG0uxE1AHzGxukoXBHdhkfQF5akv+XaApQ36oK1yac+g3kB0A0hRd
Tey5fnoJLjbQ1OxIS5rfMTfpkL8JKy640RmB80PzZPGZq3ZMatodW0W850EPIYJgvZReSPQpnQpx
F67aph1gG9umDqVJkPfRQaHrCrE8g6cQKi6iToiPxYZlWTXwcAaTmYV865VWGJ3s0Gya9r1jUL/E
3YFQkayQzjjqzbD3NjSIrJqLrixYSvhVUXGPvMbr4fPj4kOy63Qqz9W/IHD/cnsjdbNoAHZVl9Uf
AQO2qsMcht2E5JiQBtYpNh7hsAdwFhi70MvIAGiMPYIMZUHk+LFip2aq69E0KTsdMJ0DtgDhPm+Q
tlmB8kT1keaX/sRGZMODIeN1pbixC2BXHRSUdSIZscUj/USaflsZ8VvUdDiNiNP7OwUCpV4f0kLw
VS1FfmH224/bQJAqSt6JX6zJ3CIrdC4CpvQhxGFaxHWMlGpXnUxmY0Ayv+41G7HBPgTjBDfpLK4X
l2+zv3/nRggxy88dw5E9AlT9lSrLQgDAQfM52hYy9Lvn0+iWiSxbXmiUUnXaboJcWUgpZfp9qbhj
AX8OvLNxVr1vmfaPcwRhrBS9u4C2MWuQOkmnsJ/tWuBYCX4ntPhelwez7LVk6Wbv10HXDr2N7SDY
6XL9LTBHngLZ8mGHL1UU/rzpF2pZjHjWibriAvAQJXUwf3rrmFIHHYjXLuowTR4pTNf332dT3kMl
Nbf+/cF+VVVJNj93NmG++Wemmvj+UCkdtpxj4gqNR7xhXEDcjPGYxAExtbK4jVrVDluoY0+ihP7M
k8Gs/7HzPX+1FwF9A6fXcgpOjjyH4sBLBPH6bi2eyES+hrYtaGw9KMdXAqBVFl4SytW8mZk/MbEo
jt4oqvN5glDkWaxWh5EGRAHO6OmlW3EZT3wtrewx+igU8425VEXVAt2FH8qB7/V0aITWQFG1ZZAV
z60EHR3L7DJFzH1Rf1Dhe65fB14TlwNNVXP55r7gcWGTTMzxqQmboVhaE0EcoiWaKS/g4lQFz+n2
3OdPP4Mv9PiSL1eP45D3LJHq77Qf2pBQBaHzptJ9VN/l2LaiXcdGKJnNzhFdXJLuhcDP78Is0cXe
+oQoQlb3bUY/sZG76RfIlCmDKrCPKD71PnnhzOPJnIBs8HYKo/ZGIZA3kIndXZhXkQzwGtnkLjcN
X4CPOVyCp2CbZedsAKanwByZL3vneT/FTaGl7v3gndB4DgYpjH7nLC12QQoZrGST+aPMHgOWpIom
l+fSX0KCDfE4NYpNlwm9xVvDCO5BVEkoSFvyxvKIkC9amcRm8O0xk7uAcbGRI/DNEyCHXx05lWWe
RwC8BsI9GUzBdDsVN+XEg+epeVZ9G6nFYg5513Fs8n23s8iS4miktx3rYO61NR/8OipxSCBG1VDT
JeUoFXEECvi15xTR/zHdk4eXA6neQynPWyycRCUyg7JSVIhoJh+N8eKlVLBV78wwkt8wGNDIAj0N
I6wyhb9qlwhoVR2wqlXD3A0EUPD9jrGBqcU/IEbCt95pdIoe8rV0wrowJF8ksXZ4J44FNFKL0T2H
d3Vf6977vk1DixDnj2KPj0bY9FlX1w+kyzcc0GIEbF/qQF1A4Z0fM9lyknQ05uwHURCVtB4FPv56
5LmmRoN0CIldFDryoUBhlLvsP+3iL0dAOjaNBNjyngWrVv9/XYLfYZGR4K3irvjFaRekSlCNcBMP
kiTUs4+tHUimqBm5Q+QkQJGnNF8VQfGyQJrxKPEQfLRkvp9vENpuwLxr0OxdnGYz05DNKGyftw4L
5A5KGwJZMpQoNeC5u+mL5rE+uOzvVEdxoDQFTQBOL88yDMcLtVZ5cLhLfikBljH5yrOwPfX7+mX4
rVAVBEc4dD7lH4Wv9fiwvwB9bkjVO3QRsA4QGdSgKFZ1SWPAC1VZGd061n249mCKROnCBnqI4h2m
e9TyeUwOxI669cwPF14VSdeXcZO2kR3UaOdb9ltyTGexVR2eCzhtyz9B57JL5gQlquVVCbyLr7Nh
n1yeCuvds/iC6LCHZfChDAHUpR58sgh/Or0e6CYATf1LhMrm/tixB6mbCsmySwtqx+MjBZfJ5b+J
rUBq0mg57Hjonwrmer9T9xhhH2pZLe9a8sly/gM9XLj+tlQs0vfAqjcSwjlQ+Yy3X/cAQrxH2/rE
M1BDLvtBmYMvsiXXGy3XNT+tqiX9EducD2H6X+cY6cxJCS6801tBYOlWxgx5HNN+CLl30asSt0QT
M34dKmKyHXVCT9Ede96toFAlMH6+cbhqOCOH12jx7HMS6A/otNFgEb66QdnIBsXl2F8UZBMCMQ5l
UK2pq+9UiKn0YqU7rmpJbfA/NTIFetpUfwZ2Aru0ooCVHaGdxzg5wn8b+UocivUj/38eNzpJZpqW
2m6Lp2HaIKcclrGblRbx3R33EzuIOMgMFz4G5NF2vPTEIbupc37OyjjPKuOMWKQnI3LebRe1yKDN
eUk3CQUcDI57DR9w3oaftl3oZOMhYpox6+qNE3iEjnzSWjTy0Nqu0p184ZW6YYV4yvJ3G5tiQCJs
b8wctXguGP5I0EEGHm95j2q1/8IEcsU5ELfm7qDSzHjAP3DWNLv69YZK8abkhDQmHFNE2Ap3o6EP
hfmn/Mdh2CZ5mqgerT+HcmpS9YXaYDgODtHKnW0mT24IBWMYE3N3EefvBT7DTqHcZkgMEPyw5AcL
0gdozMWnG+c5DT1zSEwMrun0VzM4nkBMpw5oh3D1svljr2j82116dUsHXc+wPArvJV5eFhY83bzW
giM7EE4GXgWgD5NDyrBRgnedCzSlhjxHCPqKH6ZQM8AKrS/N6/Rw2LzEtRd2iw5EKas/SAUIcjAI
Cvx+0KKuScMHw+FSboUMYFoMECikIFvGisi3e6ShpDhZlhrLxMinRyHriSnGzTJ8rJZ1dWZp6x5A
4IhnGsqW9UH+MAdOKfD+2mj6fns7NEL/4uXy8QlpSFeS9Dr9KpAptXvXlpKQOVT/F4UIwTZGKXVe
bvHt6vmBfinVDG7liW8xQCxyH8p5Med6kxXPR/6U4ciQAOJ3CmtEpmbXZbPCvg3fjPSwptgOWWMX
pK3nB5OnBhq+K1227tzZURxKiur+g2eDGreqZlCsIjvNFJluhRIqF4QxrdWGMEa2pSoDg+G/fy8E
LD5GB5XlcZRlox6fNPVP7AUYPyfD+s71LLN9ye5tzYP1hBiXE3+qafy09xsFKrogHSndprN2kfu0
xYPDWPbuvYRBdsik1ltDTFxPJV3B0KsuLNxZySoZR2Br3v6Uw19RfnVuSCLXvd7Sn75rHStCWnNH
VsATA9NRP/THNmvfN6UgJSVcXXmq6QESPN3hgG+KxBAeEuDz+aWV1v5iuE2D7VFVxa8iIqpPNSI+
13QGG0PbFL8X2tDuzc0g0TFceb9/qHRQ5+KNxz4Z0yUW+dmjC7QeN/C+IW56GcBY03RCDVtMFfP6
dx8SUjRu8bD9Re1vTiF1gm4qn+LYv9t0eog66u4ktuCO7EnyrYCdVV85P4os1On95KV25h2+kl46
mvEQlL/5TpJJ8wBt3kbyFO3BOqF/lhYJyWTQcJK9DdPE69nDX+F0jgc0LAm50wkzBpBOzfKkyTcj
3PLWYUN2bQ09iRqPOv5l/lOFXr9DvI1sph2C6QcOcI6uCJf9IxXM/1Rs7hKJYH8JdzvSJL3FvqYf
2QfRpJcHCn0vuc+6IPJtr+x3lmo5vOg4ZgZzWcVW14QVRaZETsRURUtvpCThoZpCaV8CNLxDliYE
aKly2OZXXSovlPk0xw0ECxQ48Qs8Oql5xxZ0m7szNfUblQ0FajA5Hg/s2zGQ0zOX4g4GVNcr3/Of
Qoi3bHT2e1dQ2uwoGaiHjLZfYTanwZbopnOaSEnGOnl8Uipb0a7AVsMnPn2FfP9aBOvqSAvd5saN
ZKTk61Xs+zIK2yqDfH9ckDgmBUI79lLVx807tL0nCqcpAYD51R1I+uXTZJ2fO84H0/svfMOkw9w0
ph+2HmSgtFFDtDaXAGYFaTtBnJWYxBpk7A3Glr7a/Pk14VKQoio+MMuA33bTNqhaDPatreLbNEj3
cZP8h6k9Q3hp+/LoJWYHCbgIMu3C2sTopuAftCasAV6hkbtBDzN0HqPeIiQ7B7I4ijrC+tWoXvo2
pM4CibiBXUGlkHXcXBvWIgHW52WjnBKIlyiARAy7/pHw21qADW1aO6MC+kv7vT603B7fncYg2IH0
wD4dzjChCyYRxeY+LEUTyUIFcT8DLTGLC/QQv4yw9em+l+8dAktAGNANtoAaavYYMRutiAfkLZBp
OGuVIYgWDqkK1Tz+mauXpHEPii6ETd7/ceCK2dn1H/bqnSv+6wJ2WWhdLHPtkqQaYRqH31HlEDNO
z9lGqFXpgWnvJQpL8z2GBVOp6seiTFQPtWKYOInTnMR+DOTN2zI7mMAsi7Rq2Bx29hYz/7bgYItC
8GlJn1VS8EsTSIrC9CRtuBkRXQga7rexXJaLQe3fJcZBDCrIhlHd9pJ8H68Xe0UmJ7IHJ02C6k3o
vZgJNsB0B1PtNSQVgY+dC8Nq8VnVOEtvvcjHafgmyvyhQ1p/awSMs7TEZPxdCqUwkq+dGif7VsBt
Q/CLxm3GdWYjeVetcHiRkPExi+8zRALWHDfhPDny2SuIj86gYXPi4LLL+xz5Gjfj2p3k9u5/cA1T
lQF+UL2SulBYaZOGyYOjfsNjRIcOcRcFt4vMFAkbwq3NifFrnpOKLP68S80fIBB2Db8tANeWDbqg
TFE0iIxw9szHey8u6fnBdlPTE5WOCr2hMLh7ymFNrJep60STXqBnQjUeFk+ZvmQ4qd8HP7NUangO
XoQ2C9aQcGEAzPo1hIxQYt2qa99HP728n9vzYptSlSMl9WiSIn/2EH3K6ummqg/dvxpWL9ViHGN7
m9qkLCGg6SJC2KFZs5Zt/ObmyDkWdRkKARTPQbRqluR8Jue3rcPf9tmE8mE60fAybTxSEXIrhRa3
OJ0n292lg5762mPjRim/PjTqsShPnFgaIS1ureaBw4hoRkNsajG8ha0ni0fOnfMbXBnwCfhmE3Nw
AkMu/9gi5oa0kUURNP/of2A90vXQOK5i4pVvX+i/wZL2HXPTI/7t5bRvWMEsF2z+vlYU/xHzzpQR
MetuX77+Y5xhTfj6/5tOjK2S9Lx92hPH9AIThBRvG6Um94PUgpQSXoNkVzy9Lh89+Io/yeqAZ84I
CDnCd0GEb/gUu60aKgP4B0uyFgFm4JpXMZ/itQP/7LFF5u2Lb5hBvoDSLwfA5zqzHPnDQuHKiwec
gqeRybK92WeH+poiVqYofK1DGjmxY8EJSE+CO92FnG6cRHQBVsMXX02Mk3WczAXlZCkZT2PbYgVz
YTwk3KO2eSLs/JtyZvrRF3TSqr7SS+uUuR9cHJIr31oFYChGI4IreYFdHjFdKYojS+cmFo94/aY3
thv3/WmSObF9/cjNQOFzKB0lZaJCJY9VoKvLEOuBUlJbEp45+UiaX88iK87uTguqAKFSwE9KztQr
kiC8vYoCQF/0V4EbGZpniX2eA/MkCDVyDJ2tV9g99d995wgGqKt6VL8e+JTcPrU2fMvuC/nivtpu
1IX8hwa0K81MHZwiVaicLQ4sRm1S7KON8Q/EEMg8WTH8rw2yuJ6h/gBaa/LPT/fIyiwGiXzlLlGU
c95NORa0eb8W2mKfiPRnEJNESsHZdfHA0eBL7Htk1sXiYV0Ig7LijY60KyXMVSArD0/xEdKVoFz8
7+sWqvzW4N7VXDhcw3L8OUQ7OGK7rZbYC2lRXYvD4EyEfTDJ5Cx9yWJfjMjm1Mf2zkAPtC7mOdhc
LzcKRTSHwO3LuR1eYPXcB0tNHt3r0A0JU9VWr1yuconO7fVd5gLEBa9oQH33nlG+Az5yN4PFhhBq
OqJZ7xpD2DdFPYPs3yWvIrUn8o+YmuKiz9UelUZtf23ibczWkfpE/Hj+myqWYi4NHpI4QPIrGlAA
Jrb2puO0QcZrZmSkk24qclVKm/sPjS4xk6WXnaFXHkdAQwuvVd6xzAkF19t6hEQSM53JFvz06jmu
rYjSGfYJQyg+aiP9uPrDFND71UJezha6sPcWDf+ZH0KU28GWz+hfPLQpgySUUfTiz6AlQBk/wYbO
zPsjYfF/p/IaB8cQchOxvYxXciz5pQRbwnSrP1GH1ogJAYK9+hdDxRPO+ujRDBQCAZfR0w30S5MK
Nx725xxWK8vW+p5VLTesSynleUPTnCyn8C5jyTkx5+V5HrUqCs+T7Q8wW+ZMUBvkunweHJrPjPv1
zAA6GqksI6HTODoYTvFb3dCmWXfWDvK7KU84v8lCD/VfhKAOXCygIe4yZkmF1B+SocN+VZgur5bq
gS7fsR4CquHB0rccxgZ2GRjlY/PyWLHB9dIA9tGcIoLNs+y7V/9cVHSbtglZ+Gm7VNlHPbU0Pcd0
JOSWP/HiLeRNn/IiPKGHrhlvGzvrpykbEd0XGk3XoxIGLv4hIMKR/3K0S9UHDVZQaA0OvpQSUQr4
5f3cHeSUbDvF/e0xZx300vWZd+mr8b5zTbpvA7iaNsxygz+PCAB5YDuB7pyoDFDClLlFpAgiszyn
3XAt5TNa1Ka6nxy2BlaooTN5O+ez/W+yvVMIu8UXD+1bbcGPx5VAcWp1xLSpKIgENKxRe3986pc8
ss11DmYQMvZONvwnJVn8LFDKwuVnfYGqLGFQLJ4DVhKgXcj9J6h7Falnh1Q8Cvk5i0at0mXAaanH
KAWSum6139dMFCzuZDVZPD+PkKNhlDqGU/KlcYCEN0ATTlZJGsyRvawj3vrbSQErGoolVP5lG67b
mQdXsOIgYJEQ+gyImdtNIgy9pJXXiYw9f7PrGaHCHq4cQYUne9oUyS5XohHacTwLzo2IevNPa06z
TMGqlI4EDl0g6E5pY69SSLQh3wuYavwgT0cfNYxJTdo5a4vlZGNDwpkt/BYNdKF7Ulra6ZyeG30h
azzFsW3xcJrJJD0XgvZWLF/B2GyHiyHOjsIiAkwbRjgzLGbl4gvwaAVtocr4QGMQvQK+ptH+hPUu
mtfdUeZcnGNgEaZyxutEc25gCz8+XuHnKHwPZVwOfJdSx8T1fraprk2k2TzECTvfrzYyWhDcbXpM
bgkmFHxDS1Pz3zrifR3JFceNLAjsgRwINGcE9yLx+y78EJPVra6uVb2ZpwqbVVSwW+U4BuN8Fx42
aGH81eEcG9CC1YYzV2hirEsljXyW3ZpQClpOLFPOR/zhnRRGI1Z4T6e51+SzY2hEKJT3MtKt9m5P
vnSM4zXVJHV4wGpEYC9gq0j9PwVmggFX0zrMrS3HW+RRkykO8xBCy+LwbXbQZKuQ0K3SJoc+DKAt
sIsYH+X/b7A2oSqski/N0e1mU3nZdfBZ61KjV1zw/iXhMzm3hEOTvzBpY1v/OFczQHY+yMHMtEow
j/V+9+eFEjNyC4BIjnajC1nKuq7OtSIoajM5bsz6hr245iNYSy6EntHJ4EGl8lLtfhaOjHL6mRjr
SLC6/+F9lm2TcONCijROPnTrmauNQCBaFHpgpglo6L5Xm/zHCpLwh+enZcFhMgyZ++eey8L/gOfA
8LDm1SkHlgMO8iVuBF7hXFxZkiosKDM8HNwz+vxM6rXEGTzt++fTBt4hJmXCLt3uXsB75vCQbsQf
BHTT1dw7c7NUZ62zgJjAQIlEVTodcAvffLsaPBgW8MKYX9VDWxbRaqXijSJePkHWRlZPF///EBRX
O0lSG+KHRvQUg9AIVdYEOXxJEBW41ausi6yvyBz3ktKRWWlE0sNSuYUeZuAmp9t92RDKl2jTOCl0
eZ5Nk57VsHoFbE1AGRwG5hG+JbNtMA9VJ3rnYruofC73pTUksWoEqitujTUrjGjG2uJ/OuEJvmYY
4dA+7cPXWnNlF46OZPr8eWPtVBKi4TYCZUZZ04JLitsKCq8u5x7MR+yqlYzgXn7ITHMZTQExANqA
pYRODwhZxv/3VuKob05DB/csaA3e1vXqvDkscllHP7ALuWrxvHy3Pc/YJnBdD3rl8BiBI9ar6l5G
MUpRWcnMwdFUxdG6opo8DWnIMEdA4wJ/bZdwiF9yM0kD1x5dm8TbMvqobdzVK0bqszt+FSxHCJmP
SRw7JTK533/wJ2X9ZISHwuw1eF1jSkyGqT8CQWUxjmG84uGv9YnG1vdojWPeUZ9UG9GFI08c1CyZ
TYT/gq/4Cy/YqTZfuXglK1jLg3eOrs21NWdhiEBoz9LMqNQf3M6PZyCgHy7cUSuXLBLsf6+WW9d2
kzvKAesbDY1IQhOJ1xY5R53kWxwCSyWAotfhR3pfY4T0tjT2PGF/XPnsQZRDhl7nj20DWI3CkmKc
z0UNl3fsb9/yxZ9yjQEz/FDmuNpVKrpNLlyopE8C9mWk1uWcG7QS+kui1ANecdHWGkvgvVCIbc+k
GuEB6r61di1F58whJK2wdOXkfB+ukyaolE3pXTX3yk21xwl4hnUj4kmOratAI3eEwBxfs3YVpIlU
owHojSXeMxOEt7TPPz1D/3nh2S9eH9qPIVZQy4gr3RB7LLJNO2Qfw4Mj7qV/Un1bHeWudOVW747c
V47qF3GFlliRAUV2ocXkxBtgVy/ZqmEiz7p7W8f7GVUg6WJdQYskhkoE9rINWLPchuO1itueCzJu
YPHaH5guUbUZU6V9OsSJDnW2GrganeB5zKJFmLwJNnRyY/fij5bP9gbBpaOUhEO7kR0XjR97+qsI
xgADoZgJ1Eo7djQFKqZ1a3bizFA+eFSvsRyiGl7GxomYy0giZVICyGQWxaCsrOqxMC4TyGcEl0+C
NAWiJ2CFN9HNIUtxWCAHW8kcaD86tC5mZrFPRAkzPA0nGWlMoKgFXNdDnL/919Wz4ZzDs9zxhI7q
ibJcbHM5+kvS4D4rN+wCMW5tKEsjMWUdHc0KKZxgQ661WeU6USetb6kOVIVQSImwROjSa0Ows++4
y6xqhJP9TN9sexV3R6kCf1AruZ9o1nr+xvMBIp3zvTnlScRMf6ps2Vy0EoXUy2oOWNkm+JaQFyMy
98XqQxlD3lW9bQDMS7FS/8eZOhi4w/4Jfi84BKUcgRY9Ma8VYNZAaVg1o7Ja7L26HbepXABfGjlw
e7wAjf0gEMlHIOPnwLcqdRE5dUuPKWj36YkOveIvUDD23MGGkLgYGargEAZcZl1nTg8jxLiDV2dy
pdMu8t4CBr5EHDzipUk6WvrF8PxF1h80WNstZpdvEjI70VppOtebw2CerdNEwqxuCzSbwqZoW2s6
ffKCRzG8foQUInWpRoSKZ2BSVhjExhfUVhAC5Pv0fV/MlbOAALC//PQzNUcVREjaTpP07rqx+zm+
Rf8hxNvcSkd4Q7k5kFLq4ptnhduh2lVsqcuc6pbUGKdu5E/leIbX/aR+MaFd3OyugPb/sqaJ+9Ac
EmSgKSgnZzoam4VrxsHb0HC8mVlg+ntHhGz6XohkY0aGOOYbHRpzg8VZZ+8ThahNuKp9xdAVMcaG
/bNZuc8tGBTwOyyp0oSjeG8tVTqsV6KipLblIu2x476pxbWVEGPjfDGwAZk8J7ccQGeOa3qcUdPm
EBqRGsK8GYoS5hHsS+WRl/HtGLSU36I1AjV79caGG313PmL/AorPSUBlDu8lOfBPx2dEYYVXvLoN
l/bgWv4wpddL5Iotnn31519U5z6FLDvDSgqfaDt/XMnVVvT8/BPCvdnj6PY+o3Jty19fBGaT44u3
cn9GVytRh7BqJJWvMUNOcK3n2qCsz9AS00kiCVCLldnnTQyrzP+hWliAQSpWme95g0A6ZqsVTFF5
bl1FvjN2SFEzn8XN3jDm+VTXjdQpSbAUPsVN37Xc2fREOIMK7iYwF7dKIOus8AFaeAu2tZPEpP/M
yU+wkxys6yh5Sr5/79XTSJQjJRFAw13K1j8SGfjjyJGtbdHzXTC6L+CazMgfQnpNjs9S/JWXDd6J
gu+UU2WHzbJLRz02hWrdcjv3kc+khFqzUeIL5yeRi5ryhaXhtNqwfu4jYxYq+Gz4vJ9oGWLYO9l9
JvCsTfk7mWBZLBgMu0M6u2siYN5SpO2+D7RFGOsj5NVYy760vv1IQUNQGOAihKJkqnJV0eCLLnc/
EI8ZJtsBOXYAdicbGYVpoHfAK72ypVy9cRmBeM9T5MOwWLGxbUkugwWuXS1S0W7AoIbNFDdIXa+B
azegWgP/RrCLmVYsOhq+EiIqBVGFZSdoku1tJGzI4N7CxTSVDss6MtcxqVz7QnjiNwGh0nngW+ws
eF5me+4WUSHbImwU/vYUdmptVqb6FXMAOpe40QccrC474mGj7tVHL4MvCu0GxNZgOhwBhFuRI7BT
bmg60jDUQB+nTK9+RRFaD3wgYoRZ7KHhuS1Sq5lVIZUofzVipki1eVVka8ZcCs1l+bA5nICnEPQV
+B7nGaV8Kleoj1UXFJieDRP4vuTn//uboP9SUqfHYKg0GFVJtZC8nbdqLC3j5mKx/AIO5m+/g/8g
b06qip5J9XRa3c5WL4cD5UpfZAPr6Ku+tDlazaz66u8PoR9KTiBC1v1bdIlst4/rkePi/xnTd5ub
AktobG58RXlteDgL8zOwMRJaN/f0lj99uq1U8jdmeTqhyWR4VJ6gf/QRrJZVhp3G/a5arptzWUSh
ulRv0JBpiybKA5lXgNNwu2/X9dRNH1pazufRIRl8mQ+FJslXWYhHl78gS/wEaiRx2G2CXiWE/ooV
6HSRdNmIBrAiyg42XLiSWdpsiYtSQNcSv0QNpd9qNCJvOt4P1qwJ8x4spYN2zXhr4nCu98nn6GRm
CjmAzZzLlF4pgcVr2kR0yNOoQ0JIvOd/A5Lb1W+779VDrv0s/22RXZnYIBtoF04GMFbZZ/eqmAaL
V4NOdxII/yMyP5+/ySfJ0nPhM4GUC/H1oyh1DGNCra3hmKLcGKENQy6Id2qCYYjqVXd6hSEAOo02
3UlKRgC/eZ7YsF37D7ZeWf781ORWoVGebJd/UVwmP+bnSaRH1XdFzycqKkxYMo5OqErnupsEJj2j
fMr1Gk0dv50uPBJ1Uoj7e8cCZSx7sfM9knEu9jmVZuLfIujjiF0wST3Ar8URL7FQKav+oQl65FeE
5CGeggbW344wgUeVjCsxHznmjvgrCCVqHL5JdhDiI3ZZF4DaWwGScvhlNCwra2sdU2JmwEE2Xq+v
LSE3jRu7TyU8cVBSmVoq/C6PfFg2q7RC0o0jff0O+SyTRcFIe4c6tMv5/KCOx3qCF/fGWQ24SOXc
rR0FK1x8DVYBWsIBFMmPrgGZMRaUI3myzL68Nv49if3R2IvpnilyR2yao5WrUxQXxdggOv/NJvdg
7NCrVoY0FRxjF9h91CocdYZKRUFBz6ZBQP7JTj86qAeyl/bHJPbbwZXFZbK9imt65vwmxBxyDUoR
5p2fp+3g618nLWeTcRRzIcKsmvbfBxfR0WXUDzVQF47rRDgMiRYpVKhkSHlVZRLEzGrzVgIZEzYo
yY07Ng1qG+3GwoKPMCzVE4iGeCOxnyVggyb8lvOHsbiZQKY8jxtd9SSE58RDlZkIqZJzQ4laoudi
fDh6sW44k2ddzeTBTbV/Nc91xEdSRqb92HFJr47ighluuS0aY+4hH87lKzzhUcMQ/5fkQBfhQ5bJ
RbxBuu7iOcTi4kV1wif9DVMFGhWYnz5unAW06lGjyNEK8CVcoEinlAGMTX4DMxyOi25aApHnCBvz
cgvFsMhfU+pYTsGfSMm9P3em/+kg/5sVSgPWqhXSkdzxDtvqv9+WWJ4VDLMl1B8pgBVv/wgiYNv1
JkMdXxyh3D5GTNiktp3SS+Bcmgk51WqYOlrfxLdDtARsVW8kQ2b7ps+egpuhKVj5KDwdc8flxxcm
3ckG9luAjLrPIuf9wV50cggkbvq7dIZLwB7lxEL7gFHOm/QiXb1jGaj/AI+rVYLIWCVJB7O0Ie3C
x2dNhARg/8whEdar3pRf/WQKbp7duweJIPWm+vL+LzV6gRBpxbdysMLydkRF4dvOFd3rPpgMMgwU
Ek8tHwla4RrW6hKAd4I/Sb88F9XKZb513GINkGdBTd3x+wNwgQswk2ajdiw4ULKD6m5kj/VBmCnN
nJPn5bvGr+aG6CxRXpzvqs7/5kUUlZUXU7Z3xu+GDrN27uREliB4p2KGFidXWuOT3ltcvhM2FLeW
6rO9I31RzBdvJa3mHtmgWlpQcUqmCbD+t83nQNSGWXdAmdl3mFOr/2TIHqSAvZGMFA2RoXENvS5/
bHpS5LueeT+ZJ7kMYsxaLvS48AOMmBAfPXN5dPn8gRi2I0qJ6+HiMAj9/KRd8oFvIkb0ccvYtpWn
aGQ9BEiv6dy11DDCmbPZnHjLx1YO+5WvUyNDFzocQS1ruM18LSNxE9Aw04LaeNx7aqlCrj2uzy39
Oi8pITPvMgUhTxdjExRb5TDTu7x6Z7hN1LYog1n/P2GIFYVlZV+rLNKq9xDwvyDlA36EFawawhSH
9H+gUuuaQS4J8QYN9TjzAHhwI2GK5l7BmLrxipJELgTRQm5cM/5ceeEdtzXPkT29X7y704ncquKT
rDLAVdCtdlP7hWHsexN3hbZPIY5tygv507Y5yRQ0DlVDzdGxUfRfbyZjka3/902wf700VgQdJc9l
jfgdiqh7TTw6om/2o98OB/gLw8Kk3GH66ImznJQ9rARwLBgZqVOWALfG0rBIFaGiqox8dmmQzfnH
uXS4x2RL4v2s5ImuT0/YSS+lte3XRCJ6YdgEfuppXhb/25qcNFHkxpt13UVI6AmOYWlT0yyHX9nJ
/Dr1wVJ9Y0k9ecTVhtu+iHwezRV+fvYm7ZzRUIYpdTIYFfyg6PZShpbOR3QMv6LhUJaGtsHyMjbI
oReEi1ojGOmeoXcvOP2B7nnOd1qza2jAyqRqHcoXqQ1LWv/7aItLAgDcZWJroNi+CreG1cBNGoft
ub7CQfnbb1awwy6GqL94CLLmYZMdyivShQ27G1Kr2/Anx7pLGVu5gD6TFQce8C9nRdQFCCxNZSqL
Tf3StZWGzuQ5e3x8e3xaYtVSHdoeZclY1refON/XIz9NKd3I+iN3kxggF5ouWf2XGwsY6uVq6Jkm
JnzrgYILu4wa0JqONg/RenO72JMVQVpM8TA4FR+yZRVmxFWJU4CVMOZuwkhViATuHArBLA/LmN83
HwAX4HEhJbZp5i0LneNW7ngt8gHaQ2oI6Lbmg8gYZtKm6/q6RiWCvsK6F4o78FzT9/ACt2JHQDiR
RhZWo1X7K7vIreSMoe4dtywc/g0WgrGRfk9pcM/9tjeNFSZZOjMpGDSD+Q/tQ9Agj6a0NPwIsXGI
8pE9c3Qi+Lapl4sAfOO0DCxvAGq/6KPqENDmrUDpwkf7JyRCwvH/JCs8BnDn1jPyzHboC4I1ts+U
Z//UGUQWkZQEnX5X+0O8COUAdefvEOjfu4BywKQ5ygwJ2u88b5hmN8jGagjICr6px54u7awfmCH4
+Pi/dXCl3Galw6cUcXklIQ+Z8lKd0Jvzl50ZvRRlx06T4iwTDHwVpheTdl+G2n+CjhoCGn3u9dTY
oQ9BX+R85OQYzTk7zL7weQ8aKXRaeHeE9wfhOE9HhJLFGHCe9+i3L/0tMxZJratj4fPO+aZpBNcF
9ZNZnjoDTBT9luvIDecJeuo12sFsin3Kty0RDS8et55ygGhgCfdtOoymjXYQ78K3LD7YJyQ+CDZ0
ckYq3xrz+Po7GSiMEtQ1bRX/W5btlMw4fPkXNsTxbMM8Ge25uc9GHIMP1t+x38l1W17JbkI1x3Xc
ZjkW4j0XzM2DYAUtEa2KYjApFY9mcaPau6vJ66vwN4esK46xqX0ttRX0zdduGjkN73AZJoUlB51g
e54AOV8J4OWfefeEDby708BQEd3tKghS30BvoqRsnvuCoecIClDWE3jsx8XQr9AtlEoJHNiyGuKL
kiFJ+jq+3BRDVNroAxf94Ks7OXJhI06yromiUmiftxsN4ieAamIKidKuzigIVxeCHSMWQ4guVaxy
9vO4ovJ/yesGA2O2s+Ssq3qNv2WpzhPDtBSiKy5zYGmqL5bsq+ef+f18X5L1qVO052y1ZQwfPxE6
3eUc/J2iYLvktsQbIASUXjoqXFEnmmw4I/bhezcqvqlLVTMiEychGyhVOPqRGuFvrP0Pw3MakRPT
3UTolSoLiGN5NFhmKk4i3En6UEK4IWzaFgqi9YdR86E4oV7+isbdm8IXOs0VmYqJh5HpO7gYemgV
vsnUnhWK+DGny2Ktb+ysbcABQVL6seGyp/9vx67CqFwBi1xUlwIJ3MOJKN03Sv9L2hYhVz07q1Ln
zNsCELP26NlfDGqU6lc9Zjb0w0jHt1RWwb6BTGxUHT+OOm0b5i5jlk6f4c15bbQ3hHJYbQIs2PY2
EgCcYZp3yLVf/3cnrW1hPt32G1tmj5sGUHDFeYUfxdGHNccxbemIHBq4oJ3ZxYX15eUqiYgm6pRk
84X5Za5qKn2/v/P/vVpPgXYXuz2n7AWKF44ePLRJd9UGIBg1GbFuxhg3PHHslukLTwPUyflZHqcB
M4hHWVjOw9nWMtkjghSBVZn4u7p6PFD9HVgZUdUevOgai4syDD78PNfbjT7SyOpoI9Rz9VneLLQa
NJxYINKENSXXjF2ZhjnuCYlEbEIRLi2GzKexPfNut1PbEceB/26+2J7ldxN1DDWKtA9M5Q0GoXCj
+/xB/xj0K7LK0tJDGhgadXpljx64ykcsAvDEjf30JmOkp57cuFar9vc7Hb+vQuuvuz+axenY/sNC
lkrSN9dNtDFedw9bF1AnjHYDThUQXDthPfKHl3B7jlSuv38taVtZ09r8sPDONWPfHCoPJovP84Rk
jo/2K/mx37zo+Uq6UN3IvZY+1AgYyI1eT/zjwH3x4d1g3DaqdgzEfHGR05tKxjGcts1rE3lHG/0D
P/rmFkBSq+Bnb4/t0zbbrK5Bvdw327KCUFXp4Y79NlX6/vNqkNhT1hMvzBRoldb8SmLxLBuycY1Q
OBsqSpZLO9xkUqRWyGZAaLPH3tsWXphgWz1UO2owedPMFaLVvSt4y9hYGfeAaYAgCWxohDqJ9lAf
DyqFGp4JzW/8/iRMaBxC3hExcZnL6AALY2XACg/oP1Axdi35gLUV+cSL7kOhckI3eEfsX0yeit5q
VBmhXfvAcFg09K/lzvCZqyDP4OuuUEKakCMPJxsQvMLe14m5sfVmJ6EqM2rzYGiNVNeQrU5/zPEa
JmQes2SjDUH6iwbnL952ZxMaxCkHvtkDXKdE7X8hChKFrOMq0gY8+w//c9Y6d6JM4vrY7lQ8NKi7
ejQU+2e5xDqEO99chJPEt0mchbs0Yf9IEDzJXo5GsT1hP/K0Ft0LK+/XzbjaZK7CEuauIVLblGL4
/81DfeII0NNcRMWAJlm41kccL3AeDNrM1uF3pOdQM3i11EuG0Hyae2gZrCrz88A7ovmf5qTwYPVr
H58yzM8yvRL2Q062iNdWUiuQ8S9hmmVe8mH99uBQU0dgr53tvL+WG7S9IFBJfQc7cyXeY8LysWQA
UyLENmSlb27NgHIIHn1xYmHGszUnZFEcfymy/SIEd4G5lFJ2drqacxeJn8NWryWo+5SJZIuap0Pi
3Z02lGeoLIEE9QyIrMzlyPb9FtSPRjzq6IeOw1bHH66ZoJ7w8Y+LWoXPM8hDJ2kqrinLqwz7q0xG
x9HI6lG57hh2Xp5YikXyYFQZJW8HCk/DcOjuIi+3GZMtCX2Rxo2sfrkGyfqTSbuXzzDsQZhGcoqZ
9FiNCwxd1YvNJzDVLjg6Fr3+zwnW9vGBpyJ/n9pxe4ICH5vHe2bjQGek1tcEXL72lP5i1/QFnAAd
HYdKOoz+AMULEB7xEOdZi1WU6SFzyRCBSY87TDL0sMsQLPxbzcdEgD/Y+R+wSs3L6rnE1qZaNIAk
alIiDIrLgjEv+DWjqqnMwuvlo1Jef/OoQ3StmMOYEECFlxxpeVYtda8FGRLA/hykAHgzYWvRPNDV
eXLqWlPl0qvsLAxXD9IUG2GUF5kJW1E3iDNdGOJs/th1wFHphL1pjFwwSKmCAiUtL5hdBGpmXcsn
iFCDqRsUjNTGQRad78Z/Gnsw1dOP6sK1KfmObplQFt/HgFJ4+L+uQuCwaj1QFHB0LfHDoW2TdUUz
DYFrlXfqWWqTqpgL2mVf+l8rxxId4Hb29BhUOGXvWXXsmUpf3iYjR/F0X58CUPf3fj47VAmnYu9O
EycBWm51JlZ6FTAdIPurByQ27NbSJKP9/mVA9xQphx0XhzuQM4bsRaDGRAaVj0+3lIPcqaYDc7RQ
LlUf2AuxPYGq3skXGcz6YEi3uLjFLr7YSwee5uLobxeuPhrHe6BoBBKFaPgfhzAq+u8w585umZ4E
EJkcNL6JvGnR4qTOF/Y1bQQrQ+2rDe9+JB3SoBnhRVCMN+72IVpeozogGrOqhoYrWmWd4vxGus3c
UuDESOjW+f8F25W6vxoQYd6tEkhXqqqeVsemGNPdhOFBJMtm8Qz7wC8UzNciAQaZc6wvqQ9qafgN
GDXy+cIzluEa9FG8lxOeIpyOdEzkmkCTlJlSBeAyVQUOS9oFaMYMq+LPCU2SEXkdQfscsY4AULPu
pLd0As2LkyVGsuDQaUyttNTHOlgbwQ6wHmRkbykaWeV4zzmakC/D8SFOoF2XaaMNPymULKoZkMzi
bCMPZk44STNaPX4oy7sPxv8I3usNYsOFNzXsY7yb095X3lVkHfOXbcgZkRktPdDqjWL1Xwpl/h1+
JyOivtXfABAxWJogz2LAXAe4bvRVyz1wPvjjyShCkpthRpjjZ5j0HZnfWxl+/ir1cJiiff82OVsa
3aHz7+f+3XBRKkJTLEkSKbBF9MlFwHax8oCx00KVZnm0hA4OtiXlLGVGTDb6oPkdIj1t/65syqX5
FLFzbJHxD0W/DujVAPwKRwizFGGZgLoIko3PLmCDFRHHEb/yDaOKMpjYf71Y9crv2Jt8S4T/oph5
ouFniT+cCdyTLHRMgpoJdYyoUJ/uyAAOBzm4G6krycfgDGlfUOHViBuzuOrgHDXj+Q5sUzC+vjEc
d4oeYMLaCb6JTVkrYH+08u1yd4L9P3y5vL9gGjOMYXMaDMuRhGGguO++2A/IK80p0qjkjSTKRG+S
KZhH9JCU+puagZXKj6ulmwFPU5nScfcJKUzak84VCc/rPUehGHd02BsYC7WSklukLKhdRq/8zfda
KIxpImKmFWEzJuL0HZJvLIZaA5k7EoI5V7VBY8zidhy2dDJavO/n+hj4i7sveRfwwfkzQMxIyi6y
cuLdRDSRccaIJnTTPuiWstbBffHQZ24V7uj05xRuGbf/MPpE40OZL8RmuGl9AKLNYTJLGmAYTp+J
8P6OKXEbjY3xjhAanAjXZMdP15lF9+MVPqm6fghituUs+LS9l7kAc1s3mhxcGATX7ByoiqEaxnDV
DE8IFy0BSBHjMj8/1r3/LZX+QEwm/WvK5s7xYgtF5XItk2FgWWKJz8eV00aCBVAQLqa/t7cYR+we
Q1sMYI3xHN7Vl6cHy6uZksIc3z93ORQU+dDy7+UEbUMfeRRRkbXwke7Nr9gdtenHsYoxACLCrfHX
Mnb89hxr63iPs01zEvD35VBjZT+nv5Ef3V/YyWM3aN91cadTUPt5Q46siUaEGOIbAT+HznDac28Q
cdq82almFO4U1pk9ihOioBkHTQs2cJO8K75XIts42mpC0VixdriU1icY6qylaKFj5idsa8TaW7/r
PXwX/Y3sktl08zqpJWdqTWFP43ZI5ZOedMiz/a0iCUTWrb3PEYlYpgCr+KbB/mlq+3kxjKofmZcB
54gXrXCtU6UM3K6M0pG2Uhwe6hn6YlHfHKkhIW4WcEWgoy18AqoB2IPiEvSHErFGwu5IvTfxNZaV
2MjYARMKNkz/E1AZFI5QAKpPpd5PBTqokvoeXHEqJieTQL/4DMqul8rHpiuirFllEe/FNnM92YQT
Rt/tfwShY0UKT8P5MDsZnkBLSyZZ+fYh/hNcGG1zC+K/e8aYQWRYe+bD2ykWJoXB6MPzQdtJw+AW
cEkCLW+RTixFHPHdf9JJX6ybGyiDK178e5RtjAvfuvdVP/WQiGNo+1s30v/Uk0jOa3BtcVe5Vegt
Pl3vjQdunNsASSrn8R2erV86VnJp69buvBBPLWYiBkeL5EQveEy2Q7V9pYOc0w3PJi5PCm7SKO5N
VOy+rdhYzOlNc5b5FEtph1dKIeN+5yGXBKLAloleGUjeXPPUqkgx+TKFLFnsheEtL+Xff2ezo+oD
Ch5nmsm6aj/JT95LESosb6gHLJetT4h1ywviY10jTvGoGkYn4b3w+7QxlFzPetD1nS1T88vwExld
0igIyISYN9pov8rdFX6Fe00tnyrvtl1aRr/xIez2TWVRE40fmV1/bHA090zLnvgsSQ8S9D/QZWiO
/uLgosaGLrE3cyxyQhPoGFzy4uzbmQQ3ghJrR7NrKe6NQmBfS821CuVLNclYUc9Yj1Ex5IHGbpeb
rv1jmVUIqmR4ej4+ISXVNbWNJCnKzdyazQvj0wNrc78edbEYXoNgv4fcTBuFoQ6MvJrWxKyn08zY
88JFYS4bgE1Fy6vyJC30/R2bbqNbtwayWKbhML0yq5nexXZY+1j3hbmgFZRfKqXOdFaXjKKbyQGO
ByUtb2/EVSBz3J0XNTKj0p3VAbw5KXPouC2+dHdxJasrqTz9JBipE9RckRgI3JjBf1jxpthI8KOP
IKgdf+DfzVte7IKZhYqW59knyZuRK7qDl+p4YFxYhDxRgwHoM1u3pdC/bzUW6q8QDMUuO3Mxml/G
NanCRdPNNMts7lzahuXQxPkR9uOJr/yGabDNv8HFr/qkccdnDsvcOOG5f1rKZUbzWbHePiBXnFwH
4e6dXwH2uoBtjq3X/T7Ln9cUVUVCQQA038NLT6KEbEYW1rXkzlDEVsoFvUxPv1ARzBhLaWLDuZ5k
vU1UJ3y04iyrA/zh47GoF9jOj4yOFs0ICaKR8Q2VBBOTx5X/e/8U/XrriYbC05xCu8nuceTUGR7c
LyX+5jrb+bqX4mPEBX63zwBhQqj4D5FoKQfBvfvCxNoYTUShmtXij6T/6QJWXR2FbfJh9ndlxuKl
+nHIQarKYEP56gP4XQyK5s23pP7OIPudlAQ1tnAJ/Y4P1SAQXsl+2KEYPibmLbkXuFrHiQ8CZ9JT
HFduPpcIyboeUMV0cdeVU9PO7O/8n0D7reDMNgXs7HmsGvDrAz5htkM2EkxjJ8Sx9wxo45gwTE5A
yWhgOKJJITQVHaV36E7gfkGe8fQaElFzKa345SKN68F6KrNoQ2mmQsIrjDB+7eO7Kg8a4jXQtrJy
paykbwt+UXygIzLXrpaGEcZbhRsbq6YLd6wI8Q7dOtwWACixxcrbtbnK20m71ju0yfSHjS0ryxyZ
jBkhdZzLdh8HsrNEudDVCQCkynQtJZb0d9xYCswcmRu682zDOYHPPJuxNG3Tv8qHLRc16l8Nf9mj
XqDv8nizVbD95zKUZ2WWZV0TqsDmrKxPVedm6NGEYE421WzZ0JOQyPbplfTImKXrm1u4DlOlCAhN
SBXf1wX8XivXBz4my3WwbJhjeCe4E0TpUcLASQ1cDMxZDoxbaXHaRqB/nVuefoA6YcVu5C1TNOhY
1EFdxjr51PS0BAy+k4PBE4zibR9bLoKzCV6g3JLKYHM0X3J5Y3nttCZ6KlkToHL6g/gTusMI8XP8
bFb+VMGhvhFE77OP406wgFYbVbOQw0t4r5NDa8xEIM3OFSj63U3wMJbDztmvxVhdhp8lg8wlcUXG
WfiyqCypru3jTjfiYPViTogozz7yB9U1azcsDQ0hfs5gbHk0M6YJrpjgXlYpzUeVH9HINRcjnFrO
Y6Xq4swU2ur+wikBUAlYTNowhxG6QWmZopARZ5Kwl/nHAlo8CkoNn7cBOLyKMVZsWWO8Bphak9y+
8sj0Rr1q3xIwULD7TphrrclOG5WJdpwo99VMu0YkEoILY5gSXAPiFXJEFvJEVBAToYPO5xlV5fSK
TT4ZmX7v/I2mO3CnLxn5rUZtUnW131DboG1F/WWoy35ovTwYjNpYWJuhP7mLXH8FRDFoB5P9W2/y
f1s4dPt6htj0h9WPN+qX7ivUgVTBH6pP8OwsvFcNZ+sPfFfO+ZyrylonA2UEs11kxNhutpUCXPRm
tv2KMKekh0M7bhnduxxYuBzO4KRfyoEcXcEitn2YczXKJ1UpeuXkYOhVH/XhpTH9BWKXb25wVyxU
KCpXJLn8y59iix49fvDl8M4ob3r+R7FUtm/HVuZyB7thWc4Fb7SSyrmz2kz/eljSrYFa9wWAIuFx
lF+MeD+60rxfc1ol/oObT+C+gwz4s7+UHBeK9GBzPd/nFtdXhatJyn0ZM/jCYqwoJJME/5AkHt9j
N9osRkUC4FQ/9D/tq0lvEqV1NowlTBWLo9TZt4pgK92dnkRKzwGEuSTaB5fCsy8s97mtBWDQSSrf
y6FxGZMkLlW0/CDvvKs3NnGkx6LfRjtDlis4+AgEy4bNggG267az6d9p9yS28igZyvcEqhTbGuZB
BXLKzX/rl0ROCeYTkiAtWWi0vGeEta8UIVKAYYjuhgHDnHaKb7qPPR62kCVF/wWfONmnnVzZcZMn
x3kfFv28ZW0eZkvdFyEPQzqEz3XKaZW1+fBSFX9flq9z0M82tMDPc7gSLFsZf7ln4o8A57Op91RK
v2wLkdwtKYzA7cgIzk3+aHqYVdl/FQPr1rfQbKAlvjwwZoqX3a8Z5m8PQGwIIuO4K6EWUpwHr+uo
yTGrs7/57dVA3WEYJwgeo9bTNkWGinAFFUzZMwfuD743Ty474nDIl8ma/TsCijy9i5kuPYVb5TrG
i3ABFFgd3f0ca6hygaujyThwZCjLQKKOdtqhdfMWv9i8kCdF29nBg7HmrnAgVmWFp14DDxb440ND
Vxn/CiEDqZq3/b6MieAAn3qJC6/A9pxtjZ46xVhnx3jO0B8lx9OP0RxCa0+MgdYL1gqjvIB73bu1
9BLG01uCFxMyzAjYDycy67bX1vaEUCt4vDi2MTQr7D1uliW9Rel1+yJaWLnQ86H/nsFS7+wOZ7hl
g5iNU5DlYVh9F7JvR4iowsTo6+UiTUOkUuDpNv9immF/1ERlf4Q3GdZ5Dr08WSrk+g4kcfvQvw1z
RNbtKctzNV31RZd+O6G9kUZpBrBQZhnEqwdExLpv+TwiKSmOwmcrZXovHtzOOamTAPJeLj7tFAsC
owosHXeJNC8WZqwHszoN32F2P5MA8z6i+VIo5RR7iLCafUHy8f2pqgDb2c2+tds3bso5uOSTdgyH
Z3yULJaGjG7sPyA4sivHOp3awYcV53rFk/8Xa6oQ7sNNe71IU1e1I0b7wKIRUaPJVdNij5D2Kt23
yVARofI0fPZgc9sc4B55lMo8z3Xvt7dG4zmXq8FbP+4c1/meqzLKN/kztYGpfGF6jfiw91CrltU/
ONr3jPeEFFGNDBoFdd8vmxAb5iW/OS3H27Nse5NNVLwhWsD4jgVtqwQAh1OJ8Pu8IKQfPgkeWYkx
g9428P3wSuPk4Mf08oOALtSdBj30l7P5WZk0WS6u/I/1Ia2l8ikaaPrW/AyBBkcvCd+kQXnukkph
R0mBoQBzv/dTHP7BhIfM0Zi8J1wqdre1DD/UDWeWsYb4u1PFfyQKRoD6A09RbBGO7sZo7LR93bfc
RhnKdAsFHJuz08Ax9r2Eij/guEQdXTo2ha1cjMvt3xZTNc23n81FfvhsTMqr6RvjvGVZpg/Div4X
U4GpwPfwR9dTDWrzjPaxc6Wr2aPKmvB759l30NzRUr5EE3AxSzpbBqUfGxvPWAR5vmbf93WRJXIU
jAtgJyZdUPVV6TRIBh2QiJsKYH+217m1WWbqZhoAKHcPkBrDFU4t+jd+ecZrVaVNAuLeoqb1iFSv
kyBO1aL8SGVUkoJKn5yhfvFgWD8IaB7qKBd/grkINZrUfA3uppuuZlp43YMkfbrj85Q5+57YD1Ys
I88vT6LvE3rbcrNPgIXKjhlCTYzkHI8FAG9FK9vYSNAj17/Lp5z5x01UFFCb2a/59ez/u3rc1/oW
G8fVI+Lzy0gJ4SUC/CSNhGrRxcy1RY5sTMkEsoHYyi0OGtTDX+5Q4t9mRzb/lP8bBm1Dz3jkmECY
jgaAZnRO3J5Hi/T4aBfXyYuCIbpwkFZ1fTWGOSAvLHIIHdxdH57ECgih0R/jKfREoYYSlhJojEMX
cIM+5n5PMYYfJ/LkOYgFzf92QNG3980PEP4N62ILMNfSNj8FLM6c7ziPOrBNRd/vd8CZ3aFz3nAA
iO+jMRJRebhIw/+uLXffdqwxH5NakFvkUZImr03XtRmC6j8/yImT5k9u3jfB6Gz01PUeOR5lE+H8
CUTecjgLkytLXd1xaZVGD5pSt1VIN0SSRbvgrjK0HePwGaQDZhk75r5mSST1Xq5jkau+UPOcuQ0y
WC1DBVFco5kkyc5/PsCpFLvib6NHm3Oa7ylQAyUWsGVN6/uXDGlaU98To4MSTbcs+JM7BP9bKg5+
4GcUwDZ5r6PMw7I2FZVnhYzgaiCIafFlro4bgAS5KgUOpesJFYGpJOpcastHOCN/XVjaiqTV8wzL
X+T8+k+N2wSvib1hHQXkQYj7p30gqfhfpLnCGXyu2bZX0tVFIb2HkS1uumA/OE8+sIbvITrovPJj
rH58466veTWbp60NTmemmA3l7p0gY4tYtQdmT9OepM9jZoNiu0nyEWtMiACFgFEyUNoGNBkFGhDh
CPhagPMs9O50ejUURnVEer3cNXYTNorzkj/eXhirI3j/Vp0gyj+W5pE+z4pADkQVo7t1HjOid4O5
3NlB/fwSQmorvZs61FZ0T42+gOs7Uz5f0mF0BhdO9RbtIHslJAsATm8ND339WMvyBJp3F5UpAage
5zrYJmIJ7CxHtEcOi2GxouiwLKtFQl1H0fh33swGSoMNyar4QyUGzfA7tWzoAuExFlwICunUsln8
4wiB7JH3pwboZaoiDCt2MqWxfpfjEa6543txCi0gDbCmrTmqTycYKqwZ487A5JE/5+qQWZHS5GYi
UdHmKZ8tcViDRK08h5f/K8uv2cqWouUy7IeHNT1jNwKB3tPcIGwoVujvMN+IpfwiOjRNvY5gS8lT
qLTNAterRwjh6MyRXvo6Q+f91puY7QMgrxBTzWP1jCHStLjwz4ggt3gz45QeJOYa9D+tj9LjlrqH
FqoMRFF95RFLUrlp7VSjJYNSnH0fKlkuI6sxgpM6UJ4QdUp7yHuxvwfe6KoTL/GiXjZ0zjEL/tHh
Q0GLlz1oDI01HsOrP+OiZtAnEMJsOz7J8cA4zuB4so6G4CuWsfZOggI27jvXNtFiOJZYZxeGN5+Y
hcnXSTtf2z8jQRu2DxXO3/uCXu2Pt4yLdZZK0d9Omvj1xQdFs2Aouqc/HNGSyh+4o0LGG9ntGNwn
PT/T0pLkaZi0brZROa5qS4o3qWdexjZqxQXZmbpQ2mTHxPd0j+5E7EMplNWOoXdEgxAfv3aGX9mk
FDBX4zcLa3FIWcqlqFab4Ej9XDNJFFlirJ58SoH97pmXe6QLOmIGoCXOoXPCYRSM1WPbGRBV2yxm
wSOTeQuS0JkQAx1moAixVmriiMk3zC0SPrXBAZb2wZ5Rrs9mcKbT/1+oE6732HOxjAj1dYV3Ag6V
be0f0636DGriHgaQH3NRvnByqpxGWFDh74VD87W/lee5wfjhKQpzk5iOJ99tpTRks6HsHs0ypgvx
wM6dAiGbbXMNXHq9SwA/CXVsf6ribZ00fN9/JbC9fEhTjBPyAr5T7Rildl1GqI++UAzGRqHGxfPu
UtaQ0XMB+bKvODWmftO5cDoQx+67c1amY4Xe2c0hsWCHi5AcJUAgk4pCbt3Uc9wxnXqdisMM+UBs
xpCUPfKfzd6EAUROVx1nYSjOe8SUpmUrezrci6oqW9NJT4ajI478jJa8wo1iyTtW7mkdzKl8e8SE
cQUXqiEPeiKu5fl+O93QQrmKsw9Csp5Lk0+gKOKyp/VxdTNS3/HXHNZXUBRBKixQrCFEa/QkI7is
wlYMRFe7WR5SX3L8s338s0b0mQzbVuIudm30uPrRfLq0v0mH/Y0lDM9XbmLBlkSVGzxCInMQo1IQ
FppVamo9oWi2Bo40lBoO5bzEozSG14iJhLoL0yp2wnyzS46AKegp/4QZUQBnritwO34yRmQB0dsm
+Eh2ecuEJxUVMFRT6DMDLwHytYJkBhfu2mpSwjYWWfWFiUuDrVETlyCPe2hyNDxgNxVMaaOLCew5
eLS3X0bM0jqhs7fojygGaIMeXlpMY9F93ZNqh/ZvocV/DJRcXIOu5VbVVrcHiZd7wTKQhz0ckWcs
QnLDYwTWCTUzbgwDpd2gm/80aTAbyKYC9lCoBK5d+VOSNIGOD7mvzoA2MjLoyfgbNC//zjc7r1A4
tIVGTlCtoetoPipQHrsA0wd+qOzfllDjGrg4udDX9UL/XrcgfABfkVYRgJIzSI2UXa8oGOVWjfoM
84hHgmmsliUInJewZpAQS2YjmSnI1YxO1HrhfJiQ0JaXfYpaKXk4gyegMd4tbdb0+2f5J4hXnjsi
yM0gtwK3p7THiyA8wi7XaKtG4y+rsZZbNhxn5wV+C8n7EkP2jMAAseqpI+Z7HACM5Z0PyAllHM12
mbge9RjMH055ZHBmtPiy9tkO+vyj2PEk0Zqd2z4gGgr9higbfDNzYKQuD+l5OhoVhMwR1FuISZlD
Txa0yeJGDv6cQ3IqTv+cmh0vUOMD3p0Il9s84BXy/Ma2MCmjTg8SFR60aGNH0WpVClPleZJRQJHP
w4L2s7bZGqLyYjX/B/1d9raRLuTMDQJ3oVbRpE56aWF9UmhfMKY0xawDtYCmNSeWeItZIFKUiO7K
Qni5AvxU5lDUnHoewN2QzhRlZRHsvZb1htsffYruptYbuTcBptBIQiJOJdM5LlNrPbW5wjX9NRd8
TrH7ttPNqyWIvJqEgYGeuKKJWAcYlv5IWa4lnVWTFAGGOLlEFW15DNhZc3VNGoi390xo9+jiJAuD
EDkGvqrTvkPaHhhsrwZlH1lVBxom/J4DzUux9NT5SUlCG/R6J0OfdGFXHQCZe6CiRI/5IFybqkiA
cA2d2ilxkpsnZLLB4ZZkv5Cxp3PpeNYKi8swcnK85avBvbF14oKcOxgQeqv/d4+XnKRNV3Bfm7FX
Mx8llWIoQvbJ454S+V+h6MwoVFfTOYB/EhYewptYQDsnPHcVQrHBkldp+xDdp7ikENQ9psxkX2Dy
Krt90e4XIP+LHqqCdBv216CRK76xMi0RAi/EkGxj4g+vFKcoGTzqIiNDMii/vO90qR/ARkUEogit
qbQnbSPNUwflVFZUyAmeBLKXIhr0jBVV7lYMcdgpc5oJAqbV52HcLiphbSECB8alMWuwgZPkbjAh
yF7FGVCTqanrpRFZe21nuPx3w5cAFU2Y6Vt7GhKEYv/B7DngjhDWAEdbtd/tp4UjAgOFNbESptoM
KNZBrYjyQKHRGoCygO8UiPjfIn7KlbSeHNvOUbqKYSE5XErPMFFRQCgfk5FpUEyHGrMMWX+wnA+h
5Qm3l8uILeaPIuyU7p19aevmF5rgm0D9AhD75EepoJWJFfjri8zKhsgoxvYDaWoFMKLBHyzcLHOB
KV0r1owVVpiVc6mC57o3DI3Lkw5FOqBiC7a03fXhK9/RnLc/Xd1Iq8+TpDC9S9t5d7Dkd+G8Nqrg
9LNyfoIuab9itoN+iAwSFt2f97IH4z/L2WyoGVitH4NKG3IZ0EbtvSCBPSCxZ1wbJP5thN+VjWpD
iuwLEbgVCY8bWyU1ECy78Kca/+trsw95Q3FxJIQOsSTBAUJ+FFT3GT6ZUiGfRq1eV/Jk8KwImPHB
vIa4099DFUFh0Gp68G5Zkf/N5QPI+cjATPp8mVPLk6kGxfB6vpdEFQgQBYpme+xjcBpFpiST+5ud
3/7X3naq/rbaCIXzkqv+o8XLkHANnLVTOQr9VpkqaZxcsrLRaBUyMgXJuNFi//iN3RVHKs1nnenQ
4LCeVtiZCFh6meVgyQ7zfG1m801msiR12WZeVJyqhE3mxe8DMXS7DWG20vbHJSU5pX6nS6XeOO7n
igEoSP+0LBUSiTo7KPIKMJUAHi41XuKT5qUpPoDJBKWkDqj30w/jCHQUSjAp8xU3iYHIEJWcGYrT
OLRKjgBYP41rGS88TksyXnqjSp2CJBMcFSAjUDFd0hsuGGl8bxes88ZWu9D67w+zojNYBzEhhADE
4X2PRrqrio+QZVq36waxW2eRQUgF9b+A0+xqfrA94qR6uKua9IwydDtJqBiR5R+KKbGfPKgs0Qgg
OkTzXkIedSALj9o8yiZ6kdXA2t3hUVLGR7nQLnoSiT0GuhQ6FK/aI0/sVY5t13aP1wEPQXkDhfvm
yGqZ1iea+mUbaJFohK80FffX1CZ76xalD8OfL5kDIkIhSeEzV8as/C9qyeVHoX8QLBZvXAvljKG4
6pJ2kGp9hN45Vsb5RPCy+Fmv1JsLFEqusK7ZSienKXp5xHuKemvcSBzfzLPtLsDF0GwVV21rPaIb
S1LoouZvADTFtL7qBTQ6I8oluMA/pMlyBfCOfIkfslsNXK6+0zIEoeL8APv9BtqD47YgWkMGjbck
wqGgASmWiyd/cF+azCZzHbM2o7NUvS2oXU6SV1kVKdl/7OyCfgcn4P6VUWIiF1o1VjSG/L9WE5Tt
9TS/z52bPOgSguveG4a19k9//6LUpA5t+v7A17SkBVa3mr9eOMIHB8V8jPg36Z8/wESe6hNvYD0U
kjAXz38Y+9B2jRCsAhHXqgPTer0cOD7DvZ1TZx8meW4+zX4JqgBVK2Sg7J3XrUqj7Yn301b1EEiv
u+DNpm6/czK+jT9eymE2PdOJW884K2/I/aoOnbYXBtSjiw/PXTsqKpI9eRMSRdvT86TF7uQDWXd7
nTyUb9155aP1nbS80TtoAIfkStub4vNxbd5yPiHD3NNZcutujO0tS5fX4M/AK3rKpsuzY5YBb8Qi
YDlyv1q8keRnuYalvN6m36LBrgWoAnwfB8ZY+t4FDPlFkfhjwlcN1wJ5U/bMtjLHBN+dV9xh6y3L
IKtHzEr9V086lv8t/csIfUKXoIQxXHnCspMpi5PSt3KH/3aXxWvzcXX7MnkxLfIgJu6rp4wxQHpf
wtmiQXAaXLWY/CuAp1suYC+9ja/cKM7kXi6fkI47NxUJgErUbU9CTgX+ArDFwOc1bPZ5SEe13bC1
2AHWFa729Iinir0PAlxQeKgM4u3Y8GInAEl53cT0xSo5EgC18fs6/si6M+ple1lNXFCJMtfaa5+G
Fg699trkViaN30NFX0MYHQWT/OkGxE/+qSTZ0H8M4IYz8iez95cCA1oERyGOyhJ+qeCFn1zx/YmN
vTASJXzKT2yA/Ih3kuAw5sIpxO3AlXdzDnW9+py3IGz366hJeqDIC/WJU2YNEgvOmSghRRcjAdC8
GpQf+EyqPZ5zJYmC4vV3NW0p37mobTvdnKgHOCaCmalgdlF3R56KxJWcvGhxegKxCHKF8AhDm81t
v6XoEjsp2dSsqq8uAYCzDcTViHoyi1ChIX9RLkHbuN+LL/QLfnjtJgQjfoju+xAbNB5HBh3+2iIE
RDvO3e4gOVIewDvl/4VRaWxi/IU4dZg4V5qLFhYll1oUB5hQVXR4uWMKaESBcJUpZsJ4wXco1H6d
d77Tqcu+CoXnzrhaosHHvuh+zuwrR3sDLGn1K1MoNY72kEc9YuoxNBNXGWyZfd5c+7KmqgJiRvtJ
4XT6qC1186vv8NnitpkKlCSNODZKuaiWxwFCcQkqC/Ul812hBKC9GIHVCnbPAiwbmrfiRPiCkfz6
TNHdeG58yGo2MAP/gXwMGyZq4EyZwu9Z1Ev7YaN46BDlT2MXPy+zdIZXKqfTxhQVoVf8pezpUpwz
Bc//gQyn/g7bYtlyNSHd6YVhx8qgvfAOL2D6tFwwzfLknDzupkUg3tF5fKKUlD1fN+oqBc7b6vPv
17mMUVpnqnv8Wp+PH9z/qaq2fPmSr26f80NpWmplryeem2iAUGtZk9CFAQRyy1TKxuVulCPLA6X5
SWyNjIHdZI1DRPa61zpkhdW/oqOFxYCPWKrdtK9dHEy493inBW3vWKqEkO9sNrQKBX/lgfxd6zTS
kcMnRNFmKmh0ZdAduf9OnhhehhvDTo9SZnVYlwy6IWYbaS29fyviUeJJhnEqpOMidzk/YtgErNMc
h3R9Hzgk27vLPJ2ngwQKenJoucAh0F+D/uLoyronHztvnlIkuMjeYhB2nLbsNTo6dYczeAFn76wb
65ItqmEZqSPAGgSQvlaR8lTQR+BZZ7eE8ne3iYHVgKuUz/xog0zpHtfwkRRnLOpTxreMWoGkv/U3
4rh77utVo2YL+TCNYrvOu3Co/OH4I7nl81EBH7vBl5E6mWF5sQAiuyV3kPurMJyMfVZR1lQHX8Mi
eyEnx3OIRCUiiyH6LyCJgoU2VNCXHDV93ZFN1nFT7/y/zY0HA0PoODtdZbZhJMwqNe1qkroAAslp
ATrtvcGiTZGMuH7Vcv2FCFWBl9Mh18PjdKDHeUTbDFijMR+cNZxoftvweZ5OinPuOuDQAJHxhpi9
8tZaasHIufdOl5OdRHt5hPlhf5P/J/QBDHn/RucaJM1G6rKe1pOY/AxOoFKDnMfQSOXyezdnk/oZ
hz7FOdf0Mpn7+/8r/sHbzedscE3BuIV6NUiGxbJ7MJtRAhnGXrijLHeava4jZM61K35ewPBqUiyD
AV6R/z4Hyx66+hVTO2cvbSfzIhbbbFPr7izH3Pq33hrx9dNvDWSP4xYFqHeSvdlJUhpK1P2FQ3+y
5WQeD3mcBOOZam4aDB63nT9W/THPb4yRnDW+LAh+P4hml23SPQm0Ym3DPbH8cAHATJQemINSqDYV
MNzac3cGIa2kuYeJzAdvum0FsPKEl79C7RHoLZvtQbCNR+Tk166q5rpX5w5Phwnf7dGVRCvK5Y5F
nHz00t399bAY1sbyMRMA83EUc7v6ZgeMC8sl10P+OH9+PdWOLaISl8X2mRVKPIexFtbc4lyO+i8q
x3c7npisQfR8ZezeopQ8h77VO2T3RqXkDlBV/6ULUHHgW41NHDz3kV/4B/tA02WArtf4JzPhfxn6
6gzIL5yMabJ+G1TXEKVhkuvsaqsldSvbclqwTGJwrzOAoBiFHWb78i4IkOl3pGrz2iFblqlpYccY
sCflgFeGBPTRRozz9xjPC+gT8FkQ+UpsGZvgEEalSY/3J1uUHeUq32+wIASv9e0P3GwRt11MAwKZ
3/jeh0Y2YfOTGQbylLIl9YkG5EsS3MAifjsUsJbWYN18tSxnwL1PP2fadOXhUwoFOk2m/I56wH1U
Loarm+KCezF/H1iKWKV51JJBBIwk9b4Nh1SqFl/drlWO/eKqaaaCWGNKwBgzUdVa9h0nJEndk5fA
21ZG+OmYtWnKy4feGCIqOl+3udu2N57VSUN9C6xp4M7VudjK1iC1f7j3Pw4avu46ENZREl2AcVoX
Bynr09kDXy8Y0eexPam53yELoVh4/3OmgyJyAaG0P6wNSY+MvRVSnssPPgP9cZ2Ce3XFz+ozX3FK
5z9DjZ64qK6OZn8ALAZWsxPNTNqcxhDCBe1NRPhEHuEJyd4ugV3qCSzN0yN3CUD4Q/gTb6Ze5C+E
5CMny+YWvNHHLLxdycCA0fwiKGp2RorQdYv0sEM3Y/GoYvo5yJABK1J4yO8AGwBoRlrWwl9CSs+4
l/HlUP4ChiV4oWxWr1JrSYHaMiMu7nbo3Cy5k5MRqE1PvhnjAUjXYDiU0i2QTLhIx0LSa4lAPtxb
qeyDMsh7yBuu2YHYQnsqslWH/pmIKSfRlhojE4WeOFxsSZKe7qz572+0dtqhey6r18d/xD7u7YvT
OPu/yjPxO45145RBdXfk+7/m7xkMA7pLE9DkZ0xK181f0jE3mi4iX6LI2NjwdYExBEP79t7eB8AY
xw3g4oRVCpTxoO5UxO6Xj8cA8n/TzaxlblKEov28zjatm3gFZk5AAuoCPNiEVbjEacVWHr6mTrf8
SLe30W9b7McF3hDO44Lp5CyQNcbd1pvzYxMKFPlbP9DI9x6At3ddvEvD07yrpsd3wxtrq2mkFtYf
cAcOBo+/Wd8Nnl3CkX51ny3cT2yfz7GpOJdsCHXbkH8b9x4BHqziSo9Aozy3iuUU7gLW/cpoufQ1
2xlCFdydcYwFNR42qIfLZPnrBD9EVzHEqWSrAQMlA+eAFmXIYGkZiPHWlVuRoW3s88XQ0th5KCJE
M+0PycpV2yKPnOiZzm5lm5338TvYBsSx1zSjcXxd7OxQQ2+u228desqICU6nAMSSTa59qSm52U30
7Dlz1jizG+kmg2Ava5jQ7S919F0Y27VHIyz6bxwp1CLjhla2wYU8OA8uZdh3uxWvBG7MXwEgpHRk
ep3AmA/nx3OHRzC5NGFZK8Ry3v9taDPjjKfKqQqHP7TwR1qgPsiEjmZiTsGux2aa/iAWqLlmNDKM
J7ID29BY74fqi+2NBxhvoE32vPZWgyo2Dc02wd8HIsY9pLyt82vW/BeozrODTtEhp8/ZavRLKKXo
L4UOjpRpx5+bBUdxroeVH8A5bf+xZYYruWntHEEJrgzYvQlM+ffoqoHsAonYn8rVyi2/s4ANpJai
SLAt87Wb9UkX/LolGEu6/4NfBJBp5nqiSJXjWnfGrbawRrl8a4zg8/EImma9XQderhQUeusMan8e
2FR0h6nMrkbE6nblynG8oLGNZe22vRHZT/9Jy88czy+oeKGSjlwon8JXAG47pNTFU2UUKeJOdHiR
tOr41NNIINQfgNfYlJ3sq80aD6OUb5iRe3ESZSypzEVBUCrt5d7K2ox5cx7u4J7LuTg5j4Rj4qLQ
Y+oP5S8KlS9JJ2diAt7KAzGhFKAJHMDkm2EVR/D8lHEqgWATaYxRRXQqj6d5MvJqOKA9sksv7t/3
EJaZITwtk4266UMvjedZ9vsjUMCty/6LEuWUABPIFXImzEy/Y8nIM55eIiDJ4tOCNM5NTr9nATFb
m9gewyQc+4iLBO3nZPk74PflZOn9sVNdD4ZG/pm9zZaaEnTBur4G4aYDWg84/yOFprBrJq87Fj/m
Fa09uoFZqJh49kUR7fVh/minGDcfNwFq0WMivg/BIg5QQGykb8KAzl+w172uFjQvzv4mIuLME2+g
6e5iNJqkAvLMOhxSW503Ozg8iskr2YwnBrKFTpKPptitKi9S45TcxQna2eHbpU6vdVjIwVH6qM41
x1YCBTPh0mcR/FHKaXpcoIBs9vNYrGJq2ms+6nzrl9mF5mSJTvR5thZwFxjuyQ+B7zVadx5DlafX
n/T7sXUmJuZzhQtIifRLFIQ2pFl9lfeMYHV2QwQSZDEb4AGAh3g5LysUxgXIONmZF89LHOs/SMPd
0L5emZkzueDE0p/8uECbjhHQsbQdiw4FkOqwvcnLD/jlY6oUSPg8yf4iNCgSJHRUQzAdaqZA0Vd/
JcfvZehl4Z8mJSFecrWnPecPPpOCRt2b+NFS+U/KmahQBaCWNJvp/ZvJX4JaRbZHWRdryOvPiH6U
iZFJETvxuMr/uGiD5zC1Ev2FsSelmuqPArMJJJQ4CFt/nz1+5lFmRH7QhDtIaoHFhbAigeB2NKPI
IriQupJXE1YSX79TbGSHqdO251uOaZziecfCfe+iJmy7kB2EwiopxEY+SpKH8R62G6TfbHYPePj1
kBFqEKvf+RjzDV7mIeWWYZZdtyMJzeE/KcDi+98s38Rz1HeWWEHYSNFTrriQOEnJ40jFoFIoGJ2E
RWhgj5/LoYXifZRWT1DVHWk3+l8EM+uSzhNeDPYwl+Oudfw/hG3hfCqD4e7WZ+6AOhYz0Av2GuRp
Ar6VS1WjY4JSclSLVN11N1MFGJMURYHWZJsEGcrDsOzu61n3E/NlSv+6pnXEJ2qQhAIgVbnL4HwN
fXN+M5cCvMRycEp7ormqhe5VE++gGddJ17155n2T5zzQ0FCWMToMFEe8QJNHubuqB+7oGxvtjXIL
Akcm+gUpIQtVjqO0YSHbU5JlbqhA7836PoJ6z6fYo+nB7HgaaoBA7WgBg16QuQWpaP9f4v7lfzfs
7a8TKnaUHPPcUXMilHXQl031QhkQL3kzAOSc9di6skkGFDKr2q8MaDQKWPQpTlZBzge4hFYxrPRH
PaDVH2Q9CkZ2fQytCwH80aQxmAIORpJ9AJ7v81MqykoYdyruMPdwj5ucne5JOc4TrqOD4MRnVQ8O
HNzKVVestG10ltEXsvevhhxchEGiBsawzhLgpzT9sWcBUjTITqUKMz4jmkxpZtwvRWk7RmnXiCbe
qdrNoJtnwYxQiVeF8SMp564ordhacRVFuw0mbPHSLhpHyZ6viiHn1EqDWpeO0pLmOQPgVm60bnBS
MV2HrW/aYc9nTVrm32bPZ44ogxGjMJoWFpWrtjD5gUAtZVVMJi1R7WbcOkXCPiFTTyaaWIO9I7tD
TqJ9sSzt95FqHRdWAw+bTs5AVIY526CivOywOwqbcL+abbR1i0mmdN7fpuFDv/kMf6rB7sgk4/B4
jEnMTyIeunpCMSOpLYjz9LCq+19L3GwHv8Td5jhYEffhJmzIJj0fQWgJOVDye5ld6OJTRp+tlYuD
9o2AvvH+YsaQOz5Gs72Dm/QPjPBLdW17IMYrf3Af2dPwPIHRPVT4ANxEVJu84RHcqtlr85aShpo6
NwyyFmIB82nVoNJNPVirkh+uuke7VhoUikyHyqD+32T/IqFvSHfcpSNnvbnuKdkZLULfbq/piUJh
fiS46h1iZDl0t7AhVm/IzAG1bgbOz+kGhywyIFhpFaXwnqf8e+zNkXEySrkkyNdnaxDJVCMmvo80
y0KMNeGFKeyF7wpmjPLh4ncS4KASlOcPQEITHBdRmQ0k94rwbeazaaUQlK8FWFaCpXSQlDAzA9jL
PHxvDzjlsz7+Hy3/fHPGrj3krXVYUEg9etWj/Nq/FiqMPzyiTLh2Cu4A7ZmrCZEYoCvtOXUupaXS
OBWfIBzLad9vvLg/sGwfvheWOg7YV10CvOh277S4lRH7p6sbcnGj675pj6h0bhGyoq9n38gSjm0Y
NVTmn3bSQAWZ8abm5Ri3M0WwUu8ZdGNvQ2oIJWxQGhIA+2cBqfAPc0LmbH1XyKW8J9/4CDR9QyI2
yPTtLCPAYunv+0mLmf8OLOPXnzsYrfxWdKuBpZ7CYxet8SlhnSonoTfOOPujA+XOy8Iw5eyyZ82U
zxvEwxvS7UgvD3f8g7vUIxuVVWoNl+kAVNEU2xoPWqjCTdewJZJOp9aBjtw2Ybl5zVVVh2/reB2a
+uSIdBY6aOegtWFojdHta/72OJNpOLoGHcAtncc73ao7+ufosTyK8GDcKj11kOEJDkxB2y7TTXZc
p+DTfpjvbL7Qoi0szqEwsVOy3gJDY1aKefFxmwQhuukcQBP5A7xXGEpfadEE5yYLnBqxRJJr0O4a
n9Oa+2P2ZaGjEZSiIuYGq+y3h6If6qZJs1oyz9jdTkjIAAYW/QBG6Gqz6EFd9VcgTauhX7ia7YOP
7sLfNltxdn33w47D0EEv14klIcrzGNV9kJd0irqlVIqcrZFWRta+mmt75i4uYjORly2NEb/3OdTP
24VcQiKGut0IqVtHXxRiWF/POSo1CZ5sncqcPXQk4IuGjtE4iBmzZULBw0UMGTkDrUhw640pCOJp
4Sw++um8wANZoYfXse9w/MHmpOW0vzmAWG1abH99/bNxEJ1RgJISIxEJyY9whsCrYsqKutAnB0SF
D2gAWxsCc+Jdw+91n5Pw5K72HtD5BXCHgdwwZJ+DaxCUX8U9Mx1IV4O9e0jM5DGP+dUvKSSAD0rm
Yx/emZ/N4XMy4sXSVZJI2M2UMXf/n5slIiQ9cU0OuRhkIV+KpffFA0M9VYbJ4vvjoBLn5ocDgLlC
Li0iEhFmCsnVK8U/i3CHfXazYP8DJkKqhH5INA3LKA6KoJoT2DiB5aO8WvJVZEKqKVuCotbHcAPO
Yn3yD4WKh+weGW/W0QUixfL7yj35K3d5y4l455sXifWbsYi6CCDID0M31MPtLz31DUOtE0CXFsXD
RsS0a8KoL/hyJJ8Xbjqp+/vr+ZCHwKsYM61pEcil28AjuJeWIBl7IzVMn6Jwl+MOOleZCy52/KPM
WE6lh1P2QmNbdmfZSzlGtbhwJy0nuBUrj/IEZxvFb4zxO+V2EDXCOfXY+tcpUJ7IzwSiipGnaXQN
LemEU5DvsF36PVNDY7m9YByUmsaionOoUMLneJTaZgQMv0MPj0dJYd6Vtztp3x3QtaHVlXW8EN4E
ZV8uJadXChAWMBrqofCVxjHN3LR70ZFW9JVErmbSy6G51+aiZlWsH9T++NOnKuJqPuzjZhdh6f6k
kr0CclqYIsKvf5/5zlYIrnNJcu/RNEttSNBMsxZbh+Ja57qyz9DW5FHsrkpSYK9J60cEp8tJwGmY
wF9p3hS2rGmj1bHJnopjqFNN6upYSMSP/Lp0rFiFo+dCrjeu+rSddI4a7t3d4PCaDUrUEHNRCjEy
53y6u9fLcnMt2dNUXwc1uqEKc4rEG+JIKjOiPAxuury8xUzhsEnGmhaEJLd1c4kApyg3KfkuSntQ
XnxJqqsl9opcteOjqQ7dw9Bzd0ToKAC6L9zXNb/fKGQH4UESMHHkOKy/LivDKY6bdDzqSXJUXsMw
w/+y3W6d98vPIp8grHoPTmDmBp1CtaxMrOBVEBmG7/RBLALmexbd7fEpTyLrzfLO5mE7Z6H+1Xwd
0FICodO3AuoNQdLhrz77bFXXqRFHuuLgxxEtyGLom26dW5q/7XKswRsQv+ORerOYuHAda3eBc7o/
+T+4Vhw2+5gAFgTwHmB89X513fTHs2Xp9OpxumKpoOCNzjLTcwwwESdVGaF47DPVzSPDqeqCa/JW
1FybiskanVScTQIDvs7IYbdKn4rL9Y7h/bY59mxYCuo4scIScbrrrGRI28CAqbSvM6Z51esO2pYY
Q5WWQqHlh3uhtrxVd/xG3h/A09To+MAH6SVqCKcGDFISxnUsLGp5/e8ZGt4p/QNIei9a7DX7rZpN
os0EBSbe8SntV5BN8EVYZpqnEztjyY0osj0/ycDeU7SxcJmkXnATo712/taCGrxZab7AlthMrVnY
IRo77hRAtTbKhqC/+KurTK1LnE+oAUzg16n8xNrfPziK9JExlM2VgZltlqGTaNZVCOSF9ewSGEfd
U54Myh0Hy+cYoxdiyh5SU58svCvbuvM8XbHmr6EKmf05+8VHIVhiJloESq2BLPaHG0qkcEvDvhQz
a0YzdcLd/TJrBqwVRcpPFSl8PVNr8afdLwK+t40wkHM9NAMKeMQ5hDeT/srpa+4tjyvcovtXKB72
xBX8FMpdz7YsAc0uZbIvgKOnfFCLxMinTyRJp8VRNtQpSzk5PThuDQAGwXfVoYO3Cdj3RkcnxOyL
LsjIsWXSttaDrPSAnZ2YLQsDrl6tRzy1edUBP6nGm9quhiF8b1zlbS8VwcyyhfVC5MrpO9av0VLZ
rINa7NCbGvubI2Joz7ktFfMc+gmcfDstBGPBBPQZmiHqwiTBv1lv6bkbP14Thc31plWIoHSZazaN
g4it/wiDD+4pV4Hj6tSWDDJlrMFE+h7JHQzE040q76X6J9VunEiD233AVEUUqWNIcaktVU27PXrA
sSi0mjCIcQzG6ypyp47OB226k1FjJN2+urBXWiMMeOfwT1iIyyJpxAdfR2RG4HRv5ny8MAAhAzw2
/d7Y50m5RXjA3mkhVd8WT9m4MGVxmqRtiiBUsGXVo19FMwP+d2iAfMVNYhAPt7KcCOc3gfbbb2dT
m4haPOyZMfv7Wj3ll/1897jP6qJnzQH3fPcV3WiYDgJBOWoaYX7yI7elcFLmilufNr3l0R7UQb7m
3h7pYiQSHI5EAi9kmiTfSUIKbwMe8RkHzBrn50khf/Mn+WITDSPvg1Z7PKj+x/WtrVQKglpOmuq5
Fdw/myA06L+eKBqNlArPkJhByY3d6zAtbLVXHZjwPIfSqOAAc/gvRCefdcnG3a6MnqwUpM9kLmlY
GgSHhas8uoMfiaPc5RBnKNn3GCtGZzQhF6ox3wP27//gjFzFXwdtRR4rqHM/H9LWEClMfKVPCbLH
snahepc7WTJpXWhlngxeXrKol99pAM4OnghJkiMkvUhBPkWsMBrgJ4UC23caXNdjydyDWW8Fwynu
0Fl2dxSnreaIJ3uR1GcfnDZleM1xVmO0jEHgxiXp5SC+4BGuZnVEi9nCvvTx2qBSUtAP8TcXZe87
kxtLNp3LsEqxm0jxct9gny+TEwXgHIRuwYKTzihZfk8vCvBqAXGqLT9PVn09ZZVxjVzQxkIXApjb
hK0XPkJOQLoPkPCQwq00DgBW/bAbmmud22SZ0L6rmLST8wZnjcfuSm+ieFTE2funhbTfdF6Y2Ee1
+bEX7CalV7O+8VrcNvH5OwD6/VhnCwuZhQCixp1Vk19nt4DYeg6FgBDHLjyNxcGqI7uohHWz+1NN
KCSjYDB5DQc8ZM3HhNQ3Gw5SV16gDYol0GclJ4KvJ+pD1fLLupaSexa3nlwhgQhswsEtJd6ANLeR
F7KEPW6P5dwVipyGK2+KqrjOka8vSooDzjQDqIKjzYcuykxel96Pp3R7Om9T+3xp07+xbBH3ONwM
db8qKDxIsYFa4IgKX+2MbQ9PhCT3aJAeQE0oSdAzsnHtwlU23g1Q9GO2jbyWgLQSP9pJk8O8lfGd
RAlJp53wqA7Lmq0QR4FZdCGqGJ6yZ0cfKfcq2IIOeHBXjFroptqEfbHgIVAWCz57qnw6dTXn9wL2
Z1dJg/NeVYTBEtTjLStdA6ouo3z7S5zavAWTIeSgf2IqBo0vkA+Ok3XhacTd2Faes8byjNTQo8HK
ffj9Fexf5mJk0NGqtwQz45RVbOZzOnhfObv7A/N0lKIGCeacq9GQUHP84M1o0d9yXgr558aXtrP9
yr1RUTUpflZFJvAUPGqOhHiURYEqYbh+h/Zk8gnuTfaa+i5ZLHSVWDFt5ow0IgGdLnn+/nWNhsAA
EldJg29Wv9q1O8mVinC2nZdLE8u+6CMo6RfVxKCcbq57nYmXFv0386cN84ZsUZaDfizQg5yUaL74
gEkdjlmGRG0VsI5OU55YH0kadqtOMzEAZbJr+2FiIqYFv3s6oRNhAcgkkerFgzXi4QaIOE37/nZD
UCMTz2VMJLLoMy7egb9He9s8v7PNM0Wtc6GLey52EbQ5Ddmo5Ivv1b5r5S+X+05DUFDD6kPZAz8h
LzENXimaNYF1TU/xMMAKCg5UL+/NcxqAcueOdCh7Of8v1N6O5Erf369l9goTQGUFNrpNH2QvfR/X
IPKo3p0moenX7VdopgzSI6dLdC10vdC4F3Ydh22zzk7Jvdu+nXbvtq99lPzigg8bv9IH9YB5bA/a
mHJ7uai5rqDxxcLQ5ObjEYbgwloe8Kq/tYw4mtJvR+dsr8oq/MY9ooCH04/YvC1V//fg4/CLgxE6
NXM2+R4Lgxgh9VzlPiGyDTi4Q7KmHa5u6DTvpGHkTCuMh+M1AEXMUFytQvf4yyyz4rtIUlPTOPv7
zxyKCzCocnEQ+qU1t8HYLhqyBby0eyn+D1G9z6rYyupRq+1QhzXjjvNdRXah65kfqPImzPbo8Y17
2nJglmZFEjOoHnjITIpXGS0O9ZxzAXTtm3RnXDWFd9piCOudQdJVkLeHCDvgmVPIKfBKcW3k3iCz
/HO0+dMsvtauldKj/PvJH5zh4RLmASU8WTxV9u+0GlHGvy224cKPk2GghM7Iwt+4ttzkdFFuS8Hu
dEnrHuNHG65mcu1IWtTVrm+LFwHvtQNACm8eRxQ65p+iIk2SRtrpEK1eg0BnXsUL5nEtuL3vcz2n
ZAyvQLg4vddg2eBIhAsK+WWmegQ3D9HsRRmcAEGdj91ADbfxT8s3aB7oDBKCYUbJd+3fPbxTXqLo
c8c7qc9ufbRXYnoCZTTcu20Fd6LP9Jcu/paBtkugUUy3PJHQ9KVtFRh3j8EXB8mXk1AfOfrqo3yy
zv6OiZSORKYPf57J4s5eS924OoWoS+sVKCEP8TXlHvijEGdXU56tahWGAvHf4mUoDRNUeWgPKrZF
w5Q6JAmeujRlpc9KUvplwUbbqOKDplfze4mfr1YES8mNc+5r9TSeewAClIxqF5CJv+i4McQlJ3CI
ySmv1fTf15pqh+FvShLH6sZ1SgP1JhotGnTiqIpwB5SuKOzgGkBJ88Lktj9LeWg3GlD6Wl9AO+hH
wq1HnAGAtWf7U0cRwNM+rKDLpfb0HGW88VVNBNyOFLW17Chp81XUNq3aZyNqYguE+m4q09e7gkgf
DMsju3aiUDKFgAPNXASqx42qlMC+VQmKAayYdJLFkjEkYZ9Vx3zx5gdNZBHNGgCIud+uLgSuSwz2
jlnf3rkWHh31RXuBwBahBVR/javjZxf2pWAqQdpzwTCUT86+K4LCW57gcnsvPvjXiH+qkkXi8rFd
1MblzwU0my6WX2t1pc8cMHotd/ef/cyNHTkOJx1iQqZ0HN2WYaIuIzflg0hA7HaPfM9S76luy2GL
i/pEccQZEEOr5nHahJxR4u2pCe3gy+j0POlGum0fO6FIBjdIxTW07A2uxKmJYeYsgyin3J+9WbQ+
l3QlxqccGlXR64uMDtE6+bRZO/mPF4xo379yfDo/lULERNkOBnJcuhJmSMzvnYSyd9VVtWatN5Zy
seQdKFeg48K1E1Bmwr44oHX1pFUsxThzsYLxY58SsQD5De1+p7v+AmhtC8y9DnqwtikTVU4ea//z
C1DNQB1rvcl2xnCHVLSN2anuv5/nczAnj+XaAr0gu0b/lxg9xI9/B7HDnckvfUVflCBsagHw8LoN
99ocOT6tVTlWc7MBUw2J3kVT7J/l+jTggZ3qMGmjm3hLRtPRS/Bb0waMiKEdndV1y/ciYm8YxavI
/+yS73uocDYJJ01ri+hefK52eUxq799q54K+xpdES0uAlrA01RTI8x7362aIlfcsGIP2tyZiGJhk
XhEcSii6nm4KN/Suau8bH57UDUARohuCt73RUpvtKuMORpLcQajWwGUnIhLQwi3DwKVz021u1mgW
qEMNTTxcxkeyhj5vp9VqQ33gjphwR1o5Lzetp3vr0NcjTvaUOAOchJdWQAW2+hS4YFCGMJ/z6WZ7
ZFS6d8U+KjedXwggAPI4I1WFTi4dwrD+GXZ4CC/vsqXO4ChAb0eiY+Zl+hfvEH9MqM2SrUd7TDrx
G6xkiYq1QgduqBbMSvrAYhkZN77cqMFBzpEaz+41JTziKu0leJsoJjz9328gIlqlkN0iZGhZfojV
iZlLTRnRkSoiyrV01daPcEVBshHnDUmPRlUINAxPAReO8y3XFE7npk4+wC1oOhvyvdXTlTTYMGqO
xoqATI2iiixUF5KTtNdgB0kNYBBDVaMP20/8zRoWYchs8WUkRmcbC+4IjWcR1vbeIp3ZszvGCjqq
ANSpwlVwrmkirWfcGfg++0FAW/bqMr3S8QgBiMa75oRVt7DZoCl7Qoi799BSO7PvQodT4PjEC/o5
ny/8AM60ynTM253XyiPhj+MgZ49HsI3AL2If6gSrgtRyM6uca0lUzTir+cVisoO3EFCP0a6mtSaX
u1TnjSalugbFfoayedcRVkQZ+odS9UFDvBFmOy3juVphMZEoPfSe2RC7G958SPg+6UsPBWZTU8LT
u7yrZhLtGFaaTZlgEoEx77BA1c0w+IMh0N7pT7KHaR+GF0Hvn1P6AApLTE97ue7AMbT/uULFAg9d
uGR73NKNSqQ6U1Bs4rd9oHvz2+I3TZc3QF3Yd+W/iAcRiOYXj7Deyvey/TBx9Q+Gtxtfr4z2Xlbg
lUCuw4W7cz23It0KummbqvjRLibvSQjYRtbdVNhfTEe3s52A7ja9koUbUdf0EfuNHdxYvR12pOQ/
v92+E4IJO34b9A1mC0RvTdv4pb+vAbtY0d/85nWoIsuX5/i8lxyBK1tXmYxZIODZp0f3Em074srU
lBOyD6/FpevpxhsW5P3qwIHViShcY8JoyQ6Hq5+fVV6IRQt08HjG4AEixjqrh/U04UlGCU7xmiRW
H3sVKezJYgm6RSnj51TnAbFrgjxaE1TGEWNZjbGpCXQx7paOZLZzbPjCsSU+kC57ROVI4Yl8MHUu
v5TsCr2clb/wOf+2ceW0awZPs8aeHScX5N0cyV6okxu39e4oko4ft8nhv44Khpv7GmmsYtjrNBaO
5CyN9CpurYnr6kNcOZI5r5wiIxsx7dYLL4VFjYCeVIqT4jL5382xTzpz1xMB+KXsWR5umKHZdOjq
tzvikr0aDq9dNyQrcA2LAw3+lGd2xjxYoE2V3t/nGDURs6V3eB4l58zGCNcT7qFqeaSscSpqClIm
dMp6h1QtBxeKGTxHP3ICSu0EpLQ/NokXHXJxqOSq/PGHWqbIrdXUqcc6kJwDUk8BBjVMAbzhl14d
N1RRdxcWDtlqE48JSrmMK9xLKIrx35KX4grX2vhpOWYsQp8Y9TrdJbIvmn/eAf90IltjSwQKFpLH
qwmMUM8W1J6sQ5b9WA2fhIrJAqYq5KqlOQdKZzyBYA/ZPit9rYG2Zra8LmefVUfiFH970A7FwS3F
Gwn1vQiz974CnJ28uX5lsu9NR0S9WrFLhdiRh2JrBBAYLCKbw9Zr1hZB30GHOI8MUrzQlJwWKpG+
GvxD4/z0BfsbL9PH1tUHHT2E/1ZyKr5YzoYuF0AMmEzsxkvkhrRQ37z6nDTBgeGkbUCbVSXGiyGx
lAyRlqNll8HuldesGbdm5nh49/Vlm4V4hCVBKlDP0px7rNeIgAS/uTpAzwWIUnFE3S0xUKzF7hg4
P5duMEnL4HQVk37v8PoHk0dvg7LB32TneyEdASPWkA/2/bpHB9B4yxA1CycChFAMxuyZJcXTiPAM
flyFFxXx0tYiN++A/K1DWPNDkFNl/KOP6bwAWt0ESYkv+WyGRsJ4drvrjO9zVQ3U5P9DEjW9JElm
Q4Dj0NHerXuncwH6TECxpYWPbaKX+x5mLIrcFI7GGfVeKDdZ2oEW30d+x5yGVJErsMkhR53i6Oge
hJ30hPgPKkmbPXx7CzVAlzs9k05+lkjsUkYVw8V1LeYOP5GHeBEQfyiSVynzCywzG65BFV2ww6tn
uOXSK8ib3oxsrVM5cyYfsntRLpWOB/G1VjqxzLVi//jVP7xqeAjf5dOD64tdTWzvoBR45WdHHMMO
CebTDgfmrRgVyMRtA3/BmogsooE07nuCTlaYehcULfNtRJJx/ynkjjnG/U2U5mflooy63lLZTD8/
bKwvOdf7+VkcEnA2Bk/+OzPSumx7JNQSU0XTHAT3Zq/pgHW0HOLYk8+i+uDh+tsU7Ns1Nmz+izXl
B/RXpy4dWy+FGNGd8Mb1pgn2SzLFWwvNABRupzGAsKEC5bNBn5jpiGVfqBRIYTXNtZjwJOwsvTWr
MPFYrV26RjpXs5NZ1+7UjU+OWMuq4nKFZuYd/681VIpmLaBNmnBPYCyEfT5tEeW8PJ9cYUO8f1rB
9YQgvxYCRktrhTNtzUVA8X2GLu3zL6Udlyy1o0BREZbNrSZ2vH03Ax+LawU3JmRndEjFvxFs7UVN
xIV6+aHGXQxp26rBks+7F9p7tCxJG6R3bK45uJ6qN0Kjadiob/rFY2Oj1gryRkZPoBGlcUXH+orp
mQH/gNS9xJVJHr4YaSmEilbakGZDpxGcyxVEx7z2GU6/JY1s9H1IgegDwLm7XP3RkYlwmM9J04Jr
MPCQYfrEa9GCMCa7K0Ja/j/0+/LWf7++ALUK4zOJUHx/b6O36wwwF3wwg4wPNlaPjv2468QXmeYU
RhgJRyd/EwkBlQ+iyyg9bsBYzBBQuv3+7bUEPoqdKnNSXzOhj70psDa7rriESeHIFWq6higDyn5t
o04gWecWuhIdRg4iTdd0m13p9/kf8XIi2y7e0I2N7lKhm4SoBfAAwHJxhuZh1rXQZRwiJ2HFA6Kg
jbkLCTFuiZqyF3CoLH1hQVurH3XbMzixPf1OUhagCLG02bRRfOkLKXJb9HKtBwzM2zNxltKWloFC
S88ah4qXJ4H4AlX2jG6NDBKjAsc7RV08tn6kjtlyIEKoGx4cGqNlJ0zA8qaEhKaOlwzGESEwTCUx
9wDTruKauHElfKe6CtKBhKXSXEe5GTEWj25ydQQlfDbNg3N3xwRH071fBXv8HwaJ869Zlc5zHJBK
QPktCnpgq6c6RfYKNY0BPjvwQI6JGCAyoeMXLnrJDqtuWhFsZxmPfQEomm1HpGWtpHdJ+O5uIPVJ
WhEx9jlSx37DVDKDLXJ/WEYxvrqYvRxzR7mPL8LZB8wN3t9WZTZQGQW+THVg+Mh6YlWmNJKQjndF
ZMEfCwjLE04xnDvFtCkotgK3LI43ZHQ6DKBHjgCGgx3q+paB36k1On75lR072OZt7kt7JSrzvLzH
o0bm0335aAyhA8atpXn6MUGbeBSH7izhBEkj6zfqxY1ItEtX8FQAdHMu11LBgEOreWeFcosh+Gjk
qUjMw6TzjSiZSlaTTGMlWJLy9PXD3SDHXPdFFMuictrFbQ6eJxHrq0J1ZZo7bCi+h7J0/UU+b1C0
xTp/n1V8wEFcQlYGRZD2w0G82gXgQT7618zauo/X0tfIgzi8YaSmA6SR8n54pcUiBz4vZ0ZwYUlU
X/uACEKGNWTyDZbRlPOnFWf6tvApP6cmSzgDukt8tHdXnRKwcWKAx65N2YEGBqX3tzKQ/rm3ptbQ
r7Bn/DJwbqT5PH+EvF4vZDeACY9Sp+76ccPFCmcUv8c65w2LFpHEB1hOLWRs+84UsR/rv3SFLrB1
TFe9H6oID5suoRYac782HTB1qUSqqavRy9ms0sYktHErEHKU3DsQf3s0ne5FrgZc4pvN50eNvMpX
rrXzZ0F5q3+0XOiwyTBEir55SF6RJDyllj1zPQQZ1ZQug7oS5FC+EjMJiRrA3MbydKRSSNHvAtuU
GFm9+vmoJoxgJgbyQ4cp5VBXfInAtf4XjZfrlQ33NAUv3S+P1p4gaSuHEYFU27bT8SqgpSb/WeHp
ffy63DHV3x6FKbxrQsnDiVEo8oh85USYHBNleefgexg1ZYmfW9oPUhCwKDIr3PcAfRrfbZqVCvVe
keoV+MJG/IjWoZCqGTVmj/cpW20DIO00HLpC2/b7x0dLutgezClk8fT5mqR0MPjFi4EG1os5u2+3
qJFY5sfN4pUT1eSAcFotQPJ3KEP/GsdVLmLu3CAphIB6BJtstPIpXzd+MwkLlKcvhH/3aUDRAOhN
gfng2XBooZBKh9j7c551ChCAdTKxI4V40+j3Y2hSUUU+xMXRVUUfEjtEpq5qc+/GhQJS64baksBe
t+9yVhwIBYL8RhCk3MZuC2qYhMJGu3EsXed7/jYqq4+nT7pcCeioNvils+5DwrDi9Gb0owsOR6Xj
69M8kGQOy/IrcyJYUJw4aKgmYo28ZYZBmp6w2ncqNocZvL/vsQ9fC8/+5YOH04/vGLUrY3ks4v+a
aXik4x9VCaMpJvwGgLGuCpDBvcxxbQaMpiujWX/Cf2gJ4mls4c6Q1Apd0et8uuga2dw2jjQhVCrn
AEdsbP0l+oJ8Jl5PuLO627AIuijaSO0mwaHchYepBZ2a8RFb0LABHlTCFXnQid8R3x1Jf07yO107
05cIsxPXCUc/yTGUfqkuQOso+rjR9Hw1y9aiqFHZ25DB0ZnoMr58zw2X8qULqqpMF6zAtIv4qiHR
lHKsxMvtAL/Y+BMijH4qEqUJcNFmicwNKPLqN1/tSip4MVCUSlAqtfRJ45KOd2QZT6A+65DKaMJG
tpiP+2UmLuLjsdi2y9l2LelZCXEmoofA1bwXdaj67IVMFK4IuXj2vz8r+kU0sPg14qKeWsWnCwKs
FP97PsXXNRzauLxTu6AfXFURD8cypMXIkMrHbx+FvmBTRH433I3sSFGI9NjLhhZllcSoR+/J9USv
oQmwHRmd+oucdD6vJyRs5cwR/kf7zy6XUyIRL2DW0YyyYhNn+jvnNc1heP3V3tVOb5n5uYK9p79X
9sZ45Xo1Tg1xPEPdUBqgi51mohzYJ0Hgp2uiWm9zSWy4mMDmBsUoL57I7Tfbb8KQibo1A06B1886
XStYP51YJAjd8ebpJZfTcvrWVNe4qvOuzJjtuzhwCdB+BQdIRl6GczD9QYbbK90sZYMMI2pEXv3+
34sLsMGFrmD2jShS7PXr+5U1GWHlfMeVZX8jvnhodQqQZ0zXHfp58Cuab6et6Feta1mABD/J2mK/
+JqwoJ4K+unHskm7aAvF1AdYUOMlXqbSvR96+l8WEpfoomQqZxTQ//zuXXGtlJ9PmSymCdGcMziS
NbkvZo8MWmKeWuuotblbV5t8OhLwpJY45WA7GJG5d+MWXFMEaKZl8eBmx8knSwAIQTS3FtwRGwIO
W0bHtEDvx8gyP9U6/jZaj20v8uVhCo7iHtQOG1v2SzK6NDmJ1u3pPXUcIV5xP1bTkdioyaUXwcGE
RVqo94dU+P8Rc7oFgQeUiU57ckWEnJ64a9cqQKJPSii6l22wNTVXgVGNJEIbTY6FY9iapk+rrFG/
JA5rZbxj7CMpTiFPQ/V9gTJ/f8Pq6iZPmuuTw8MKDq2wtb1/PQ4/FtBbiMPtpXAkuGJHh/RmkIpS
HB3IBN+heoZdat9bdpAXOYxNpwtdPEtkwXDCvGOKx0AamwSX0lUsqbrjjLz8+ZKKCcQ2NBMIehth
2aDsupYmJP0Jszu0avRhsbG8xX7Uq2PK4UHJ+2wge+T0jdgYfE6NB2fZXiujdlqkyNETkGEtb1wo
XI99w7wjFrtPOZHQt+36nhEYMeRh+7jdcvfRhpxvNEl8X4rGH7ikh0VtvWcNCG7aDakd5rg/zeXO
0M8pVOmQ3RVoCSWslhOQ5qFRSCP82MbSx+Y5+vXyzhrwwh4HY2j8NBYDueTnHFe3s65ngRMGTyIv
h87gzeGLUURma+7XQOnQSPWV16memia6sy+BiuywFyKgSSvck1ArNP+krdO+xYhiuNl+02Nlwv6a
qOG/ZiiTM2GXJrP9NDO/Tqz+A1mKepThUd45LJziJKn5LU6Ty/up3ZAL5XsTSOPbkKjIQJ+BKC2z
DVFXbj4CyDmh24R+qTwc0Hl/tQ2JybviWAcg5sjkwHY4vn4dhv6z5QwG3cUDynKDhI4/Dv7Ikiua
7eiO5dX7QbLR5UlevpM3dmGBBI54u+zd+M+EPM7x7gNCFr0rHFC5AL3+rVWvp9Nl8s5hnFrNbnb2
/DXTCXMv3HJCTytAaapkiMdlJJwc+vUAC7vGcqDUtRlK7fMjbpY5Aw0UOsc6WZ5IdM14la0B0dEp
IP9UDHCJaD6A0nZlIPW+IAJIVKbBb/6tl6Hja3tMdM7DMZxdbXiOiQMgHJrsoQg7zRwD6f87lmhm
y4SvOEhWkDxF8MmnK0y8bOfiNxCkKRqFuHkee0V8prnYA+vw2CNxoOgKKYeHiG303G3ZvFnFDvi1
YC0svjxtvwXh6UwjTyMcEYPSP0cp89pDfgj5LxT1EYcRpWCtgRomGQ1w9mfmnrs7+g0S4gyWjmtp
ParFu7+dzrQjU/qujyE4C46OEcBJ3F6MmtoEB+fiepWU2LGn03vzFMcgs/6z7gHKCJg9CpOPgKck
1LdVDyDStC36etWudJVF5S34w2IdOxBuPVRcrJC0fzWT899ow1eRRiLNYnR0uBJ3CopNOCSYnTev
49JLgKDsEF2FKgN3Al3yM9qFIHrdGQ8nvKKJ3wF9HpKR0DQvG4QDUZ/W51vo3daKIL+lo04jTF2T
H3BC6E2mwy7fcU1hakNcmXOrgbwowcuHTcBgCrvjIYwo1/sZC2ntP+CAvq5le7ABRyyrJQHETWTi
ZBVJaql9j1wYH2d7RiaWCiyTQe5n2Vw+RGoCPaHtlqO4WRNUezdmYnAQ2TPpWnFMJZaQAcm0UmIR
4Gg3qxdnKLA5Vsa7hpP7nKgrgAKmvVoGIRU31eyBMkXvP1RjF1egFYVxVRhTKZInYJzS+kJ7IHs5
fr+1WF8FKhJZb5BzK0g7Fr77baGR5vpGzvAu8gKIzxHvkRBuMnp0IWgQWHp+JwnetDjMHzmYOQ7E
v+aZZTm5mqjXcctOi3rR2844IXtYASiuVAxJmnwLtqpqsiGGLmGEVss6Jw929EaNZa1Zxe2+oRbg
T+SIMNeLYu7aS8Zhsx+07RxYIpQ9n/fmqdBx3apQbhAqXJ2Aq3wOYU0R72gYvxPT3/YL+LZDPZo2
9jcdNzklppRjAr2G2JUcZvGcLd1Xt7ltvf+1ScakSnSiho09RC4r18GHf5jIIwTLhkbc9XXDzGdC
svWLEK6gH/ip78zCoMyV/u0CMtGX1fNi0oFrJhHkeUx5SeA/KwGFcPPdFfQnWkryrpYRaiWrOKGz
EHj1BasdU87+ymmHoCYqHFRcnyGrNrVuGRMhWepPG805t5h/dPfVRQdgzp081zfppSSI216oCPjZ
R2+D4zFV5vQJZ4TxAlPGRaJP1upBkhejspW1kE+pLSaQvUtD73r8393gwqz9ltsJc9SrUh536xhV
HzYmWQxKMtW7gdqDD2JeTqxa7HeyqXls0ntooodVzG3NcWKZdnByOCVNyEsZgq3orpfnt5yPOQQq
sBWLR743LJMuCO7LFSEvTAyz09feflzeLncGGTwETQ1AkQau4Y13v5pN8bR9qp/1iCX+DDxEtSDg
4mAIHxvAtGMA0vfeDw5FtLGiTVCFHQO8U3bPu5d5ffIkcj2y8OWlN22kpTTfZql+M2XiiQG+ub/c
4bBMyiJktVpCDxEoYti8r7dAhveNDu1ioUFbQEZzdGro+UBIMxyYWZFD+cmiH+wu+b2mbR3txnyk
sJuYX1X2gXFIUXSugva2GGVnuNn8IppiUgiveSE7yN7Ztd1nVuoY2i9u8iZJDsHIwg7Eb0EpgMYI
eRYemUldmnNcsa/U0b1FkYLzCb8T6Pz5a8asQfZVSdI9zLvC2Kizjm4v86wi5cfuzv/VWDYWVeFc
zih8aB44xukheK/GXWqm9mbWtCDem2/FDvytFTS8I4Gr9DFno8E+ABfV3XgzSoqqtAI5P+vHxt5J
IgUzHfFuVmP0vX1uEocR5Lq41wnkEvFzO78snrl8OCzKlkDn7Tpmdj3r6VxRQr/LLfhJGMFF3LT+
kBK576fyKgQAd9VIqCzBR+eJLdTg6lqaCTGTD40y6a7keUFII7I/NhWJoc5if+ar0QesneLzblrS
hyjMkiUZjop0KHFx32xzcJ/OoJnDG1fAHDM2xQXZndUCudX28aYD23IS8scxeT2Ob60ZSgYPX61s
UW8H4F5NOdXS6NguPYshhYxAQGLW7t0Oqsuqrft1leMaVfmRqj0o0/dbPnANp+sBoEF9zDSh7E3/
WEGIEX07EOlxoPVj+ym6yZO3FCow27SaP/TfERPefregiY2vVXW9ff7JJd/pvgfpCUU0rT5pGP8C
JYgbm8BgPTkpRrA6XlmR2OaJxU6EMoM8DggF5dbpcdWYr3N5LvfG79syiNfh/EcGHpEtNTSMKMjq
LiiYoC8683DG5ofRRy01pJY0Wf/bucJOedf51+X7Xzr3BXKQh2txKmjAPaTeevdLnENpyoZTDPZk
PGfd1vZV6uSCfzyyIQeRM22oom4WomFVY6WUbQtUPV7jLGTy9c9d1si41572vL7YHeSapWILR8W0
AkBqJ9i/LoP/PFMaYo8AErE5CrizEXvbdOzDfQD6BoTojCm7DrrHrUmZTW/3CG9Ue5P1tKPszvZ+
CS/sGpejkqUbgrqPv4GTUq5yDYjtGY/y0+FBn9slmkJ6ratVFmAl8+J5LZyWEwdwFefmvCK2hnaQ
gzVU6k8Z5QZ/kIZu1Nz3O2RdrdIUYij9iqObqSai5Vmgbfu2A0vbXjllmG2g8Omale/Uahv7B/vf
LLwOvU8EkPj6rJmilLjaSkdhq0huo+brqWOpACYFHwfVREX5VXDkzkYn2mDXuJIFA0ch3AOIPx5j
OpXZu5/En19UK05ZpQs30rlElZRIUWFP9nBiRuFf7jipP94Zl+nnz1gO+nXUr20AKengyF+qvJ7J
KQrvZqxuTmgLUDcokEzVWoJ8JqhtIAOrJqjFRgcK/YO5qdLdAvaJYebeeLl1sllnfPf2l7NFHMZS
n2F36oRcRjbcdcddkZJam6aEofH39TXsoZite78x/uDV03k0hYF6diB7qIO24d03NKmlKBFiHVU+
r8PiIBMdtItiVN45m0TBzpjicr5Ab3GOFMlJP7Ob470ajOgufVm1q6evPVa7fFKO5V5B2igLLu7n
TxbSDcMDdyOMUyzCqWgDUcxLcX3MJepZ1IyGn3vV7Yry4aDY6if0xuqmOUcnALWEJXDtFWm58Ohx
Qm8qwI1UgWI2apMhUQ/GnbqrevlzMQQn96Ix1+mGjGxAR4VdkcVSKSsI6Z1qwpYRVygAgjOI2xy+
3MsFv0j1k+fJE6Tf/5XD/F9jBwVfFc87gOciodzs6HElIlKNauhS4IQXrwQUMIT1EHFn+ILeOMX0
vxsheqAdvxeMha9gRhWsT3Qy9ENnVsU88QitHsC5WhWuSjn/jz3XKBsnierP7NYHYdDS3Jvxyui2
zzrL4QVRWPODaPwJhIrw5nNBNE2yD96nZpVsJO2hvyqCGMRe9mWcmtl4e2zvZctPACXBR7VlRT+F
jTXhpg05P2t4CspEctyrjRW/pdX/j9WhfAhGzIMZ71XM/kfxmjoAQoixnCjUlkLY7q8X2cmTvLHY
30c9s8/Ogv4otuhC0vk8xl6K4s0NnFZV7JYfjOJ486qszy0GhBkP4lajqwOcvTcVQUfCp7bco5AI
Y9x2+F0CzxshiJsPTXjT1W9GaXkoC4IQeihqnS6H5tHgA7v+QLOoizGghw1Wp89KCySbt2MkY5M+
kl5IFK58WkR6PJxkaFJWsO5ErSRmOOHfL9tY6XwLopyAS4nKnG6Es+gVShR/7GMaDWmggUpMPyUI
9PH/FjnE8HLRaxxmOcpbpe/3+jvwCixbmajt2qnapWghwa8/y/u4WWmMBMgdWQqzGFJLKkWc3nO3
yW52NN2DyscY10CAmGDZxK6omSJ1YoEI8Wk8kzqJKZTWZMTXmDQLilZsViyy6O4Y0tZmCK6vIH5P
s8grjKsRTegqwRPRn4P1H/Loak3PH4q3yqVtW6UYbkUHPgfOK9jkapZGuvGKwLLSYFlj50OiTVxV
DSAxtsMCSZDkC8SBzTUlJwoCk7JLiJUkGh1Ac8nS/V4YUw5Uk1gXsRaqZZjXsQ5ae32RGCPupv17
tMdDZ6hQFWBpi/466s7y5/bjmf5U61ts7ZXp1iy6Qa7VNMQrT/CrcYnUSUHbvMvZnVcdvK8QGzHc
jBmdLE0sz6KMzidaNKpJJmtsTB+RvYsUIaZbWmWMKXAc93SH8PBB3TqHRsKBbSxH5E22/6EfPezY
BzsRX7nTEnoRyQ+4/Rn/qhyPbw9DhsN6uV/0GLXFVJZH4PGh7dwyLm1M1nTtzsKihd/xAcQr/DN8
GXiEVsU2yf3WQ8jQC9YLUEhsamrVm0ELj0rVGwOc+FAZQNMY68+6cQI5wvUqrUXAJQDr+Kk5Q7pB
nqge5O5DBihoyfTO3gV2hyTjFEhv8NaQ2+HgZlTLCIwG9hI5x3FePmzhsozjZwCqVUKpwDk0mFHh
AbTPB7/OYEwKEZGLZd/ds70ioLTbz3mnSNXQKR2R9hWp8UsoA/p2A7slGzEQhUQZ9YB+oBKUHf7G
DESTrRapzkeBxxkr63gJG0Ij9ELX1V3bwdzzOpOHnOaHF0twfYAAivwqeUW7ZLcg7nJqRBo3CV/5
wvEKatUmCKiJVf3ibPAR16EVg5TMdS+qP8gSGcqTzFb6EmyFBtk6ZMkV0hxVTtrEGoYuzpzOXV8K
8mACZ1SymfnsbNkqvFcgX4iAGd+8NvJI0Huk8H9XTUYqcSPpkFnji4UwhNsheKYC6hck+5VXKjGe
95zuC4QWdrk3/bg0lnDFInos4nvAlI7hlbkH2c8RSM9Kg4HVash32fHyqTu305tI5I9kCY6MtU5D
GlqI4W1BwTzPrJpGW1H4OySVi2LaEeNC7SJcjrOQfww0X3dXN2m9shLRLDTBsn43maixxuOQb3PP
EoopZVlm2Ax8L7hIpo7qefhImjWdP1iHoTFhldTiXSXq6uO6d4bEV/+bGxw8yU38EJnqu/RXeoQk
gjKMz1dBt9MgOZvorC6xE6USJHj7xe3quKcqqm2rxp0z2zgBC9/BO/HzlUb06/X6x3dQD8kTu+li
XPVNUFHYdL76MbKtvGXTbAq+ETSCAF2RrJVH3AYSQXkE6veNvx/0t76Cu8DhmKgvLKOxcfPmJg4t
6R43BeSWuiuelzSGb378lddUcuOmGXmNk861dKpd18FNQxZ4krXiv0TI6y0CpFtLaOtgCqmnfJgA
JvJHjEZP8BG50EVsvIKGmVfV/Z3CEUtp59Nu/unrpVclq/Q7uUW9LY6LaTMhjPInQxDHMLg0VMM9
sf8xEm3nJhshxb3vOuqiMwqfs85RoZypEdFr3EruOkyjXoItAGyZqMeq82npZtxn9quMLpPSJWGV
Dfn/vJz7yCBIVyU51v/sQLA01nl4X7C7j0SfU59EwdpqdD3VHrncf/VONw7I9SQEkMZF/yjOC6Jx
vM4Rle3BF8lyKHW+q7YfqvOZ6ukc6bEcDx9ldaAllc5iFP8YBup7TlFLlh/G9HS1x18vvdyJiWj0
qWSk69WwmYpKvmse39YxuUjDsqejUm6Lm5voDE2y6Ii/mkD/3haKuiTrbABomiiGXd+V2M1zLOck
5UPenqvmlusaHst5UHsFrVLLKmr58SG+vmkNkQyNCFzur0G4kWoUmH6YHW22tSRhIHo+8guuXIz/
1E/yMhqNm7iOSv92e5MWm0d8XkhLJQS8TCiH/PkCxEsYAJM0bgjcvql7p3N3aOJahkIaZg7RjOVx
ymGEUb6Y+ZvTLsGORK3OFZ62FI97cgg1Jgza1FUveE671MdOccfj2kYQ/ycOI8YgOuMeFIHU5d/Y
kTO+opXHPHmVjmlmKQrmeMXbcKDIiPtZUQH4J5X1ol6UVPFfjpKUHr9ebLQBT7iT5PQf1S55mK2z
s++WSEDtGLzLbdNek20EO6cL97RrGB42zOOQKjBoWvY7PX0SV4EmizFJsGfcFNdJYHVmN0uF7cGa
TEOUC2PJWwJU2RAfRxGP8VSxrd6sS028aD2ak5dPFD0M3fCuYueMxg4sLoQ5bvtNcD36BSUOr/pY
MMy/j4PvvwEK2YO/w6J4iZECtk1HtY65R1EMfLFEqzCoQ/IlrIkj9S2J0WUNHXhLCQV4fXkJtyuS
K67KYUQrYdWqu6AOcWUsDUXSdEYlx6WIji9c/z5ocdaH//P/hbdBizbpmJFDm/AzeFL123beaTy9
AKQiOWiLSXtdhFz8e6sml6Op4NkHnNIZRzIqGqphIsV24W/iYjPU7G+a/5nJCTdEwn7Ei94kAT44
B1ox0rhVPs0VTdZ7KDicg9ONb7nRAFQDYj299RefMdjkJgOk4GMhUMgdo5oRiLx30Xhuf4ec0m30
FhHTuQPBCaXVx1Y+sZy556cmlqBsYkC1sLs/41PUo49FEWz/RTpeI/rPITaGNTv4qorzWiVrJyNk
axoSDCevEjsC//RIEqJiL0tJn4cmOR+YG+bGtYOqQx91R2edabzXZeueywVYWsf2FcZq2kfTbYhx
fLTeOS8GxJtZ3HTD9Jd1H6Dt2KSte6iQBHTAT9aJuw1vTA3RJ0mlyBA3GdOzTiSfUicOZDlToamH
Gb9m2PawdFtKaAw+7w3Mi12jzFUulzGpkGZio67/+9AQPrabUajx62shtJjYeqfCb0J2CP1ILC/I
wBZduRNY3kCmv09EcJ16hCf9C28I9hc1DDoR3x1ORS+79NdUiB/T8or+noj/8YPUbchX2uBzC/Gr
rvittQmZ4uw/TnHdeAl2H5X2CQ/Ie87jbvjZSOQjCu42yIfuZPCKPDbEjjM1zWk0l6AUZ2qDvGSo
/O302o51Em0xkFeESM1P1fnFmkkL9COPYfqM9jrXs0Fa2wBHJFuvDaRl/Ss9siTcdlIxgWr8uMOn
+NUVdw1WC3HccSijFwgs/u5Y452rAlBewHgA0yAHXcrr1QMtvAGyYpYJTVQIrfHpsy3/qgvmF/ma
96aR0Mr/+zuj54a252YVtzxC6WEttrGwO1e6NU1MdP7PsdxfyDM2h0w9zRvNwkiClnzueFwJezJe
FpzZM9fhsnVZMYfsnV53D9TagbgGKq5Ar5rsMu9PfnDyn25UapG9Fow9iH4149ozWL6wxaIC5OtE
qZq6FZ8xG7e7/nr+pGeMJpeVxBFUMepnsNI2Xv9MSCJM9hyqGWhbQCp6c8fYpAVLX6XTSyWrB20r
XpQfJObF+2pWjZ2akwe6iKU/XwzlOBxCLhrJTOzFva7dziqYQJuoJeLv0Dmn3HkrE8caA6zPvnXi
V6mXuayIXHfSfhInMDQPc9fGwaI3xWJLTYtwFurxw1IV68OLtk1pvSFeAV4HPQzZZCXHrnWz+Rg6
vVp9FzFwbLENVD07RXA4eXJy7MCr+lwZdTj6HVPjZmg2RxCTnDqhcaUIBqpFhDWlJFLniywq1qOD
X5Ew+0OUbxZPtvQeKNuspcYGDBPXcG7jky59di0ap5YYlYSmr7CL0QOrLx/E6GeBJXE7eCOdgJQg
m3Z+9IxlWM6jn4hArDafrvYzwz19EN6spRKGpQw8ncH/B6cICMHtrGGBW/qJTRGtMNuMbcIH5SAd
VAnGdc9mJVbE+zF3qficGyN3BzKEBJSS93yD4T1w4oq0f7o33KlymlLFwrDXjiUrkfjOugrdLoWs
er4VCqdX+Eurj9Jvu5WlBmeHwHICP8fHQPQvGuiHeOxpISYrTihDARq6Zci6PzzhqYKqS/cICYnk
wK6OOVmtkXM5ASwNupzCOvnBFJVvLRJGbXdJ2T3lKTGsA+Z6+c1tkxYOkHU5/+nVkHbA5I5kctQP
WuPo+YJQvjMvTuGiWclwjOfrilbCpkK/iZKd7dlUDYWyzL+hDDXALhfc6TjwUIqoSCo4SL/lTfBQ
NJ/gJedYl11VrkgHTSRWBR1VdDs9+J42ieeQkEff1br4JfniVQv3it18YlQDMwKsJ/jGz1l3oYsE
5GY+gdcpOLT3Nd6sqXEQhgi1OfBYhoVLqh61rZUuTz+XCBYcptuPsar1lersT9LIZN8YHULRc7MW
IFL939tgorJlad8uz0JQ2l+YY2K2PTuux0yN+gV/5MLRqR7NAW+I7c5ENkq/QY4of4WQ63Idhb+Z
TbAWLJILBqpMuoL/NL9ItAe/Gxm9z5xcoO9p2xx3qpXN5kz1+QkTWuAm15CKGRLFEp8qo2QJqQqa
PchCPsRitnZSC9kOq0JlJtfojcRqm/IDiX+T+kyft+rg/ubQsLEAxNU4KkYRPkH/0hr3RzOC/gBx
3rTDdvOGSP7x7q9ve5lJdQaFGmAeI4L5z5G/lUSO86jDcaucJM22XoFHz+du1vvJJOpszYymmMAY
OYlAYskGL2QQbXGK//3uW2ZjE0IfsgW+z1zB62L3tt4gM1l7DgqPNDGLj7Hq+ErIPEkNJre1eF42
paFkT5HLJwq+jwhEgzGSBhDKtuAk/7e1PfJ+W5w7S298NLaenbUzkA6Ho52qeOpknHyTnNPgCtmb
cEq6u9PtzqaI3IWXRxaFnhG90akGqhF3v9FTUOQtnVH/m69Y4vKi2RyfBNaUJf/nLxd96Bp7u9wj
se/kD3n7UIbdD9cnEbnGvXJbhIHq0bvb4gc4U47/3thkdJhsg8V8GCf4QrsfIXcUh2vcZsmo53G/
N5tlN6hDpANOPMopedUFGnL/RjnMFe4QB9K8hq6VgXsbRmyNjYAfRYF6N4ZgnuOTtQJ+8RywMU4j
P7AZ2XlTc5tfDBZhcWNX5HfCfu0ZcjR7zOS2V+rkzr+q9E5yDBfNN2gnT82B1uMjt6uzNK65AJBW
5Ovzls9bkkQiZKdojmq9Ljkno0zuOYptFxr35bxpOTuyxGi1i+IzjQiTX27HHblJAOeJ+JZaigde
gq8NNkRuOJRpDIvGGizE0aNvCigjvdj5X3vH1kx8I6Bt7uat/sfR/jOle/eUEaF0PMLZ6wPSevjL
rLS4S5UmITCCOiVYTXZ1GJvygjlXY5CW1NMSXN+2WaBfp6tJej4ZpEhd3iBlWr6wQKgOVNW6JsPS
3EK9GRqV5tLnKbtq3pBCnlorYRIGMfPUsmLjYvNzPFKQrD+g8hivZt2dmAsU/fFdloFxnYa1rntW
Dotap2ZngZBnAnN9nc3N/pbIcUtFVXpU3oBYGfea69Z4J8L1EMq+B1mbIgNdKqdt83bIE4TMZlbi
szU1TOAfGRFFp4qOa1BxnnKGgiuE8rB2pNQP/rgobgQ0cQTQSW1K4TsgiFGcRJRmF7RIip9o+KIY
FF5vGM+oZjB05VuKizF4R07cDjTN7/ejESbAVhG4sCctDKW1S57yl2kTU643R2VDRkibJMANt7go
BZTcHEfF0zP+xuR5Z/QLcZDMXTOoUPgqd3ik3D80ImPT6ZW0KjC2RBqLAtp+JgfAO8uBlLTx/INg
rGXuB/yQRuGoyvhFZkZMKLi9CszBQjgscRcFLopsBmB/B4O8gbGrf6/erIfewttoA0IRZNTueY5g
t510+Az4gjxLn/74c+qQRwzVNtnhLHRTpvp79wl30QDiiZA+eWs8AiCx3vzteZvOVIjZsXfMWNPH
G/aVIoQIv79x1FzfglrzU0qtmOkpClprGpu+2g9BznYcxO1RC4BenUNv4y/3kiLbpPLWoBdzbENx
kF3Fwth6QkSFXnQV3TFxZjzpTsTw91kXXgcXGiHtQmFYguJf8Doun5YbRbvclU5VnIilBElx5aHE
4KlpCOMQevrne+kQPJyEj6QRHok3RJlzkzfKqfYpW7qAZdslQqhA2NoCve6ekkSvg0uZED5AzT7p
rwKN2AZjj28TXzqh1OM98dijEiRXAXEWjMfp5amK01kqjgNoHWHn68tNNP6d9yGthm9zLgnWliBs
m/jMdObfq+MjIArQSJ04uSgzDRSj0URwmic8u3Nbc+7/YfbfqBQEk8RMi+t89eVzHQxF8MGLSYZ7
Bqna3tO0iUY34eiUNLB/5BOm3QtyfN/ijmUbmfiN8vFREZo46EwXJYdHvwxyBX3e+PxNQeEZs6wP
y7raPGF1QMSxzFhWsNlcMHdIuEUOzWF4orOeqVDeJU+3mgO9kT061RttjYcAZFp2za8nZMfFz7+t
7ze2YJF/3e9IpcNzqFHIzAfDsjqLPc5/NFHA738m9cN08Yq7BMDI/raaOR+WwrnidjJADqGGFlMj
YtpiVmxHiQhXAODPFzRPiXI7ucmo8rezGskEfZNc1GKRQnQP2z7RTnzyza56qcDZ7L8DK80GLvYb
5DLGHLiXAS6kbxP0nt1eICfCEQe5CoduLprbU01F+mO/AMqf1AQfPzA+hl3Z3OMbEcmyQOSIj0Oa
CgqCqcuKCBYVVDue7iTJ6lwZyD1LzFvBcQNBOGII1272ESmK5/YS1+31tyljujqp1RrbED6MwEEw
NZfAfPOJ17xDBhxkoRrycnM6DxUU6H7kx6AWcz0l1cJIjBnzwR/89UyX8xGIiVPTwEpbN6evjzqa
oCUNc7HShMiLwcqK0G6TZD+yn824yr0OGdzZ//d+j4bm8BOm7maWhgwsPkE4s5roxnkWwgUxcZIe
CNk0RreAR6py7l0goYU0LMrlfpIhL5Lf/4tRjCwBU/1dDMqODrf45SJwSpDjc9j/bphMdW4h95c9
ytxejgEgGBLkJ1Y8UTVb7gLoYQ+tdjZjWDZZSP1Y4OKcoT4Eikeof+wUS8rxfn5cHX8wBxsH6fis
XBV7r5/UmeUlbv5ffUGP8XWeDI9FLH1uBpAoHGZak6w6Bf7bI4J6ICNY1fB5VhNfxc0n1QvbP/KV
Te1btO913UB5yRG8l80oefcUtbjt/4cAO6tefXDP7SiL+WXUP7Gkjo/3Y4WmFbmAsX0sL9ZlP7BR
tEjpD5ENcczTK+BObhft4lFPjSwoltU6eNj3F6i6i3aoGJHxB3Kx1nRqcec2xiqRQkjGz8QiiMKB
jE5oVRwc/GyEGiK5R78qqPQWpLo2j0OzMmawaUSHrvXzG4Q41MaRlp8d0LtmbIWtQu0L1zuN89tl
YNvaKXrDOD22X8HVTqesi2JdA/TyQk7CJfbL09HSyhwjVZMIeV91YNq5zHoi36sGJTN47vxz7rMT
P7QGunNQ32RxUAbEkr41+03cJXQ/OsJDAR5bFv6PNRoIv0llkfoQB3WIUoiN2Fa987VioamreRoi
3L5rE3HaanqqZ3wfMTZWwH8N2/aaQar3aLqu3gcGRKhlk6663tPBLEShm1F1l6h68RTdvI09VHxE
z3F3T/ayLQDFG9zKTwfNMo/PIlnZLYNbTB1lIeAbxlUc5uAWnnic9EzKx+9+4KCZoG4EbTs6ec4Z
TfA4xa2LBPvhsx7MMoJ7jfx3uTpDF6T/qb8yA0Ymo+p6AccmPG83p5htHn74+jXKthvC16h95C6Q
moc4fn7vjUAZpOnncvmxMPw6FeKF3sWgU5sHSz6mLCHMhemBDdjPsypyyoQrzZ4ETOlhHYQyJANo
sBgt6ADajYiMwunbMQ8PIaPZPsmpu2ENkYh6k900O/EBh6X63Hh56cpG+EKqXKGGrFAaxlVRYjdx
Bc6mFJbLzYuNeTBVoUacxdJRfZOyYVzrXgqbCG/UBksBOhau4YwOx1vgtzWvgm7wOSEYleHDl47V
SeJiLPwZ6Z1Wt9czD1VaCxfHIKQ4tedq11ELm0AUOeCV4LEEzCopDnA4PxrGwj4gB6EId+OS7KGh
ikkme5DrtEr8JEWbrJy0RfXkXtp5/4eRS9rtzrF1W3PYHz8p7J8Max2u3BgXttufkELIKV90nduV
8b2EDa0gCe7U2hqYt233Fl6Fk07SYe7zSKbNhoUyp5ZYslcyKvEvo/aGsLzBcfp7e+xAxWfAHzqd
x7Xj61Tb1IiXxqp5PF63Uwdr3PPjDv2/J/S3N8VCC9SAzi35N8bCctPWUh6ZpuhQT7jauhjYtxM0
ldsO/LB2l+FTzq9g6ic8HIUZ7lXlqDdSya9dHufGdZjdooF+gskQ6I23HZmu1qrt3g46wwxCsC0i
2jRs1dy51jRYNMXQlwx+fsqJHsZSTdIkuCXxWIkSbzrhfGeTeCePDBy4jkqKT54FxMjvvHw2FT6c
sZ0X4lhVDByNE1bLipmUE7z15n7QKDXSgQcZfpNNHbMjXHeAjih/PjZidGc85kkG++8qPSJV0UJn
+lm8bbQwUDIwuuR/FRuyYGOjF7fFut3x/E2wDHZL8TDhGsqSIkxhUFX+G9vJYSasRQyJuATODnvr
3PD+N4oWKpYYY9zsho3VP97vz32ztI6OB2i4DrTFbytCogn8WT7ZVWA9nrGEhiqxDiFSR7R6+0ON
8XDT3wRjq15RvOUlUiPvvSxWEwYqh445u6V/E7qojNR21rgYGeer8gBG+TI3h0YJpheYkbuFELnI
nwiE+zT//0CiYE+8Y+q4M+F9xv2IqMJH4Yn8eyeJVJj3VFP3P77Kswk9hCm19eOewvlPTHzjs6cW
x+l3bc+10yFz9yvpzcUYIAR3UkIa9WDQX31bGk64zmkzKiFuyN+x0MKY5QcfMzC9Pj294pYr4Cdu
NTSXLz3TixOMtiM2t8I8Zx6FKjyLAH27cqRvvV04tZCqVyJnwz/u7GA/NbXK13foLLEs7QqnnDlN
K7wbB4yMtcvyuPYFMPB5nJNaWZoFCSqjO3yiCEygizkV9N2Pv7NuGC5NVcqs8U0lo4XrCP/DTkYk
XzBHyOX3/F54SRH+zbPwTaQjQcHFLngqFH6CLSUop4/lKnNwuK1u/QdSJkQ34puzWMPtWpJXI6Fb
liD1ySDiXF/qaVWLYziv1wGYt+KLFk6xklvFPyp2cw+7lJNTPXbYyaHEIe4/V5BY7ujUq3RweOqw
Pn/vB+uSjioeyBWm/mz9ohn0ILeL63y7+YnoILEw6AuKyyRSQ6w2k4t3I5adgCFpHMErqihR6qfh
B7vpOkDGG96alzg2dk9TcFIn6eKXXwaTbKPnvtVepuwjqGSKNthlgIfPrXqJu7R4yoldsndS1AFd
GsMS+nEpOMH/TDbd6on3flUgQgH/zxa873j42fTb5hqPxMLlMmy/mbfbmmr10p+iVuiMQBGzOyxZ
erKVt8Rd5L7jD+yUWaqOR/JtgwgUxoR0u4Bdw+sUp1LeSp/cimaDVjv4CJvafHsBjQ3vI83TpI+T
ciiZGr1hKWvKTnFdH0iVFD5dTeQtVJ5FI5HkRcqbC4r48Ec0fPJiuc6mciFeV/q9Wmljv2ZKxdqj
ybQ0NHxpRwsUF4sOw507/8xgCGP6PkGyV9dsQAiLEKYTLRP69DK8gTVoE+N+fJ1Lpnl956jkran5
2xFsNzFCZ4WroL/N/cB7H3qtrwEDN5k0S2nyy4ms+Q5H84X4be9ucp9bCpDMPdfBiOBseR/+kk6h
i02sjGbrJ3iX0RimKj3SWhs4pYr2uadTCoHJrLIg9CXxfvWC7fZJ/xczQ/ualLC1P/BEKPxiI1Fl
szMH1pI4V2G+Iuxjs0H2YpCLuBviKlqWcf577NElurJ1vgNlcUH6/FWNaYl8mw37NveD/H67p37b
PPI13BsxiQOXhYUaH6k3hLaLtpIcBw4gMZlVZwQYJBccjt0dRNpII3tPvvrww0upxrkEmW7BH4sx
BbsN8C8gKndN228AXv7E3ckMcJ7Vx85Xfj1DpB16WZuq1fGkrGS+m8r0lfg8xCgMUPidq5fbt8ij
QV3NZNs8DtZKqghh6g3vVuakRvKmpGbddtJVihmXv5OWNSqltozfS1u0vFmdGfyUBRnTmgM2jC6k
mIUlg3cUNw/vslUYmiNK8V9rACys0NQj5UDDPtdaNwVWk3X23pIuXiEOHbDYgod2MUdhpiYI8F5D
efRLCG525Qoosexk7cHRkRtVE4qM1r8m1eZtBx1eXZbxccMcMh6cD3crcNy03dkRFBuHDmHe9Uec
7JNbMz6XUH9V74gnzKlYf6+t4B6+yomRxxsQhPfPWMhnpvEDZH2DBimRuBAsAZlzO9w7NSpiOnT9
q3i9kaJKra+I8bLqFKEl4wIONiKG4gE7QA/FOmhA0xN1fUr/NJyDnyMx4yhUS69My/PE/6hr9PXT
1Mis+fnDkdc0V3k6T5X1Qhuk3wgF/2irkxkz1rFklCw0Eh39sicMpCl055iCkTLsmeL94lBUW9JH
CbXD5iE0DwOo+PJL6GfiJUzTwNpFEzoIK12vNyOQTuklnKuegvWEyKPaEs/PVddYY67JTXxH8QoB
0FI1lCTF9WmDAaYkKHNc3jh0cjPk7zpE9njEPQBBrcnxl9CA+2BGJFY0OyklWILG0c3YRGnsCdHB
sgV4+shXBVhL4giielRsQg0eQTXiUd+QrUkB5gpPe07K8gb2suBtzbI0Mu1jBd2eAOGyHx2eQNCQ
l1tk+tbiZA6uxZPOtdwXGMWxGIFAUPvWbXGOdPKDUshLSIpTDDdbEbSVr0UCqL8VaWVwr1vZl791
vBsHvKbvA6+cK5re3y6hXAEjb1/Hw6Yz70Olx/K8BfGCkIA5iQ7MwhDfj9hFPqnik0Bb+JBkGQqQ
RotxetnPCHew2Tqo94rmvwBPcYF8o0k+uLMg7vy3WksTrB6enLUEtNu0dy9DOFn7+6DJqT6LcSJV
Xbj6RxBj7I56L/TOyO7UV0E458SsR7JpFxp3r+EFdBz4LQARN21DOmqgTzkIC6W0Yb9AwP6xrjKH
SA9FpYTuikYxLTWB87ZTAMwjp3On/1GqPErfZwyt0rmTi8ppNFlsJmjwjjYPp7fxUyLqVyuU18yi
i+AX0vEa4a69ZbJwyOivAA8J6MXjUDmM6miC5eXXSQsPcw0KAnV2p3xicCO0tG71orKHtjrC0wDZ
q44rV46hxRYsfdRvgisZ2A0sanbiC19BF5XbW/cLU9xcguKP4S69pRLHE5cD4/uIC1p6bFVzw9/p
m0RguEuJNF5qBhMR//QIjEMOGi9Y+6EuzwVk8vIcpCLmFFThoERe7+ezChaFL7oj/doiwM4C5Pw0
tC67b0bKIH8n8eNCjgJZabZoqQUp3PnF/YjP7D+Vi8rES8VIO3nLhMTHkKsbbV2U7wo+sH/tbP8n
356o8oPxHWxCrX6924pZ21DHwO+PLE1UrY871rALoBd5+vwwCEuzmM2R2p5+lB5jfFKH81YVwLXa
pXp4BXAEF0KIIpP/thz0duOjkJVJAeS012ZCDfhTg71f1iP1/AACgGNOjxtNxVc59ji21eQsr1Nv
+cNglEsJ/dCG9sNeFa+/JUns9ZbCir0VS6Pbt5AyNomkz11/5qcje5ipjojaDn3z2O3uoUxmLiE7
dPP1+Roqc17UqihOJbUhdikE9FgV6qKaCwZ3YiFihTivDsNAgCus88YaG7BE2cdsFFQjenmeK3uQ
gn2ycI72FH0VXD7mpm5JC7PTfAZ8Dwk20QlOFBtVv/S+IwC1z6mD8O5FRo5cazdXAYiFBY+zI2jx
d2crbfT2HymWXZpCaYHdvBVRKBuEyYZUiBLPpK3XfeG00riE/RLQI6bs0FXi/AOz3pOSs09iJW+q
eLPJ5lGnicEP6wniegArbQA1aa3n9InjJG0mbsNsg8BBklsKVGK9BRdEyBbwGj+0cYkXs3jIntBi
OVAbNMy9k2s4Hmg2vwxGY054ZIY7EVrjn7smue8f7wIAintqRPtNKwbUVrrs/wCM86fp/qDvproA
jOiL175bBVhUv9wlk1b1EVLhfBJP433XAa3eqlETlfDo2KfSdqrLxppaybjoxYDC7Mm4+FlqpaRR
SV9FQh2jCLxMqcdXvnituqQazwboU4/Lt72T8yPZYnotPfGwsm//jm4Ss7nW2/GOLmFJT5bMHAFA
qG3ZmCiuoMUG3Y2ZLEvM9VeT2Jm2BrUjyBCCk9zcWf9b4wHmI8uXS4Y1pz25OdXW9zdZHxinXczf
0l6zSWEqemnOquNXkGgt9ICO2oEnLJbD52g0WO9EeSIKfAXvc8k7FN26BkVNFPKpUxeBYCd3LZ24
DstSrFdteQ3ZESyGfefMyUJw6qvWYoT3+ZmToqr2d7A19k8TwnPYxvtdQksXDEyzKYwndNLHe//E
iGde3GLt1wm8TW6zTf+4Zq6AbzFedzUv2DqBBKLbpWrkNrMRKH3yx/trlbTcNx4u/vvXXa4fsi4Q
xCUDwTlmtrwj6gfS4caKWmPoMj5P6CgDAkkU06rjA9aiPB1yfq3XXeUzYc+I4XdtqCeo9u3gmIIQ
ALxUfzYtPVqr84v0bzBtyAEmqrt0GaMSANbCAaT+d2dM+7Lx2WwprXpv8/inxsN32OfMRAVq3azU
yubITOVdCvwHoP8ZHqbscrS7nkuYyeSJDxX04K62dQ1fXlvMhHnZdMTsXleh03hCG3DxIFlfMSqK
WgWJPNs4EDyZCNAM1WaAFpdy6467RJtRAwcGPkzLkg4wHWvw9OEs8CbK2ET0W9BiovHSa/nNP67x
vDU4T9ifXEjjyRoiShVlWDNm/dY+HOOJtZun7WxYpYSb7pfs9UAiz6Xs6p4uDVgh/yE6IKj7XUUC
4m1LeM62nYYKh+PV+claIY6Z7ru9q6TJf5esNKuHeDJEBT+pD2JHpLNCfvnaTwL+WDeEkU5QcBRA
HmVhxliY5TTqAvJXWHS8D1iAEaL+/OBQKC6fvXLKPsd5YmiH7CsFFR03xbazkex30ucMpvepLXOe
XiOLzjVCQsWSVqCj6v/mnY49GoDbORKFJujaJPSGAMDgFjEicfiSGJHOFJpgIfUqONgqzuAA8e1A
vjZsI58lTgeBJpLLK08GNvUcWJGU+Qws008RcC+BAbalzAn5lXdnIPMBfoGmBQfySuwaKfVVnlt9
nOac/ZDty6rLvXDntJjnZGHhFvGI8GcIUrL1wxbZ+t7i9JIMtbBmf2AWk5B8/Oj1tZ0AUA0KGHfn
MQ0u8vuWGvUCtU6+3uY+KJCVEoD/zihRpQHiW5gf/nWPILPlDEYOg2YwaCpTxtMMKxVwn/CNhYtX
aX+nrC+amTAbuqqlRLjd6YRwW4LUizFqXiLlotjnhPp6Rt3iN2T/UUaZunxn1RQhn67QuwzWj2EJ
cJPxjB97g9J+v9jGuP3DTi4em1i9+Be8Ik5PMAv42ILBB4eF1ojM+4C2nwSdOWhS6lq5itUdwUyB
HxdS2Rxpgn++ivxed6BYoYlvH7G/M2nLGXjl8//0LVmqkxhq3UnGL4NZh/Yk9h0+mEc/RR8uVg6g
SBFfocl5wVXf0gvlun78xeLh2Ju3Row7FYL31KH2orusNLX85D2GGY2fORqR0Y2k0e2PkMg3RMti
fdJhptFScAEv+5AS/QkcCA2lkeVNufeihP/5FHuJ/QYt6pSKXrPoUQ3RS1K7pL21TKGlOXsucEz0
aU+7lUFn+OwllhxQ1aYHEbgmA8gHbwu7wxrFK4EUT1QXfSJhuquMUppP7qBrLq06lmXzlEf3u4OR
acTYZGXOAMUlegvCPh4iY7g3YbPbSvBQ+F0ItoyB4e+aIFuOqYe7NLjl9r1UG5ht4YFygmq+rT+V
mOSRJrDAFbs8nnVfmJNA205JZtstpg5foZA4T80uGUMupMzln7HaNzeW40AG7wPFxWNYWCkrBNYF
GuoiFk9bhb+W2+AoayY4kCtERB6wV23nLCaUbbvHnNNxKbZbzLBL+kRnWZlNSQ7JVNTAzGD7oqvY
EkiLCFVVfraZfhsYG0SHD9PQYnxhZEjM+DtOL63goo5Ry8zHXwZC33qgj3EOMYRCaOJ6pttk9Cc+
8yL3vkA1fIwrvWXn392vCSBNVOJb1dFSSyMM7ajMoHa7j+SoCxUjDgcWr2+URA168m9TJ7Xg+foc
11jLs4B7HU2RtwF99yEZ3CIpDSNx8gQ3rSjpGOf1y5qeVrcq71a4Bo94svyaEybfGEtBPNH8+hPg
Nxv1cRQtCywz3nK9LLWogt+vI5C8B9nBUYrueUoigxN4+3LkY8HIkXKXAZC/umUJmvYzmpIzLoKY
9nHt9MtiV1tr6hGxgMHAUSNcAbs64EL1SK79ce6iqG3Zl/WU0SZf1/elo1KQaT3R/RRjc1vejiLv
/CQ9gtRJxqc1MPQNp21Z3CFR8yWaQAhObC9eGQY9ZzQGdZ9YeL+NCjpCJs7yTDBygMpFB/x4EfvH
EDYp33RXh1/Lc9hfONkvi6J62cwqB0x9u4oc6r3FQec5SHBpe5LRls0gvzsnx2p/zqLQRRF5Z77f
LuGFIEJyYoAUMdlD3jUmW/enpyFrSiuWXWNGp7gz7tsXCIL7iYrVfTcBo5WzoeKc58nvNpN4MoHy
WLtyZBXTWnL72rRyrlV5ejX2xcC8NUU3HutoIrlq2Ap2gDNIHQ2xMZETCsjqzoXWEGfzO8aR2EDZ
bpdw6Hm+cLsLbYViSZ5r4ByTzMVuQGjk868VAo6/8y5vluhTUq5jfQW4Gt7CBO3o/JzW+rHrnZZw
nIv79eqWfsnKOT2KullgBQq7C0zYOgdWeU1ZMfxld8VZIZvwXhWNwm3HMl+1xMiLLoJ3A2GzEGGR
ld1lfLRJN7efolHH0RGlDAW8EotyOPj3MC+otuwtF5Our7/QPV6T3p/9O/qI19C33/FOs8IAdB1D
OlNPr2C4slTrQEbJuKMvX2ysIahb+KRmVnqEUFi0Hv5QuGALX8ZrdbZO6RlZfi/EOvP5DAwHrYyu
QgjIaxSz/84vkzVl+0aAytfUxaA5kHTo5l6FgasoQEYS1EZBsMeftFzvg00U04/bAf0t8zaVYTTa
Evo+dPg1x5fBjRqzouHIr5FcyD2ltFrwhEWHo3a4TaA9hSVXNlZdp21sg7poyzG+T/mh1+i6l1QX
PSXWT7uy1Xw8aT+DD8gmBgyzFV0PILpmpQ1AIaiYD31wd7S16xsWbChnFNdpNkZ9+WiziOnAnJym
1jyOfo5DiBviqv1hVwx1viaBjwlri20Vs1IGiSh1N7Z4HhoVWyblCVUGlUanR14zok6q+X/AdVpT
2aY5CBmPU+UnAygXx1+Ef2ON4sjAixZXz95mcrTaiWnKEkXVPFeYEAWHj/KLfNvefUjc403N9DGc
r+7nTMKUdfCJoEG9KHwEIRVsw/xE7Il/siS//i0LVV48gFoXWIw/SMi+swlj2MdC9oB+n6vCBQNe
7orroxVJV0xHZk52TMM6z2QRdmQRphZ/BdRNpV+v0dTgA3atEfRjvvPldOphfRRjxgAC80lAUrDa
yp8xrOgRGbB3ViZE2BOpp9u3RU2LBljpc/h8gLC0HLi6ENW3oU4WM1QouRsB7MxSMV8UTKrDXW0h
956JTy+TY2jFGyJZ3vqKNH5Xm6Ebyt0L1vT1E5dBYRLePF3OF9gUBgWEBXpuE99nrkL1CZqsznv+
UWoHHOuaZ+XuXFfs/p8/z4IXSg255k9Gb4M1CJRxcbaZyuDrSPDECi7ak4SDBfpu3Q8T0Fa/Fvm9
n5p21S6Vt5k2jmErcTgtq+I45FVxZ7kxPlKxyQ6uJwX5o7M7cWHw1pFlcLGNM3RqDDqGS7LykjcK
pnZ8zERPICNIphY7KRuUl6MkKtzurhCcgbPUzz9YTYk3KA4Cln1+MBhy6RH6LozIRaPnscr48vPh
ueupHyhT8NXtPvcJhRhySoXPDlENbREGq7d+9uvwZXko3nengXXsk/+9XqZK9cDopEGqHDQajvSF
AwPl8+kBKtCosIjkUeLKr/b//7LgUSVwKnzU/jxHBlCHDP4P9Av74rg2qsBKz4bCOcU5lZPUUDeg
V1VOBkAjBxOh18nq9khYuAqdF0LLY0y9UT8/v4N4iX4LfSia9GMc8LEINC2AeVPUeW+x3nnidQt7
t4mC71Rg/lj4tkpdGF5O93D5TIkSaGukwW7DddP0QMB+KPM87QPrr5cFM3CIAM8IJp7v7vV4zESd
JVYspHHbcjetlf3YM9LGv2lOz8yK+XAxqbFg5c6v2UdOLqaK8K6noXCXXLG9YbBdUTLWqSL/k7IL
wo6sxREJ6pRqbkXvfyOVm+pp8S8VGxtqGzfOuvod3xUVbvFU6WLmu9uhIf8Pp0eawXkjE1y+zaUb
U79ePQTfdU3JmAcqWvC8BJh4i/7KTOvUX2VVmlSqBiBjgxlqCz/UIa4YitR5g8V1HzEFUxe0VdLK
y6PwlGRm2wNC5x77UOzs/5a895Elsji0VBN9J6xG/jWN5kXyJUy+BzovZruOWx/iNYu0Xe2ZOgS/
lJddSUFWvvJtfdrCWkOr6LRFuP4gWFZ+ThCRZtabvpaYttEZlZKzolYDgfAnaVVB3atMTbvGm+rr
r/JiAXmAvmMo7DMyfR5w+0ofjddYmi/YeVGxum3QkgugUL/SrgdAnRF3lbby540eKFSzp/L9LLwh
A7t60m08LzbComKFi0ZxCaCC4MEU+wzzGb3cERkqAtb9g5NRHB7GK/x89HJnlX3FYLS9ge3jovSY
IwJrAJAGJVCAIAS773KqjN0Dahxtmlp0oEXxVA2TRqm6qcAufCOoLGIdOEmAFY909UnCUlnPJ3Ta
w/Obs9d1+al1Y3gyU/TrMNZ5nLZjJZKGD01rfuOkwAPu1+IOMIG7n5COIEXhYTzeg3xt+TFmGahT
+w0ptBCjp4iLIqykxNFMbLrwCknZ+gcfZHcoWXt6Lwj0aYfm/GzsQxaY8wPTOhhoQQ599mC5WG/e
KaUY0bd4UMnx01ChVqK2MhYwGyxf/b3JUgoGEkrgJ5WU1HUvTNVK35vGjqNqMEOEQSkgi1gUhWkL
vpVLW1aJuQXF+HfCp02ERFUtYOo8f8Q9fQEo6GfzHJ+Uip9HxurIty9WdPewDqIhOh2l4DK7uo74
Rl2Wpf8/hUELCf8p2Wpr9gEMrZgHrAs7Jfq+sbyfmUUarDpiS/ZKAuEqN9PjL30tpjxpvEeytRZ6
vW2GWKzpi7RBT59QS2ZLBpfNa4Csc3yKrvTtKtG64VednEWt8I0eYZpaAHsifqgwPuW2lTPvWK0E
/GYAbLHsg3F/52ZZW3UWLAhX2U7B1SZj5tcEfJdOiyXwmJJgpqoR7o2SnRrwHVO18uvC0pw4tgEO
fKCqZ0Uj+b6JMFDKjsnI84/6QKft4H55g7m9PPjfGulBDQ7o5XR23sBG/N6uEAblpS+SZflK68aC
0VqgWvB+MciyBbNVKfRPDAj5muyYyfTHNbQnWj8h5+akKs9eFJcVXNOpFh4VjVSQjlST6Sq1XVfJ
GIXFaJYtPQAIeX8GpDvnwPNg+SyNleMez9SNfAO6nQWlFJSxlE5hLwIrfGGq9F8gUEYrf5vkxSjb
Bsn/IYAeNOx9x/JVn9Bn7do+reDKY5JvaMVqsd9Y41xVswQLfSkMA8jVBpmslolWTQr9WjZklDNg
nEa7J2aTTSsFpzel5KP2CztKhEdbOP1LWPEhf1sl99QGnTnKH1yXf7jxH5qUmIpawijf+yWdWzf4
K5WlPLKGJ+79BhdPujFJRauzVMytRN/s3wAtJfWuZ4XRt6iGnFma5+crarmVaiw+XZNOAgzBzdfm
2DddeN+Ow6Q8363LuEoRvw/n9OF74Nc1YLwtekvM9LVZ1W2CZxMTRHWiuX8BVtoZPCv5fggmvouT
kazmf9myG6Aelc9sNpL7hYjOGmpQtp0052zLV+mv1K50m/0f+AoDZwlx1OOM1rCgdgweL/EYR7qH
g2z7CDS/m2BlwW18lcXkujyDanr+zaMVCJ7aNwOoMBK5XfbRY7NcNv65hfyQnjCkZ9+Jf2Pm6oCb
MUN8Yq6odQQ/Du0L3FNIAUP0DANkEMvgsx0FbF/5vxtdl5PEsT99ckOsDjp65rZ5fZT0dSDQqg9+
LFRfJYfczu+MGq0oZQP8BFqotC4Pbz9v4v6okKhbE3QoPaxOwGQRA+12doDLR9On/VUhJckiqZjU
4cBcv7J9IHDbIEoYFHl0QmP4fcG0UQ95p3PwPgnuHXHIQEOsw9+G/0Rh8MGRKu7kvc6oNXgdkvSy
3EfizUV62ZymA6ohPu/6LiFdov7ZLSZGjqpbRjkkpKBm0ZsB+ULx4PZQASqwO3BfOeWcYTOMz7ec
u5X3mDnukzBhWsfgQ+At6BFx6fI0pKWwzhQ1x1cKrkPNrNU/EsMgbd2i/j5eOhLreWQmILcagFB/
yidlg68tcDm0cvGGleU+PeGRhpOUsFRjsbpE+8StHVEnqZFfiBZ6Mfw0MHCyRKYmoclv7qJKf05K
6hG48WrBqrC3mqAVRdBzp2vVGCrqTN5YWHLIHDcWcCp1etG3HgKH3G1vxu/f7jeJUlsMEt18TZfX
XLrpJkoXeLQ0hmRynt++4tG4tt/L0RL6CqBlcfFVNbmqTrriyX5JhFq1SOrdR1TGpEuGjn5Eg6nB
X2LTHxZ1knSq7X1ckV2ZpNHSxmwTPAYL3DbsKnsL+zFPhoEH4Mrw6eMwaXuvibhYjRRHDcA82Bcy
j+h+xrNfSF3/8HlG2pYo7X//gPV5wGwl4pRSVUu1pEyfdmH9ZVs8KVbYSnWjt9M7TBn5VVdT6h2P
JgxsbDTycJaxSPdeZKSaIEVZhDuuhgUaLDNQGdgbFZ5Ghajq6BL8Bb64/iE6xzP/CrXrNMCJgUTD
JmdViLLfvmAmrqesibEtpd5RK7bCvwFHOHseiilfL8p7b5HpXCF9muE44HwxIBRCVGXHg5WOUe/O
FkxPyFNCd5XCqur8c4dkV20W40lbYHChbnDVkpPktiUUUNaR7ai7DM+nzOuDOyBRsNmabDgX5era
zV2w2Gt9jZm2ni9uJi+hiKd/ZFv9JBC6XnJ0U87iXq85i2k5CxNs6CVNdcthMJpTfCU9wswsHsp2
lKO8CdjjmtDhwmUwvptB68b+zWjVu9JdYpuwSxah0Ys0GAD9KvGP/urN3mgFiRxx1ZcJ4U/PFaKd
HzV2IuvR6pcabaJu6AfVvAJc6t3uRFP97BCJHF0pXlC79qtXYq+dIUYm+YlE0PafqIaTQ55IjFTX
FGRqK5+AjkDQDQoreNXMXTRDX8HvSIOucVOQ3flTqoDJct0onqXx81Uuf3sX7gI0JgoZ588fKGaJ
XIWKbLWhZdRe3ekLNpi43uUbCOwMQGf8W1avg7QT7so4UnfF3W5bAv/i6g6/2dd5eemixn1zrUYJ
A02IZEPmGBmotvEGHE0TgziZM/Xx7SY955lF9wV5RTWVBGMA7D9kbW0V5VwiEaDq1wJcmqk9CCAc
e1MApLEa0PWw6A5jI0ULYEjaQ7lrlNjnk+fGVUL2g90hS/0uXS0kuZ3ceGmyxBrzKvRFiOBqsU3F
brxbQ8xG1Xs0V999s+/+lr/eoumJ+0eqdwjQlYf19qV0frYbg0xtsx8QKqFytRIxTrenOY99YZNE
I3isS2HbDWLMab58QSc5YekB3tzzf6/HCh/BOPDyAGxhd55xvl+UFoyP0LTYCFGsMRKsbffz0oQe
IZIJeImC8YjC7NQzcxoGqdm1colrh7qNsiFp/l7A+n60juPGymrPfOw3nhvcZ3zg5jnEgGNuZZI7
tuDfyvdCuBr1+tIvDww+/Wis4VuGmBwDswxHB2088KDd+jPEqsvSecTzV8gxyl4wEZdTgrZJZ5Ne
qaI/8XhXlozZ79iPF719RYywijw66O6foS679uP07UHsoukFmcD/VCJKsHM50tuYA+MNee0sUW8b
JhNbaRkCtOtCTFvZzFOcAJTsVVEfS+rSx3i3deqxslAM0XW6+VMwAb28JkJ+7726PGnd6C7N3n8N
A90W+i0ZRYl9Wt1Sf8ccowYzAHPYzy0fDE0myJyxGVVbvXMoAiKEFwueRXcNnR5rFnJU3hwuI6t5
T8LCkHBDjc2anR4+Q9HXCa2/CBgiXXAAHq2gFAQEJQSytfWM+1a5VmcQ0pvub2Krmui+UEBbLy7P
sVv8jbeVWo7n0WG+JR2sw7Nd/JvSnB+HuzNcyur3rvjcbgsOSOmUIgTkeE6uCmR9B4YKdtX/aIQe
XUkeMUtJVHd+b8rRZ/AZ5FoyFeVbSRyOmDa7xvjrUeU9vWJ8zSbS2mxy7iG64On0M1pmvzBxhhmf
uNLATD11Ng9EW8tsIYyD3X3eskaHW6PrQ3gdEmhcIH9eeQ6tB8sOfS9pdxGRKxd7r6jI5snFIGs9
rktHUOjEUUz0+PT09NnXkTmRbK6q+VsYt1+pewMAmoCNPy3qQn+qTmcmQ/R11c+PBpKnV42UcbrH
TT7uZZTGvEJnClFWEg+PyUw/5EFBSSw3k0T4IMQjSLtKOf0qiAGo1Dt2f/u7iFDfopSCwZG/n7q8
yRwBYXho5CGq7wJAYAwTXOlH3g/iq2mm6aPVjvn2czB7KZVYQd/8/R0L4e9NDk15rA+jcMLBuuPx
gV8N2CMnNMKJa11BRc5LABa207xKKbmkltIGnbaiTu7nBPXK95+S9wSBNXDxIyn3FAOdUu8YMJYS
YtnxSsSyBl6PBgEiRriphJbC2WupwbRkvqLZtnSsQOaJfOEr3NZekKFdIRf0A4Smo56KyhdoxN2z
NU4ELwGcVtpXowQ8uur1ECswwpD64eaBtg9yma/Asb0QVohHU2rmTS+yYkdo3o6i+gwsA2bRwhN6
SUbTCCusjP3YOeMLbvS9sER/2rQYj9f0qx4ogcY7h25AWryQy3DseM6S6eIxBYYsF6qtVwc7NCBW
GjTu8QqcHVhnii1QN6/vw/fLFTfs9BrYOQcZ5xlalpk0ZCs3f2BfZyzO9CLDN6AXZuSpbuaBpFsx
DjjEqG4d2TfivRw2Mr6hNHRy0dmBLUj4Iz04rn15ohhjIxujSi69WWEXVh17CFITq1eBd1xDF57p
JPv3frZJM1gWcR86uObijfMsYg1A7UtgIO1RnSfVhH4BvMXH/Ky6rEMkEhqL7LYUf7/PstvGa7Tx
k4dTU466YaSQRhVQBgX9W0HRzd4jsbqAb1TtpxuT+Rr2iQTcxxj6spvp7YGdP/Q5QoXQi8d75wJL
GQVkI0pMcweS1RB9CGlxdZPiiYTT85az7D1fEJhwN1B99LDrsZClszz1H8JBYlG2X3thkxZ1Sp8x
cbo6JRu3tCgVVD2IN9uLhFCuxYNGqlxylTBDAnVrVVZNAhQ7MmE5zNGyJU78Luci2CW011hXJtym
Kcx5BX/4QWMuFkxuavyr8WgILvtxruqCD2KjyN15WmM18UcOywgK3ufgF5OsTldF72kNcYosVwNV
N2rNtsGhXtuAqRJNo/cI0W+P9LkhM2d8/kw7RoIrB6peIHKO3QakvZPAUiByJxWjZdIx/EpYEOky
egzVRnf5kzmww9msbXosiCZVG/PaI6CRBX1DUQfft4dPXvBCCHdQqSWyjUFBcsWegEQ9HyxoApYm
KDe5YVtVGQlKyVk9yWSlBUKHMq3fciC9z6r71qLRaeTEGp3aiQwEfWlG+iXBaTkGtX4dlv2jLJbL
PT1xZavqHAp0snJooI/jVH4rbC23YIOsg5Jul4ZkLflNB+iRfai+ZswyedH6lgpaMLSmNXJ5sBf9
eg+EM5Mgwj4P/GNUsykiZFKfQU+9gwqMYX5c53iIZj+/aJpN3Snw7kmm929fXqXJzpnrDfZfgJmF
gfZxcPPm1RUd2XIyUetp+S0dNBH4lZLgwO9CJd5TfJOvTZz5p3XYNvxrieJjTsIBMemVKIqcm3vQ
JaHY/ncWLFgCdOtvHOZcmVVbw74ztD6mpT5ypNRsyo7QbzUWpcaEPSlaOJCKnOKSzI1b+ClsWW7D
KGObTjEatOAIYcsMMOIvLZZTgyN3WFIz2TWaRdDxGTwhyxGZnZgO03zIdHQLD5B8VFfLOexsMAWg
Vehktn/iHm+wGIGOsCsLi8SzvHk8VIxdF3D6WscHTTAXmUH11WhUNRVtMALSUI3AHMW4tJTVeUjf
42q4t4K+qeXfD6zSTFgOIgrvamzM+XJoGu7md+jZmgCHoenYVwno0HqKmINmTteoaPRPFqc9zkpk
pkjcVo3m3ma0i9OglCaA4NIWu/CbDwFS9VnEoa7ex1cWOt6Q3ASHy7LppJFfPbPYStu98MhaHS4w
DZorzie/p+l31Yl8adIKVJ65InufphcjUaD9r4K6ABNRQxRUNMrS8hKqFRuUPMryaqVdyQsrCbke
k5aa/DXPNNwtOL071m9OFUtV0s1JLeM4GA3PrfiL0TJ1iesmjPJKJ5/onXPcxfW+4AbbS4xL4tXu
aDkBineQLGwh553+2NxvzObZZ8GhzJafngSKwKGuoJqmysnYe6/fgmlR+wgDSR4uUBWZVxCgGSDa
GMXNOiGzyVW2/zEO+jc9YbTCqi1IfSWfB4VZxSMjMnjeFhBxWPDEn7rs4cRUEpeldxo+rE4e9W+2
X2iOHekzj4R2z64Fhht6mHIKXN3IwJYCuZ+uJSeP+gPVgvSQHSblPJbWjscKpeLlnF4qgf7REN01
N/iW2TN11RZPlcvXkZmqyMU6XlkfdjxBsPWqBHLmlyxMcm0hzkNeX/q/QpE4PvL14oYuhLbgW0Qy
GN885tdNPJceac/1bxcBO7mp4PgNPpZDCvD0pKXt8+QXS8dXAK50Qa7XT4fnRDI5ELpAdQcYYOW7
CdtDN+v6DAjHM8hFujf5oJ1P5v+UEpOkhsOwlnEDo7GfJNUTtoMhtK9SUujBqYK1v0JILOpd9KBN
6B8/eFA7cCQp850AghvGuS0YsEyAgikwB6uYALm+ksB60gSf7mV+1zGzk7QswFcVfih35cvE1WtA
4oVdbYSFWOVQomoP6UMXL7cyami8ttWZ1CZnv12SR/8hitpfoLEmc3/vU/8UvFgvkdlR2UBI4WxI
Bahy6yrvJva2n4dKHtYZslmYDyP6ZWze5jcnI+wXcIvreF3GhPW57O4x4NjxRyD6JZxcEYa/YJbh
Yx09g5+mtFwwovAEnr39yB0JAmP/oX7Q37bali/D9juj+KwK5bi+HyBM//H5JCUYyaBmL9WPmMrE
EujNf+JLY683U3DEnGW719Nkpnl/8dg7CuSdUsFTJK7vQJqhzFcbC4ZFDjxKN46M/kV0OWBn60rI
QYnHmTJKEo7uQFfvScrq8NiioY7jMKrUizIT6aK+kiOb2ZDeLQqxi8Gfckg7N11c6KBcxTOsBphq
6YBH2x314GMVBYc9z/S/MLE6+nyTKNuc3S6QWu0F2VGlc4fU3HcURbRyAJorw0YyxqgcN++oy1u2
N4Bq/EoJ43JtAkL1Ctc4Tr4yrNCGwA6gVjIoPeVPNDUHmZCo2jgZVAmD+vZQSgdTE+6FK7dBvccr
IVOKjIJYbm7HDng57sFYQASfryY/SejjxFr+9TrcdnSj9hLR/p9VrLIENDBx8dGRyr9UFya2+IvK
6rGhFsXhbexPTU41dPG4Dlip+Csvbw+54zbf8sd8nGTsDxRzcKdTRskv4sIAL7wjv9uXfr30D+QL
bjaixGI12r7lcJKEwigW+b99tBx7TQUoGUSHBf1Do32WtadpyxRT/uBudFtL5XJtRVwIxnHYAiSs
Dkxhm0AR7FkxxjoH3VFrJ1OODWfRZ0NU4tUlwPJUjwK2Wp86hPIj0Dp/sWaw5xkBPrGj2yl6Qoe4
8Qdxu8YdTg6J7uc7r1Pyj0iwBoexChoOqwaFKNsmLJrxp3CA6u1dafJGhhZdJYe81f4aNZzrtyBb
3IvgCcewFAZcRmzG5hfCX6/OpOh2rWZns6ORRMupTPyCwdRAHx9QiuqeNrd3F6erZewajboaA4Lv
uuc+wNYImKZi4wkRuYYtN9gfs7eTbhYgEGl6ME6F5DLqi3wviju0EBGBgu22K81SQ+YDUYHUKQY7
s4jwoBX2gaFJ98yTxCbE3wlWZOtUfvjNhrRbSxCNKoFHJmceF+TLqKKeGY7dya1r82jKNe0Zix+s
mvoUb5CBIK9s166J0iUQxPJrjrW46s2T/ET5g6nqLN/mQ8vOuj6zwmZbbmqaBaVaHpnLkDKlb2cy
urfceYPqOgzrHec+LeXekn5YKlHOr5XIx502hwBlqZQ2BMtKMpYwiqZrd27e6l8qv94Ez+tyk3gX
dSgYx1M0maU/zTP2rxVnKD/f//Rz8Q2StcNTVgYUJzKqcuf6fwgJY+AD20RK/BlNSeqU5TFeEDXN
3TAhKOEYhwQTahjk0CGs2bJifo/3WIDQbnvdaQrDVDUyP4HOZOujZMBXmPweHU7L4GnhfvuPVBDg
NG9rKqgMi27t9TOh0apEw+UCqQ4d6qdVY4XZCRF5Z5IIBEA/IgvRMTCfEAvUgCY6Q0Xso0Tr8zGl
GEOxwO5PmShzCdYo43/HU5TBgdOLqAgVtQL5HQbhH48Z/dbYebHCbHL7puZzvf7wf02LP7gzIBUJ
kB35P+2xYJijlgzuKHWJjPDm1qU7zm23tDd8DgTecfOA9/utIv/L0z1vRC7ztqtW5K7iPApylD8q
YwnMexvKJ3pNksjoMRntUSfWvv6X79gQubQbFxamSkF6cZQpN8GfopVa66MXE2NR/ZOR6B7bk9FN
ehqUuwra6bRwamMkYCMzEMNBsuXcfokvOxkqTEgG69x9fprIfk/QtmiuBRo1EzLBywZ2jBB/5ila
jTrE7z/0GOeXP26ja23g3VEEHcY3NZkhnVVcBl8fvO+qxhPqs+mpGlcQTslOmXXdVNlWToP+Jv/Q
urSiSSNAhccsMiKg+CXsQ7LR+s0+cgu/5UPx8blMoHK47wkIfMd0nSlbGM9vsiNdw2YB5Qjh+653
j7a+pz7sAojaDGObhFuDMc7sC2qjwOj1yDElwVHiVD60NmHz02ArhNGoEnn62kNZ5+gg8Sje6vVj
8PaXH1ikg8YYg8xpf3HJpFJqYMq6nptk+IaGuIxT5IPs4fsfYLHvd6HFdUJHU5KaKxAdRzt3xgFS
0+0WdAfQp2DG2J7XKjR4vFtzhYTjmUUcMfo0G0JG5O4QuA6ZYHjGS+Y+pMEqxMm2qPBVfUy1a4TZ
+1GFRknCg19KqNTFz7Iwm6N1fVtNMWKzEpt8TeX+6bQ6ePHCPkALeRxcsnTa+nVmQPwHlduguBrQ
jzLTvJfQ2enBi1Lh9C6I3ag5s+7ggsG4K8klU3fQlB0vrQvgGbyaz1D7wS0eTNxD06ggumhYvTA1
x5QsbQ8VvJFJqqiQ55uFiSERgilrO6M8P9vUezn7WlEdLkRNfc2Wv4ygEEMN0dV9PcIPrmSm0xcf
/dgrDxxPjWdDlvtcnr6I+DNkWmYGXKa+qva86u0Onfs79OavBBnmqp+Y57YfLGVK2F9SVjf4Y1RR
qs69Qqnwtr1vmH5wiYv1sb3d+hzXw4ChfWivvQzDLHsvar9yD1fTfITRokMqKsFL8va53xSq+2Bs
dUI6Odd5i3jTWmcGKBPCjb6PNW4+WT2tiXH4L/0xkNIcDxhcENLEpCgSN9+64T0SPWHrAVxGC1FU
YgsPdaclwX7IrdqKa+OczPwmbogpL21zTbYGW73MJm9LgLzgzQr9d2Ha9xah9ABMbIiq/QXuvpRS
yw9uMegdT6wBLm2AVHn3SUKN4oMdbrJnVbKKxvZ9HtH6RbeTF8PPBIHZlIyfAa9RA6Jv3kOZNAnL
5cr6ipoGvfouPPNQWdwxGedrRapBfBhi6NWJZTDTWMx3HQNnbCQvmQfEkwR1afFjzNCZaDfu8psl
xWkRkEadSGcddGaEnCtZ5mvpN+a4P/2r+NsNJnozMsMQCyXng7FAiStnqvCkOOOdnbpN5w5qnmmz
hg2raRrWWFijwFWUuyTNpiAyJHAmeurl9ZcThSuKGrcJX7Ckl3cti7KNFceVPXS7AwJOAuamqLUq
EF/IifVquuxUMjnz8IBuIdvKNnf1W5fO8jQZb8jQH5/MiScVkFPv51WBhvrmG4kPl+x+NhsGdiOU
Z0bbisT9ZS9rK3/iW0aisphvu/m8wdWhzdtWnLtc+mrO6r0T5gmtnswwtWvf0IARJ9ndkSuX2q40
jWxlzE9hFDc8OyOnQzgsenPIakB53ExLZyMaWlFkB7bhJemb6iCRpiaF4qmj7wR8na85rAVM/AtO
5RFHQv1YJN0RPKyBA3pUtens6PFhFW5biVdd0pf3zvUCet/Ru4lRMtyA8vSkNOECDZ4LDcOR9voz
rjSyX1GpmTA3LhZn4IdigLaKZMh6TJPtLTsM10aD2vtqMvJPFJXOR/aVL4mK4zIXavGiBZ1RmzRv
hfJuZJBM61eys3XKqptJzlXwhi5mgWWzezm8FHhBvjpDEAjZ5m0qEYuGwLRKLdMMFm4KfHO85w+y
CkvSj7R5vWZpcPuvyHYB1Ki4AMqcu3L+lr7l7GgznWTnZsOLYE/G+YTclyl8C2b4n+pz9zAHeGcJ
VirShkQxlyVYqcmxJRtXWcxLwWT81SKJv8bxHyjG0S3YGFKhd6x3d8Rt3ERsM8AiXABCJxxp8Wyd
Fs/4o9Mqt5ZceatWEiVznyDnYGZEm7ru4D6iwvCo466wCE8K3pmfZ+QK9BldjrlDcF0RsD6aOYT7
DGMhRmPYfZRGltTM+2y+sxVK+00npb2QYnhGFjpDtacml4AvKZf9siQNeAYEpyBxAYIdZL21n8BT
EjZwfjTRqpJWxJ1AfjTtXXxDFn7QJNvZregnmyqjNFC6Ut6lxKs5PdFg/AvCa69D82nN+DPrNjfC
6VW+Q0vKbf4aMaZroQ2RMB4lkYOmyXj73FjCsbYAKVRR3nGgPkTmfKV3Vn0H8oUe1J7y2hIJcnV6
mbKgBc4wfGQNTiJiD9Mk2wbNlTwMmy6sza2PirOHvu43ez4o7YxShsKhclQyk9R868X4FU3WDVoi
otQWD9zDY0Xkno9k93JVn0Cvqbsz0v/Y+YIp5Lg+FqUG2kCpkEqzvXVHOlB+cutP+02UM+A+5WQy
Ja/1XPEelZim9Ha9NloiXo7iXhDKJPLQi2LpunCKaFtfKofvTMn0cnq9bmHxCzDOAepwZNLFrjmD
PBPG/xU3n8VpuTM81Fsldb7CEQYpVSdGWzpyoTgMl61QZUi2aJOUZNTse0ikUe/ySbz9BGbO9WLU
lEB+b1vp45VT0/vzhh5aWppKXIvlfFrNjlIa3Xf9Sc3B53jtXQcK9EgaS5IMQMbASTPGEPvtKu81
Zws9umw+LoEAtsPIAAJw9XxaajE2IfyhS5P2gQ8Hs0zVq3wRk2vq18N37BhpeIGmwwqVdoY23WGW
x4zKN8MIVzuvXl2Ne/ctzUXrcgju33HiHu4JV3HHD7jDfU44d/NYMbzwZ98VRjPbK896H2mxFIg0
bcQFMybA2P/Bizc8QK3xslpjDsj3daGNVeoPJQ6g0LqffRTgGpohPpIalBIufwE80hXwUVLqRzZr
4OalDjkzukXEsnfqsjatY+fxk9vX/DhJ0m/0whc1vGlZI/lhOudlOShni1MtIrVOmxIgQapuq2kx
ouNm5UsVVpc+M6hElUr7X7P62STaBCpUVD0r2PrVygvx6V9ZQdzVexdxE8ae48ALJUIsw9Glt6bC
JbG/P/9tEEm5/DXG3+IojLt9eqdzYf1lMPmOSsEKzci9tePabyfkUpmGdwAXPR2rEx4s2OHEYELf
jCWntWT8sDq/BDRoE+9ILyN5/sdFCdyyF+x0yZo9WzglsbNw/jFpFBCr5tNGwwIHIoMUSEik6oQt
DEyj/0+X1gn2jHbdRmx8ePcduSbZyNCcdiok2uBphiS0RUOO94Awb4cEyqH+Y3TXawRSyqGt83Ez
N9NZ2NsM2BtBxs+Fyy+a1Xar+3wY1yld5COCCquI457JMqgZp9Nm0wQcDtNwTe8XYz8rybX45jPR
oyBzSwq7F3bVlCEekjkjwNsjBw4yYvnzaosID3LoMAwEJHXrKVwhhCnXJ/HAl/MjF6LCpZidE7tS
k/UQqbnaf5J7K92fjbooHOAsYIt50SPv+x20wh/E4iWxMO4nDK4Kp9X5s8RjDSI2DaC4xSDDodQa
6dn3HZ9cUatNOM3NwU0r8e60bmp8rwB7IstEmb7wCftd/oGNMpyS+2nHqOcUc5SNtGf2HkZM8Ifb
8TUAeKOqUMTTo40LftM/ksyfVw8fpLofcn1Sfv3Af2j4kJW/GvB46xsHyoVRaDahCL2iLvmudI/G
Y1aYRezhIVoI6W2vDrRnYKtXygpd5p2a9A5QrWZMljud2Wp6+6iD3d5T0eVSfvwUmgNbfjsXW6WR
SurT/fLTyEbZaE6FNBJX54uZL07aoB0P6Z4ht+bQfHKhfe+UoFrXrgaennHXZRCKoNw35xOHtjkb
Qw/FVLVmj9X5EkEgYqwsq3FoJ99jsEoxWOBhV6qYjFL+XYFCGX45cvkNyQ0p7WmAOwW1DGV1SbwF
12HyJMeo2v8K53MH8vba0e0p8rgpP8jpOyS00C7jWeJD7JtypmGINyzTTuD3MNt9e9PojxRRv5PE
vJjVV8dvN+/XSGKLZ1wM9lXxtT2SRRvUqRqb8ka0EKE2mLu+YHBh6JGyKXX/ZwflIwoK0eaMmstu
DhbP7sxVH/YRT0lfk32KRBVljornhU0QDd3VWFP1bVSqx8uD+rpbMqMzBpvIKWA+pOzYhyHZkMGK
uHpuUBeQaG1gYR4xJJdM1+vUAnmYGz40lVuEdCiRbzhjzx3SoGGh6XlugUatbFG+DwWMn5wnPABI
c2CYuYGxFx7nBDR7WkAtJFISZ0JxChgxVImW4bKzpzUs7CXbDmIWrnGsvry5YDZ1JEGd/9Gy2r1S
VOyOVCOlOW6ao/2UvsYJUG+JaOseg9dWpy8PmzLZ4iVimDbcmFbd9v1HMTF3zA8bHMwrYLe53nf2
LPkMw19O9lXsEjsK4VAXfuvf38nF5cS1Ea69Xx83SrOzzo2ui+I19vQlMDYqfFnXsIdf4p2s70r6
s7lkGnDqiJmLpqZqsyz2OQ0Zxg7E/LN5a9UrhjRR4uB93nxYQhwrR244McTLul7UDeYqMWXVnrKM
Vu34r/5z07wYnNpR28bjbFKgkCewXzrNkZH0vBEnrKaMMx6Rng+PFhZspxjQd/IKEW2aRyf43muv
xoL0Cm3wvJldEYRJnQue1Za1ZZrYapa5lSwTgOBbZ8vJpSEsKbxrILIz61dlxCUqTx4pbety7C2Q
AGCAiPBFKzOTIMMV3OvEKqEp/6POmtNg+Dso3hUGddP20s0mz64vLtdmtDnvEkSaL/xOBRRBHIXH
0pKlLQayDW4omJ/VjH2oXduiz1OurJJcbCfrvUftcPufQBsznWmCwVAwmRaaHu8BWSEbxLB04rwT
kad/B6KIcBOZ99waaprq5CEjHO3/L5ZF62dBdzCYpoVcclZT5v4jh05Qztok5H64jBXmJpn7dohT
Vp3FeUIw6B0it3I0OY1sDpd5ENZZMYAUOnmLrmyCUtYawaPFj2HQIpY1KUbzvB4wVw0/g7f62WKi
L+V57VuA7S11mjbd0torCKVQsaOjP6jQ9SeHwGyPtzmCpfS15aHG9RpnybWDmwpDM+rKu5LrxzI3
u9AW5I7oCJRRrV867lf54yq2y8RmAK94KpZLhYrehYiNmdzI7Mq2+fCeiivNfzIGbieuYYcXgmMT
Lkh1QQB9ROkg53BNaAlgaQ3fxwlmbhCv08+vhdMO2SPg1gpoJ3m/J7g9fDfhFp2rAHU3O+0I8u8g
76iiNNectkE6nIdGypQojVbCX+LYlxqdkf5/i14qUuj+MQvXetYvUtiOPpUq0yp4c5nZuEAaQMMF
G+tMuZN3enn3OanZE7VWSPSvxP26TLRKjuoQrVhh1mEPyTFkfKv7vXSlkcgYE5oXbOKl1ZmOT5xJ
Gr4SRbL68jZQTcSHtdSMN6QOulFppYKbcCDFRHj3/+O/3byqjpSJ44gkLPUdIf5eKlRKHiz6rp9b
vxWzeLViJKP4+1Aks5BegdzHTDXsC5lJnMElvGXNBZGBbtUIH94xcPqAtuewJe0yQ9fDHf2Mg9kx
RFb/oV051OS5S7Ed1hutV2DZZLdVgUcCyGfv4Ng60xo2IE/LTZqRdqzPKIGohdkDTCsItxx1g2Dh
V51l4IlpOm0QPuk6oav80Qv5Bf/ZBVdwJdUdy0LlqJmKInJYlRQ2ISiyRkI9Tcfp/F9XPZtgAnpd
2dvxJqpQX9dnifYbW7x100ZXiBR8+4pTMcOlKaBepntI/AsppGf5FH7ws20mD8t8FCP93yRgxwJ1
bFxiiwN8gGkGXNr8NgL0dB5gjkRmP8gPYnEthMqdTaYz/ZmJQyWxmDgq6GgC4YBrjveBV7kVGmQV
1AaIsPQ8d5She0NFQ6GKaAD9U+CN5o2Eik0nJrIoBMn20qTy+CdL4pi20Rr9JIuoh5AW9MkgWg0R
5pcQP3kJ+iHLxE1ntNswxYM8qm6MhaT90Jx90N1mtmmqKejoyQHxSUQKy2n10wWP3QeqL4Sw+uU2
Ec3VUX9wxCIxWa+74UAr/aQ5K/c1g9DSxPPkEv4/55GY3S2LdJfc5uUQxS80TGi38+iGQkNOvxNr
5P8QdCJpnFsOkHQpQnspfhcLVnpmGGCwxth8VK45DI/kYO0gcSxHx3MWZs5I7tyNBoOjl8AK7KTu
4LMhN4TCaIBJHuyEex1m18BF1anODMNh9ItVvYGd7vdOwEiBW3dVjA0BXmQsTlRzxOGSCqGmP8X6
kJNSgtVNwetlMUun0NfX8HSMR+4kIZktqZb6SCssx0F7KQdNNw78Av3Lx0gi49LEcFsdxLC5coYG
R+i9I/vUvgOVQDHUP9scnATVP8vAOFp3Ua2z+JfPv/2U40syqd8sjiBQaAAHLtyUOwYuZcVU5wdT
RDLg+v46Q45qkJR8oaZxTCci78xsnzRJe7FCiTcbsRIUNT/JM3Xn2TxhGmo7Nb0M15NuAPBuG/Yv
DUvDK82lgLs1ZoD2ofrbr2ZkWFkBiMehqgtmctdxgMO6OXooOGSfBuIzHz96GCWm4W8pGF1GPrKu
c9BeI4LN10OKBIt+2t1CXRXLSyAe3RUZHGPXmKubYasQ1r+xi2vezpI0w4qY9oYDHjIwON5c3S1z
f7Hc+KJBFrrJbN0TuJTarkOMnma5cdUqT+nCF38axIqq+QGbxTc7kLf1XqnWwKBlM0PS5mhkY4Kr
VyXZofkLt24tgLFCGwDKH8XQND1hmIXUSqNAQM8DHf789/tKcvMYsJn4gb1yzdGuStVo70P4F5bp
KGaqBdYUuaxtsalZvzO2aM7hVYAOEk6iNCIzcHgr/4XBi8u2riKVLNqmhOxPAtqefQn187MFDcSu
cpQqzGY/p5fPhLGUZW10WOtwy1pvaR9cDJjBADDq1XK90ShK1OchO4jRGGkyLqwBc3iJAR+Jlf+J
yTEBdl1XwprSsHMZZaOpLrj9H0eHeWUVRwLlxGMnSeSwAIFf8ceP6ZCEeu+6YIblnDbI0kEX6iwo
HU2rVYeS1VMZfIXtXUS7IevFS/CQONaLYixXwplfY4+4Xgw8A/krNqR0FKEw3fyR54dc6+E6e7bX
X29xE425kd7RdbG51RHaChKhzS8lWJk+c41qlihZbsgseZ/MJLRB6MTRjWGUdS0l702vsKo1lKAG
poUj0hHnm8iVnCIEto8hqWebYPtoxXwcGnLpuCHvm9oKR4i5x1r+7fwGfYMUQVgB9mswgO5f32AM
fniSJo71PvYEmzAelxPRBCJKfXBl88l8BO8V26R8KoRfDLd7MBP3Q8CHlClf7YDObjN27EO26vkP
I9A2HJKe2v4kZnCwAjZje8fHUFPkMXqb+H6jVUQCGyvrGgliFooJFk0fqC5f/IElJqyMLw6Pxg+S
1InhtXlgEln4SyAEnCoJuEV8simXf2G9C+JFl3ZruhnpcPf1DeVwaPpKKwkiGQNU9ZxrDMkiQ3FR
uUAhmaZBLLEp0smfuyTTZbhhTRF6iL4BTQpEbnFE/Un7KmTdxMA37kV2VFiBcoLKQE8OnnshXqs4
dfudxvT0TbPInRBO2C6rHWIZ0a2xiJ1Gu+8rQylOWi7Dyzez1e/sPfr1GEXWoRSB9jPri1m8QGZw
wzipmQhqf23zxLGNP+S1qkD+ZyDEJRaO4RbB4i0PpN9EuPZmNuXksc2yEuX6BuDjEAfQQh+NYH3O
kTI9sNPEV3ZLEgBqn2sefbgsva56Xs0sswNwaDZiMxN2/zKZeGfry2r6kezIGVOARPygj7bzMIaJ
Tz98JaeAXe+VGycXQkCeqPmooU49V4tzNauqXnRcBGsdo7xSAbkKo8BjFW8uwSAEHJAFri+Rdml9
Gy/psKaBLsachgo3/Ok18kk67hfmQsxB4F2NFguGpBvXQJHS/UKM0z8EWSxSHADnQZYu8Ya5UlIP
LK5JPHpRGKdpHFbZpc2/vBKCbJo1FJXrCiFU3XMdo/rmLFhqwjroMndL3Y5DDE181h+LCVoVcEr6
whaVIRoTdU9GzqkjL8Sjo0/aRGSal1bhJ2c69SC2BfZ3vVarz3EJH32V+qbn5BbqI44F9LteUgQA
ML58KiBYWQR2jS0hX6QYN/xvAWxwlhtyFGf430mEFAFglM7vT55KTSrmfct5yX/jmScdOCkAs9pU
1wDtCnjWmwVW3cQolEnIK+DTqEjwEkdBLeUJzJBBtZ76hYDSDFY9CpyzrG7Gi79Vc9KUZ3mn6DeA
p3qhXHYR/gHG0kFlS+ZJCyTTd5BlNoM0Pk6TeyqL/TY/epzru0ivb3sDzYyQ++p90fq5yTbV/6Rm
BKhyq8Cq+KlRlVE+7E4KhoyAhTdq3dXIjfh3L+teZqsquV/ib3IN3wpk5Bt1rI0mk3/gABIzcJCt
1E7yfcxcuiK/L0hWJJT9iKDVYQjHNB7ep8RsfwQ4u84JLqQOB0cs6mJYUPYIag/K8mEq/DqQLKVP
k1L03NUQhn8vNJErwbvRaOTLCAPkXPPGJcfac0AuOdrJkW44UcxkO2fCR2IfnlKW1JlFdedFQhTi
RsisNgIbdUIGonauYykAwkWRGDill4xUWo5pQJ0fNy75cXmg3N2ecBD9kjBfVKAcA0fHLMNLnbkb
/BSuLSCjh8IuWZRPm/qwLTZgGnPiGFmt7q3gxDzG50+0cOgQNfYnFWPScGwIshc7v/GYh01s7X88
n/Ydp6f+Mlk2PRp9LGjje9UYdDpgCatvmOvX0OubEiPXI60hEBXeW6HXl+DZtkXeFFlmUpBgnOWu
MWLLhwCL8H8ZuZn4hiWRmSv7WniksRW6LuoTblNSZ/PCNEEm5+MLlmS8wwSurrbVC5t2L4yIxEzX
aEvP6qjgYWZ+hKXEeEx9Tr+sGKGX4q/qb0rH8IF/gugnsTH3xp52D7EzfQYB/qRQPI5Wxs6yDtGP
wMtVrmx1px5Lhm4xOrz3PuiR7fKEqz8mT72V0wrai7SsUMr5/CDrTrck+5k8Nmfaxp3RzOej+59Y
Mes44hVZl0iYyDRmtN3/YX4RWq9Esmh6ou0bfCFdP2eX2p9Qvfwq3EaB2TwjaMPfVyHKa28I9IUo
0ASFKAGJy1PHx9wO+eFtG8GKXhj7n3Zj3VjNvDrDc16aASO3MZDMltWhl3T0CrkDm8ZIx9bjVsGH
83GtZWeSVTTJKOinsT+ze8Jj3+x4ihopw0swBz7JXjeN8a4J5kQtefiZe+sZlKI31y+YB3PvjYbA
bYsXOJcFZSelnEnBnKyITzlNSTu61MVbJ6ECYYeX+fDM+21ElxDp66/w8g7Cm+x4lbhbHHxFbRou
xi6ffTbEHc0Qq/jG9ziMZedkjKWNiY9KGWPVoBwGH88cyCWSccTwtw+gxc82b7XhEu3d+/TQk2iB
fO6VsM1dZc0aBXZw3BVShjeKvLYSByh1sWJcX6pXx7ouxfxllWrFnC/gH4MJjCxVTqdArUlfZCI8
38OtE1pEzNP5qyfRV+H73atoplAfNFRmkQfy4AgScgJ82wsm09nPZ7icAF5qEyPPahk6NJoDwb2u
sKBPzD7Ki4i3OuzYxZ9twYcXd+SPC4oVW7NKl1r/XVd39pG9WrbCi3WwcIRZeC2zG0sjnxy7u9TD
BIHvNf0QamovNUSo85ek80OX38ne58M0vGawC44+E7hu4hTh2dg2ZntikQpuOW+zP4uMyMY1ABlF
gscc5ZyN2GOpnhw/4ipUdEAg4ImQ8XHO4NoacP4nHwhC5Cpf1SRg2An0z3KrNDegCpIquXtwI7Xb
ox+j3yAR4L1Q8eFd1qzRT+gQW20plTgQFFs6gLlx/IzmzLVzru3A6Ws+rFmV/CYCPDHOjMWBJ4cH
r/qt8SdeUzVXOCBKh6p6rG+QnyJaY7yAPxJRq2Cpu0Zrns9iPQxe/YttjwV5AtNuGMyVJrSQ3yPE
JSqgFAwFDmKBkJDlvY+LuD+jY2L4Hl+KNZZWg0sqL69jqY5ck0//TE6yEzBFCQluaLp9BHK34hy+
ZW3NNUhv43jZSlUMYgTsFC9wYQ39RPM2H1TdxNcBp4CZXkZiiHgcb+KglzQdE+kkIXyr1iVmAR9t
9/rsZwBRR04ADQlMrJ+jFYecR9LYO/mLDe6pTv8P4sKIgjPrMQtW40MZxGzVn14cSJGmhTlA12bk
Cd3nD/d7WHCjHREXnE7cuQ6z9OBVPLEQnSVmNMPVKUnatDxuvcfSF978LmhbrxA40cK/p1j7+LbG
biiUTPqpZYET5nzpdc6h6ZtLgXJQSduWj7nK6GC1YSXfoJUdwUmC0/2nMPKYxMAiCnseSzmwJNap
xuRCSatwk0HuXlwip6xqGWUCkU4WEn2gZzXjU/pJV7SqbwGOom+z55AWC5lelQP97XkbqekB3gzC
ov1EvMzM0i970CsCE2rymPOu1EtRDaTRkS0uMX1+PlN+DxFYQpRL/h04F1auqrMoncJJGer6Rjoj
d3kb0nKomX3mQFA/PcktVMBQ0lRTHI+Q5P6XTUnygh5KX6ZACtrkAhurkoKm4KFKAZzFCcDBxrNL
MVr6BiQfe0iskb1XOmtjSNj7k/x93LDWuG/w8QwCfc9ObWT+bU3cDvw1OYFZ1EC/7jML3zQ8+dAA
GqmRo4jhC/3PizKV638maV6vhRH/ZjBgyLIrlcA5bmneHjWNEzoequiGV/Pb/0fGDcqyxEYZdIiZ
ZMALggTXp+m9YcRHayscL1DKEMS3ngBaqwcR63p0BKiwqPeFbSrJCKFwF/zTph8tbV5RlxkEuuFX
5nNZuYpXxThtNqCx7Kw4SOzVevDjKXl+G9Sk1leWhdNH8A81kfsjn1POKON6ys2aQus34024ZJr2
zNvwry5xhBCAinoqrroa5x3ifcqXfwgTaSeqBmWiIB9QieuUtP2jXFOQ2qRHKWz0kBDz9r1WcD2F
bSHg8Uh2bcrAwgrOPmN+/uKYEtNGK+3D3HrHKCnPe73IAzKndLdklZXyeA2guizvHJy1NEYJFYGq
lEqit3jDes/wc6JA3Md5U1Xwf60yDKCm/RdIcd/n+9UJDOChqc6wsw/pxEPW+ivUEdjTWLR4GgW4
OaSGBXFNSCnRBLzhWz5jOExEpcLBv7s37Wik+PO85YFOZhZvNDHR+MX4E3bFXXB0yudN41Nhrlc5
QcIatHz85y6HXZKOZDxW5BEB2L4t7AQdhCDKQplFsYDZikzeN9DbG0KfjaH9JOE3yQunntwohKz8
U6bL2CizIe8OMdKHWwnP9QJ6qtD2vXYbcmN0ZoJiahwg1NB6A7iHCb3FhlsVX6T+ZqGTKI6UjbrH
1W1I7OLGW12GXSrU6AA3kQhsNT8LQCuOKOFZPR+MFdLLhaRvyRKWaVaJunsLe/7jm8vaHjq2zf96
VrY8HWa0s4N5+Brb1cP09s6nG/u+vsus/dWSSmmG8NAtgRIbUBN6zKLydMcES/HqgSPIS1uOOHHD
tWTerVbraiCMOfjcDBarVtFn7n1gFS4aH28RhFLLEtmtlEc7I9j17p9BaUqkGsQSrJNWIKEW6Xde
Bi1/VNm3pavtMynWPnC4RJHYM2qy7vKSxvBbWI/TxtUD7pj+R8fYMiVqQZrt/dKv3hVc18Xj2RmY
LFN7lhC6OxSugjaGFlQtSIsj5M49IH0jmqKAcQz1MQzBoysEpkQBnE0vr8/e7s2+aNHIUPNqr9iW
7wIgui99miwMtI7o8rTOzoBVW4sJ5qztsuh+fmLdL2iQM6oFtFHVG42CFNMoVSMZLh7FBW3odC2i
mlF7YzVLcSgSoSEUE41ihvuP3d0S8qzzkCdcT67eOv7xTgPnSYcHBtiaH5aY9lNwzgX9A14CigeL
5JHO3MeHPOsTn7bGlcb85PTgITOmufb5nbgvf5ZnXrcr3HLVQKNupkEVlXTgZEW+9L9IpfCk+6FD
a3dpFSuGG3G4CA2Ol5YJmLxCUS/BSxJH2Rw3fv00v7rUIeO7wjQxv5QcZ/E0o8SeyBu/qoOQ0COP
2bXRhtVd92lQO1m9YyWnhb3dQHyLhGj8loic1zwuStZ4Oytlg7fHx12Csroo1BE9dyFtuRSC8doz
i2vaQC2AfhycImBTxci6MjWRunLckbA2ZJONYECm9sQxiCfn4bhEhh/nWMX3rkIg1+HeMnLD8p7E
jY/S6HvAcwCRriJaf4UK/X23eqhey/GRw/V7GTEYg73q0WmrzusgKGJgnFoou2C1LPqrNqhNf5KY
6xRGwKtqTJO6skKg97hRleqO7ZRKQy5kIO+QO6Q+ff9kkrnRJCzATGNDToynUcE+C13yt6fPvoMv
02WhEBcLskMmyYC6L1tDdIZRxVZYuOMaz8ZWRUTsCoNiasVeliKrtrX0FMe4B1bcFoaGEP+vBWxb
hC06lyN3Pt9Yqx4Z6biZjUPjv5aeA38VvbelV4qSKnEJ/D41qcziles74vXC8eZxEsmAUURYMucB
2hWqYNe/Rs476izD5LH/ypnZNKx1s5pq4102q3rYgum9v87iCliCEqV8xWOJ/bXXRXz9N37Is+uO
61nd5f/JspenvXddk5AWAwRpq6nb5z86hb5sNpzoua/JjIDwVNJuk9szWFTJcJ6QEHXO1vYI4023
y1caFx8B2pXxVd9xjIwcNFZzxh2e9SMUx62sOtnUxcbcD/amVC8Gj5XijVQAi9lru704vSdIkv4n
w0uRVaniUq8bXstK1pqBUKFRYmtZ7n1wSkuFlIBlV5WzLTuZrMLkUxwKn+XASefRCGrqSFDfjltA
TnPG4/S891F9wtXl1lhyZXVwk0zQh9vUsyDRu2rrYRs2qT8kGuGyEtpWh+AjSW9+39VxgIVgmWFO
Ek3l2AYmNag2Q++Ou3MT1pA9gkwmzOfceULI7okVl8S3D52T9TAfgas9G6n+KtCXyo8ujrLN8pps
zh16/n4g64zObH+OBK5KoxxGVx+uJHVi782efgAVgy2P78RsZBOkQkhcWcwhTzj/R+Rf386Ap5ER
UDYRI+PMHl9CuXZAfaN7ututZf5ol6FbGivRiwK9HDYXJdjzp8rAth3AF5gCIRIIGnmRAJqJtMfU
d81J0gwBQtNaVcQfOabwTPqoaV6vlvbOlCzooZ/Syj9tBn6JL8eC0EwZiiFbs3OzUIYe3fvCNqNX
rdcRIZCuqH7pkaj7RZ0kGkmAP3Nqe3xKODWRJYEFjsQkfsfsyXVvwWCgqKBuzoglMg0yMmvv1Cpd
D7ZWa7LZ9HHKhhE4/tuuLC3xYrSOxdMnlPPtPn7CpdryBC0RWjhiVUHO/Ows/IM+G1MOhvQYx5Y1
TKgfW7G8e+AxmtC4UMF7Z8btV+hDZIGKRNTucf9rMUC56puMAnLBjMCt/zLkY6ckAqqlGdxy/ZIg
iM/IOLquJXrkZGW3Q8nXG2OI8KaXFWUaAbwjGgN7s5qriNwEhadtOhltaBgZi77vG/mCHARUyMbw
4cCFXCHmOoVsM9Q/UD46SAEq25+RGEzobiC9Y6x35oR+jT673+kGtWMKbok8XqZnp51D/Bz+KKIR
E/tI2YuLlt17xMFMs9D48QF8yEszoW5ch6n+HArLSEAVB2e2GmwB1+DkvYcf2Vhwg/4mNDgzXtzE
ZS8RhRikSFgTcsZwc1knxiMwSH+PK1MwUCYmZmiM+P02KLlHyxe/LE7loSmy3B2M1ltf43JXpaVJ
Ytzt9NAZND7yBQvUly/mjulC0iaKVrvh/kfPeSwhwDUgn8zjcZqQGjFhttQ6Pc2s02bIvIgsFd9v
tfJv4Rk4CrmmUFLnofmGP//qpgJpgl/fDkhdba0UMQSxrm8NMuRDbshC8z5q/+tEUQJYYcDL01Og
OCnaC6NkheK9p23r5/b15O0mmFMu+6g5emnPMiROpG3RqF2hkfA0jGjUD7VMXlxFg8cSbvPECk5s
qDKocdSDGvgAmJwA316gPsqiH+uhFKD9gdxvLvlUzlAOZ86fJAGq44Ysr2cyp9PaYJhxUsJyEvVO
xNdHMoyOEVeq/aUGszl6WoV7+3w9nRvC/KEgVejR+eIgcyNBNyicWrT0y5UhCRs2zoe+/D+mwleM
GYek6T8tM944meEohWh22s3G1R92DSbTbkBZ2FUlyMshGW+HRk0xwt5pFro73QLkjlBueWgiJ9Ic
PeVioi1lCEN+I42bzXVVY05k2bF+E9ZkM81YVE4qzn8mgYT91BIetFeihtiQRTFBVXua5x96clP7
h/tQSF8SZwL1as/cotP2lua7HmzQHFj3jt7vwyqFtuDAs51k38i+AzILsx5fnh3ht+Loe/4XYZNq
1/z7Tmgn85Qw4/Alk68YEVJNo4QTX499ebqY0N3az+DcaQklU0sNoDFxpEOfKdg/AJ2ysq2MOKK+
bIDGE5j5w6mQOmXKt7R0s/eOq3fZvD6OrTaWuatNvCWIUY43nsNSTMQTAmSD5yFaN7BXP3T21DE0
L+LXmV6VC2ajjQZJia0EVXtGTdiwoeL1MYJkG61ep5F68tWRy3LekgaHvFy5zgHIbSC3Hk6AOLLF
lKb3HGc9nEqF3gCrIwXmCTwGXitoxp4GxmrMArPrJT/meqj3i/u9Q0xoqfGZeevMDmJV+6FZoHt2
sWYc8wgOXQsmhjb2snm3WuSNYoMST2raErZn1Y9ryjE69YgsVcwKhXyYqpv9GHscgeZpVaXcd3x0
AVtg7U8e4QhvKLBzu7u8agnJod0/istsHrCgGW83R62KZaR8+W1OHZnqazMhIi1IHkemXmmW5umE
oTCzk/HjGKCqoOEx9Fl40rZUosJnVRuA3F+dWnjgTCgfrTz0bJT7ks+MRzkzd9qWGLECOBQSdZ20
ckgvBDFb19hOnuzuStUET2wyH79ckhvlEJj/PL7pXRMeuWq408wYBOF+anOLe96E1itRXSTv/F8Q
L6rYk6AqsKDgftEVaNrW8aY5CXIY/eIm5qD/etah77D/nu9iEHxoXGeYON7XDs6XyvvIf0tvgM/7
wN8NyKfzHDOHL2XUsFnilD9KGVUG5S9uue4kjM1iVtdBsTlTSCQV2/Z8Aa+oMGON7dTE0/JOyRIe
FArPaeZyiBazpLwNHhUwWXdyqwyqOBzyHFIz+1YGIphsKPbVd0Lv9pK6ccXArVp7XGswzw/mAp71
+29TZ2mIBrb1NLadCH8M+zD9dhg2l6fEtvRLaoEYNwFNhbGM9Yb4Rdj+z+NCRiZos0H635VsLGgz
8DYdpz2lATWt1ObD5vXlaQjGZSrbkrLBB2JJHkdBgWX3d8eqU1KNCMzGeRrdM81onh/IbelPGZ1q
rJLf6k39mT77U2sc6bBh+PgVFysIUxgbOB0AC2d+EGCbUJg0HocfviwQ0o74QhFXDURnRbm3oxTA
p52LIJjj07DjN0YM5T9EMua6ISBzsdby11m1g4NRwgUf40D8IoJr56GmqQ5Rb46JiunFB2ek94U2
eYGJB5MTcVyGoJRqAv/nBjYbl3BzXxJLKLf4EjONEyZLb/ukVial6oFl+Sq4YA7uDATYbcwNyht0
K3NRuXTkTy/notzQeY3P6cA4fthRtslokFlCTcRFX6swerY/KKfvw9W1exFMkGe1QqwX1DWKmxaB
F9lRQPhB4+QL0gkuRvzaN3MT3QCfLFrZcqXqjo8lE4s1ZHi6W62vAAp7hA4TthQSIwOpRhVqnmPk
46bTF/RydObPvuCxKzB3Z6YWIO8ezaMTQNRpP2mY44+CSetc6mGGjHDhFzbzICMt6tanVcGwSF6M
QrsG6UOJiTq8eKrbiM5ukJf+dTjsXX/yTjy2sYoF2K4hKGXxjQep2u0IfLV7Im9s6LUGLDxHF7wz
EwRouLxD2EvmS0AIwJ4KjWbkmNtkalmdbraTkNNHPMl948LMntnqfWF3k5+3BYjNIYq3P3cuBX0B
HkZX3FmSZGy90WRxytZB+ND6f1KnPabhfIP8ZU/1qudDy2mtPtUaJxe8LBW2J5oUJ16m/oCo+p3r
2DsrRYseD+ICNysDV55Q9O+31ZC6r4Y8pEKWAjXdp3ed36R+JNhq/o2tETPIoWeE/A+MxvjSSn/F
9Pzjlxma+QK53MvG43//QKoKsS+iNopkGjHmx6A1qQJLiyA5BKLcbWkydYhOfb4yTkCzl96dr3Ah
bk5vI9CsvoLw7y/l7poX3JtxZYVZuQ+kc9YFVDhT5edCFCHK5Di5x680jE8uhjeGibvNhkgQp5ro
FBnOpbxXx/+FscKCb60jiTAYHkRDxqFPCAqx2XYWaq0xUDfmu3Cyhqf+eQEX//oaIceIWUyrJ3OM
Esu4PP0eG3KnmN2kYFCS1eUrDg1IrNulqmHsCM5QP+L+R3TTs/RRfgbT88cYtKMJJWVH+0AINRKo
8VXjylYqxwGg2aO708D/jv941YsqB1BEjlfdd4/CFuJUT0vNQpX1MQqNdNaX1rNQ2jsAdAMI/mqz
pX94usPje9tve6VZS/ghXzXlLwf+SJ+hmlX/N66jPCum9to8PceMs8QXRY45dS01gFJorP97bxPZ
XoGDGOsqa9sAzbBNWq35TPXTDwcq7T582rD9ySAevmGTFtWx6R5e9jrYQS7zeMEOPG0tqZRuI0IF
SesoWNONOt3OdDFmucu5Rqs646wYnzJ3TJeBCZPiJxiIXZ6NfJ3hhxCvQZb9WOhVftgdvPOuYc4x
NYLFVkHWIklJ9dz0TGVaft+vgN7rZWZlZ+T8+/VH/PxfmHRFCxIjY6hhyjxm9OwJO1bIlBEGNrP0
83uFq2LZcWsrLg7ISqo0P82zKr56yS6YN/84NuW1e2AwSqFI3AiwXi+61QujKIsikBZRhWVYZbQx
9m8C/YbN4o6StLlSQv+5qQWsnM4sTCwCLDx7ZcxZmvfnrJnnMN/dmucaUjVYny0fujo/rU2jt1b1
kWMIKvwu4+r6Qd72YKXCkWc3oZZCiIKaY3Ib347wWsb1+XsTCImdLBeg4Xhre6XQdaoJ1VymA6pH
6Go14kCqVHMomAGZ8OXYMoN8n/erp/fd7J2lAze6MyTJ1gKX5toU3kZ0uzgc+eUHW0Q1hP7Xv3Vy
yKe6egDCXsQaDVljBgOXyQYoj3oe8TA1smVE3F5VA2lkLDKIQtEoU3uzwRHMa+OzGsbtEW7NDl21
MqWEbxfCeAXSzPOiqG5Ll3pdG0RVl3vapRcfiaIWKOrjo+ceNM1k8Kzr1eFtGhqNvPGFtVTLXUvr
707jJKK+v7mlEmQ4TXhYcMU+YRSEOPxHGF1fxNa2QEcTaZng/+hs+h3jkTvK5o51Od1qU2xa8koj
VIUwfRTrZy0U/2kp8Mm6Vxe8xRb2GER56SbubKHeEXgZyqyI5Ria0l124dojnJD46Slg++eDOWQJ
JaKNJc31i06rpdFLXtSbPcMak0r+4K/SJU7XGyMViSKbNintblazarrulHD9KfhKjtKz/DjWnqHr
w7z8mia8W9FpTTb11Zdc+JtzIABSIpih5Fzylo4fj6TlctbLcz1Z4nZ547NuXbLDMPRbpxXObaGT
lUIbbK0/Q+kJ6n1GA/J+Hoc6kA2VI58etXAIFSSp7DAoQmXkSyf2966mWfMuZBuB+mY7dfhr+h0q
JthPOEOnGNibQtjC6nxo3qEysmFkvSfO+NtUg1MBne4kAt/e6nHpgpr62gIt+kPxJiCrA+ifZdwN
EuRel8pUv0Q7uGSW82qpGi/NH/xqIpf6pq180voUjNlUdaYRDmZx+mClTx3lmQiBlRidOBmmXTbH
LLCYjHHUarfhZGjL7L1ZEZW8v5uZJeLZ1YzTPnF9gKQjr/htJ0B6Z8BSi3dvfRVYDLi/fHkTPdsM
bSBexNkkPua2qPIZrMbvgD/7smZejDLc/f41jvgFwva2lPB3R8VAWozBC9+7GyJi5+M0Nk2Ilrpy
z7ArGMxzBpLXejgccnprx7Piczw2pkO4SRBWuprgO12VYweSTc/KbWu92n5C+OfS4hiOoiKlAy7C
/3WZtXZMaCly2kubCFZLacT+OupzU5M+b1LUUSkMWqrc9huZIgxdy5DUKvUWL7BYG5IdCb37i1l8
XwWgpDnF9GjmdDkDg071UKP2otJ1X2dpM6fJq0QiIGGlmH88ifniy6PRpKa9XocdCknFmBc0MqCW
a4yBlU9zYmIYiE8wXjwcZIhaUXjHW3cDsPivyq5T/kSnoTcOQGvDl/WazjHng3HjnE6NjLEbXWa1
pAnyRgyl6ebDY7+He6PjhuNMoXNAniebv054oVQr1YE3i0VJ6c8EzhDta0sl1qXr3WxHxTc2WRId
kN3wTISPILcDJUJtqgl2gDHMwN4Sb6yJWdyB7MENFa5NjJclXZj+SlogF6bTmxJjJJ3hVwxFWj9k
v6hKaKkKu6LoJ2znxmMxRuTIhmVQaDPyw7nbGSX5tQOG8HY25mIB5X+SgDzeIuxsRg2wAIhjPF6/
KcfVU9gQC9OlvHU9C0ittJJsMI1WPFdEtGdPXWuA5Bcx6YwEjpzyW50cE3RH2YlOtyy1OYYrSx/E
4HbrAtlhGCqL9hBlwVyENfteEej9lOsylWQhCaUEUH2ZZqI+fbSgf+Yztb0n55LslKa7pVcWhE4K
TwLtK0YYKMGT6eLMp33R9/kf07czRlJEsqHYWdghz+BHabGyPpMx4yXnlkO3Us/6wsSg/Vp6LdD/
IjV2SwQOzQgy3ap7s3vHMQiuxS5gcJrICJRHVraXH+Lp3lQGaLpfEsggujTpm0XIExanfBARgzWz
OiJb4/PZ+105f0aEa+GblAlAvr6cnoPDA6GprieuWP3VHRLa7hSYLkoYaXIC8gwvyRuQP8enXZSx
uc9EFeVSpmX4Gekl58XFMy5UkQpbTftFPeFvkhMgRho7R1bVhWmHPWDJdxqi5RDNIKNmRID+6IRP
Um3ad7TK6ZfYVJIcKIoEjJ76as/85XUty75AqpclgVgxJfUJg3CmMUHGMnn9Im1nXcRfY4BL8Nut
H5cf1nt658y7tRNn7LWkXm3s+LkzkRMGi2BCvOekrnBXpwTvilgbbo/wC24BhcxZ9H2J2AIefgGj
sDA5OVHYih/WixXOUcwJw9oT/vPcRmZiY5c1hHt6hY8pRIxo0qJpv+qw5UZMxR6Os9obOkJ3V6U/
Co/CYxOZYA+OR7D3CruqEjq1/wnCd/fta4tzkr1gEjhu1DLl1m8RTAdmWJXfxmxlHq3VV7p9dI43
RBEIPPYvEN060ZSTdDrMHzfvenybp8wxt+8ENv7umktevkTwrLUkNgiA7odNiIcpTx6b5EPp1tOd
lECiOfRmaHsEcSClXkqTxumcuOL28XiY5XoxddZl2usmNpjgVvjqpqfPQSsKVljGodKDT/zYNTnX
Xpwurz3jF8931QrjdN3uOu/eblRFal/ebzefMDV9SWILVdTG/3dQZbB1LhrXXnEdiG3qVbVi9w8n
3x96W2HiFhYujnu4DzBrCcfV1Py1GhwdnCQhs9mdwUmRr1zghC6Bc4vCmbECTxrRFQzy0oAW1z5d
luWUzb4cH3R/L1tGE4lf3JNbcYMB+T/ZmBpJJFROKLeHCtni7pbVpdNEwMLGq9aB+xrn8+z8M023
tbIAw9QiMtbnLfZFKedn/JMj3WSADVUUTjkF4/Vr52xJ91753DKXdSfjCHj77dZReiJbRbkn7wmk
IS8MScpqIuWqESkRQ0AD17rQtmVI01KFJc92DPH2AY+gPW9zJR5eCAbXeeoNGTGb3CWc01w1v7iR
seAbfhAZ44+02ocQboyyB0v2ebFHcGm2F7yLVH7TVzIw6M2kgHNY38sHAfIhKfgJfVOzIwWPRLFu
TsMbW94IqwhlVf0Jd7zhfI+eL8KQXB7Ay7oEQK5akigsyEIejr7cAJ+YRCPPXUm7NgKUu+0/PaQT
i/Y1KJxNg98b6G3pl+4mQcaf3+j7bFC5o2AAcfIhDhLYY1FsrTPRmtw/85E1qLZLY5JXgX+LRU7S
avpFIlKEO52Ew80d5sjQYu1r7ipbpCTDItyv+Q4K6pk8Y9TUYVEIeox/X6/jEu5FC3sjwsP8B/W0
o6efnXU/8FIP9bU5meiDXpU82s44v5yYWfs6OtcMlvLlrmpQICM5Jbk68eXk4LuttR/E5KITvBLF
fRItx8Yx5KrV9PHaPUkzhBsvh4tOLAMjxpxyDF6GMV8yU6DsZw5XDrGpWnZk0BrREYyWd7gLaj1j
kCE3LZhaPzVrYc0QYSowJkiGFbsKkm3yRSZIJ+ha6iEFSzAQ4NDHcWVfukpYi5s7FMQln4+IHacj
rIZVw7IV6NmAYsg6Cj6/iMkeuVa3PcwCwtJ+SZqxA597j/1v3XQ5foM36dg+px4c4sOV0NvtwcKa
nYh+FG02qDr/E80o43UK+T6afOV/ZbSvnk9D6nH2ZOVqfPEgUgJFg1HDK9vR0PDQ/6pwdgzHOQdL
7/PKd5MwIZYltj8H34MkGIYFY/PTx6AfjyVlhnMCvZLxxaQFA1PgLUAcQQuSAJMtujyae49RDUQU
qkheVnRNocN68DqG17HXe2s+fp8NPTG/92F+DWvP2GQCeUHcWv10TERiOE0xWQRHKFj8jR/3dAU3
Y4aPdNQ2qDRODwoxrOYPjkf3IyZgcupuDyAI9idCoe35bYnJVP8PIPG6wuwPwvDc5bmDWgDj69vl
chsvlAWKv2j9JSLQxNN07sh29QHdezVXjvVshjaCwFGBLc6eHUlm7AQNkcqszkI0iWAF7YxMtgK2
UPZdNDkcJtjs6EFBQTgBnIs/XJE7v289AQnTdJtFL1jltbp4dqvTIQzaVvQ3WmNVWhA0oMJcwaN/
oz+29u4F8ruujnNkncofRbT+JgWkw71BsFy3XwihtBVHHGSOMWDbdzvnPFJaVkVvjpBOAT4YhdT/
to8wB2o49KoOztts+hyuZADYY3XQU5IWNZ2/u86I431nYkt6trrCr7GKAABb30bEPmA0shzveW/t
7RfPk6Q0UAxSyoYOisYTCPyubMV8KqSxvY/nifop/6OERTjpsSx9W5LGr8BvJV8d/HThw1JY58qU
Hakw3+pI7DhC1KsLcmFCrSOsQ7ax91QsGeiEtckSeNp48QK6tarGyj2PC9VV9USaBdxJQ/nUXB/S
EgEmfZeoRz1LAipQ0Q3U+Ab84sW00aq4+t4QGzp/OIijis2hsQlKRT4cT71IKGV1HC6twEuekpzn
5p8pxNvfblYuXDRZrY4kI8Olp8TOvKbXwrutPJ1PQqyrplpJW6eQGIjuqKDk35ZxOLQcAXHhYEbQ
efGWYVc9Eo5LEV21QrFwfM9rwCjjgzwzXLVXM2ySBJJhJdvf+VJ6j0PS+t8nTRW9BoBzMvPmekGb
H5KLFFvGKYSdLnV6uEK+U6MLqxovxS5TRwWzdfTnRT0F9ulD9ZDvyOg/pCjoa36NCLk1c6H/+Nz8
FlipKwKAs1bi60kPhh23PYy333ILsfQ1Oi/d7IPzlmBr5Sx9+gGf4sOED0Fy6PJRUsTXQTkun1s2
OivZnhzQZV1jcpvjoRmW97J99R9KR9PHkFEDJu7Bc9MJY3d9InamQVgeOTKLjmFn/YH3aH0YHy5b
zNqLlAcT5xqYGJo30Jl1W81tQLDcKMS6Ih3Uky8BHO4cDVR9SIltbeNh9Po5oNXWyG2AXZ6OM8HX
d+d7zhFmtWfQQNPDRNJLWtAe3VHMDAxHvM0OL7PWT/4C1YsFsmGcvYeajvQE5IXwELO0yMxwttwH
LD+dYQBoSvVC6SDpA89gXVHRDxKcMEmLHrLO2XED+VsrAYSZe+Sr4Tr6JY1JA0YRMn/pyZmXHqFo
/fuSv3Z99NyYlbxnvZsknce62niOihE+kQ4QvcI3MDlJhmPy88ITTK2yoQn8RzSm264OE9Xsw8Dd
YaMoDJUEldmzi8UNHCmmY4AKa8YqUL2CCGClyJRiOEVbu8hbGMBX2Lxotl4ty31Npph+vJW0ZkCg
Vy6JKfxJwjr6ReJxk/qWhKJ16gpVcKb6pv+3AuzHU9y7e9VU2GdMCQ2GXryzYZ/MC1hKb9wuLwH2
2j1s38L7EG8+mjrDIyJ034hbBAwIevqjUCSH3MM9mAFqX4quJEfRh/YLnvNMIBOGZQe9GwVv5h98
gm1jfhXhZXuEWKny+CIkGSQRqwxmd7AFCpAlg/SvPrC3en89jW1NWvpjRfgp0D6qQWXtADUWabQ/
4UtIgZdjlbk2tJu96DoCrGFUyCoX8UBVwy1DJWuTcXUQgkY2q8J+1H9VuLW9MtOh3vuVN/obiZjA
WZluv9pIamNP2CKXSfcgwq65tZNEUhc0Sfw+1uioR8Gj6uBTdpgyrOMhxG2/UWGmS6vf1M7aadBN
W+krS2w5q3uCJ++Kx+81HD6dSFP0Ke4woAO8nDOWqkZSGKxlLuU92vXModyNf8sK/li+raf4srHT
MiydiP+Rb9299862yl9lsfJFy+rVkmSrQStWcjorrBT2BC+Y4YTuFTsT+E+XuIdU2c+l/16JYvac
YQvBBumh7GZXXPvY1PMaeml24SUoywky1oJcxdP5x5rYnx/TV5ZfXWJjRPZ3jWYQoAhpcy1hvu/3
1j6cJsgFxkltglDA/bIrrBcqEaSsw4Ccam52i/T/7aawf7S3pgPwF8VRxHvmFzAljQoIjcPmoVt4
+Zko/qPyIebK5MpYXwNW9zwyQWtI8FPMl37p4UVF4em4gpVAPa9A+ZFkwakxhl8ZpD6gdCg64PGL
Q7yxKxBVZ0Oh+qTkTPRfn1cwz3DmkOCvmsxX+krbi19Pl3ru7S0RUtF9ZcpJB7xlPA+shCH4UQZ+
+716y5i+ASWPTWWxCs+gHCIoqRzxV3awlZWPeY86lPeHrvn/ypmZWqJpONhET4Uh0BlVDgGgjOa8
527pViEmdpinXTWFy8fb8GapAXkX+dD3nu2CpfEjE7SL5r5qZ7gmcrPhmMdzYRwGD9bB4TDktJj4
A5w/4+rz6IdYfDy/mf5hMnfEnRLezpXB0jUKn+Kdq+BwCg3M0r6zqzg01bqt0y6ohx0JS1Liva+O
3Jzqy76v0lPUv6L/dxJgwq/kpJDGBxsyUHTalrMxKK16f2vIhGLghD9nqjrol1GAT4YhNXSQrY1G
5LxehcD0FNX0Mi4asezFU1hzVaujcHpsExbkIyRiDluWA6UU2TjHzIVuoMqcCkB0IXr3Mjhwid9U
5LYmwwEQxz+yMNiSR+21OGiGwPIVw9utIEkuA4RBp6b7OjA6/fJSZRK/VU/TX1X0SF4IN+CJXA0K
UQHm0JUBQjF485M1l8etdVJCclN3Psd+PiSrEvsPBnpPMsnLhqfagjHTfeCJVglVsyka7oo9hsq5
rsTaV6/iKPczMU7JpBqT3WIVJHfSnBzir5YwQ/0ktPt86uFLGn3dDHpC36PI1OyXItMWN50kWQ+B
g9PaQSZHK0T8HzSJVXSdlrcRUaJPiWCDsowYogWL08kOdykWjDxX2xt3NG6a5RpYrvzHR7qd1bbz
48pF1UXqZpw9T0Sc4WTZlhgq/48rAKwvOz9EqOLRUaUpzECwR7+NE9/wnt3hgVHZUjXHDzEiNIEi
FdhurPR4F9zJ3ifYCb93r55tiJD22HF2BVP4rJn6ALm+9EivFTKszXh+yv6PGBFXueXpOp4wocYW
aCv4deIOZXNZ+h8stJY/FQGH3n2zF31q2+W09TNtGkkgzA9KVyZTqjconQHZboZapIMLv1ee/neT
Rs0W4F/CeAjA+Z+cNeWSpXQo+HkjXHfcpAquf1bqk74qAey7CS+xr5o251alVIewqAq14p/+ZOe0
FoxFrY8wYbxs6qsAAEthKSbIevOEhDLPdZea5Ef9S+f/oke5ZuuwLhiT38myD2m/XMbzMUd1pB90
525us75edZMEG7QBpSthW0TjMBmCEAcRN/njoKDjOMyGLQz8j/cUFhnJITF9KM6rq9ZbmB0VELMR
aWSbkA0HZJ5ViljU7WuEzXjCt5XZxu11tvoaR/Z6erS/usIp4sJsd2u19Kd1ROV6lisChsZzqIwB
1/3/yYiojBSqTcnkUbEIUsjMHfdUpunGDjSI0/ujXMn4vs0zj9ADWTBuXrwRlQxHmpq+2kUuUB3s
LNelPO9ibjF9NW8v8l2O0DOgsGf/D8WWY2F4oHdkyRSUoA62JxOYJbfFW4fHQnvc6V7Xmac/zATD
zCONDlSscWFOXvLv8AFXdBq/ydVqXZugHVxxZDUbm0GBVyfKALrdhDfrbeKZfmmafWWn6u1oWmcw
qfAqexwP5Kbsv+W/gqhW1ah3WJpvLixFitPLL0wMDqzhuUQLbVxoY/Bhng9DhTPp3Q51dxKZ+NxK
w93FuzLt3PJOqKmxLLStEUnp0H9HJOW+9szdR1lD1zvdFRN9puic0kEdY3AP1zvxKbxdXnl5RwPl
NdfZwpVFZtIzzjH2hNfB6CzkofCeYQx8VnX7qsR1/aQZG8TsUFaEmvkI5WgldFuIFbAsjbE524kV
32IWgNgHpUyxhrdZ2csirDUkAgrPGUg986vSudcpejecUhyLcCPd9C5wcFQdZFesWzYYFoC2Q6iL
BiHSUAziH6kqkzA+s9LOn8zuUjP8JrVYzGmG/AG74z2iNE/SZR4oripIpST72hf0/jY7VaDvgpc4
0DhrVegxkbI2fmEt432D7itC57nNSTRou0mMbpE9JZiU2nUxEPVTCaS1bXuXtiwiM8EBCK04jgnz
AvFEtRzr34X+EC/0ex7JY+zAcKDMkja8JFzJBpkC7dsJQzL2aEjZgv76ICAttFxhi7Z+qRqed1LD
GrvegifYXphIsahxZB5skabKH6vsEwutb6DtVRjTSZLH5Vz8UlsrV/lntv1zltgMtBCyilH8vcay
9E1Yda/QrUF3XVjeL1+6uzJPtmYAEAqtjNvnMP7jZumrc/r148LgVFPABBUSjsQ3jz9JhFLL/9RD
kJaeb94r3gnNdnU5IGgZbm/A6sJECfETGCp1Ok92+eQECnWsO/720saP5//bkKNdH/beulWsyLDH
5qEg5in0W+s1FnnxzMA3k2vCiPsw6km6HqMOvdMXpjGe/8ir5qAR8uBRFtY4ofnPTkMzuNIvOCad
UmgqPq7q3kBHTUwoGX3aaWiX7oU2GoMBcNeOv9rtGN+OE979GM4LzaK7NU12V5qQmD5EvkVSmGU6
oybRFD0KjTe51wF0oQEMLXcJuXTsXtF/lfMhJ3esUwfg51mYVLtxU8XUoQMQN4ObYPOuqVRCOoS2
mnwDhr88LsjhutP8Nq76f7Y0zF3QPHdeDfi1yUxZJzdpx+SE4wqEMNXUDwFRA71DtacJ7dZBymIV
IxZ1BlToow7l1P9mQeetoDTPwQMZH7SdNNT20Wwmg+WH1+nVlfSLewneFSKtv/NFijGGqbrjfK1g
bwCPm9DSo6tXIShKF6JNktHfuD4U7Gvd/k9SaT5EKcYGDfPKP4NEoK12f7b4jhdiinFOhu33a/He
MGeEMGQXzeR5OYNvBqwDI51F0j9VoadajuHGQJI5bA3gKttdi14pExZsC9gs5ALoTAe7Sw2JkGcD
Uup1baW8c3xS7/ewW3tU1OzYQ5kU0McN1v+Cfq/bural4DcIy1DuofUc5k5IFCPOlE9Cbu+GPYrt
MTGvp6zwdWfoKa9wqobny9JkDrCKsnfEFa9UcfrAhGgLdqnhM8hLz17BJdCXBIfQULpIIK7qA+WY
PwEdwD/Vo0dTp/g5iSblV1sLjMeSTcdwRiv/fQOraHpDWP7GcO6pdXP8u69Fo5wX9mOPgnmiS5ZF
xirDcziW0aAwWV2WgIviod+rGlKaEuk2IrxSrF7Ohq7G/1zOO3nMHsNjsFbNTeD3ORTVccjek2pe
TS2bBkQLKi9kTUTG8hHKrULHkWOKxmaTAviH3H9yLK+6trLpeXxiZ1dEDxBjcGfso7BE/Bymm93U
AIpvtifSjqV5/u74j01DrWTaGfMe4jS0Yha0Mpc2TYxkT3zcyNkEPvC2khomndi17EVTV0td3pcD
psoGxtLptuig1cVK0Gme3F3kfNf73IiID8hVwK3T/bxcuqJlnsy1I0mCmKZBIx5wc775yPkF4D+M
HvERFg==
`protect end_protected
