`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
katCri0yoqpW3+zUv5aiiW69H0EXIXYDC1rz0wATFs3jxeTpUnYp1/4rcAGtL9Dm+bfDTVKP6kPC
3axWrQhgsA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QCA8J6idKASBB0vaCpPEzyzrm9HjCQTbSTfLTYS1qUVRSINF7HoxBsLxEHADIF+GxYJowHlIssF6
UmltpKeCwe4cVf8GPEYcRe4s+KkQY1FrdZQgLBRE4cM3VS/ynt8EPCfPhZV/91Rn62uXIrA1LBZq
elXsGMsNt/l9UvCNdJM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iSt3ihBegRniE4SleLG2CxigzTtYILT1cLTttwvOqlEb8i4uiUK8flSe4xo4wa0c3qWn6YYBOLbf
XfEm5BriZh9NvKgfkscEN2vX4gmpGdm7VhZ4r3C/rwCTSgiwsyLzUcrjh9Yly4eOe3pQoXJGjmFx
pkPvXwhg12dePwnqqD8qo1WZ2ZO9dZ55lceJJRnfmOyvCU+oeCBqCKj6+Y9eYzcCUpzBEi8bM1US
EL3UdGMjK5Unkmt2uOW+gEOQTGsGGhgkvIC6TSIO7nt1oo0JXhC37alVNkglj4OHuRxFEunGnVRp
CwCvZMZlsBY3s1TLxmnERze62DYxYQ0roDlMtQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Dk0vSc1xKWUAdFGPIT/2WnVUPSVUacHeMdz1UwhUirdniuk4xUNqBfyRlnIaYbHM1L3aLwjhK91x
6+Er+lG+wEr8RiKSY3Z6zUze2mY3jx6UPcWKAIeP84HwdIjTG+d0xMsg5PbvmFzyB7IyIL8mgeo1
N5YxjUH+pQ6v/PvG7SR3VKh/9fIxIpfq1tC5RXhe/w/j2qaryyJsAj2pHVPzV48TmZgDhP2ZCJQO
sYqCdbgeuEImDTC4yOzN5u0Co74BFZ0/RipW1Pp/m1qjr8wYSOfn3TcEipD8WTGfN03K1OVgT/+b
Na5peHVDsa3xmqyfQ4InxO/VTscGZ3ChQZiyBw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oUeLyw6VJGYRB3sHvaA3YNNCqWYv8aOainUgfREyUzP17t1uuHNz2VJPSjtH07/MOUmSCsvTungD
wqc8wyVC/93Xr5ESuq3f9LVUmDiDEP/C6W4lDdMdYrzfD871w1ArE9HyYyHpADEpda7nUDq7ZkSR
JOyy8CEH8ZPh7+4P35tQv/I07DrqN+slOqqE6rpG1mh69Xut0/TBMli2MghYW/eB45yDQD1NLsWG
/bLktNgUiQiOe9ChAKW9iO6uXvFZcv6xxY1s2OKthUMu3F7aNPBv+NEWFIQDzkQ9G8ll+4aawB3J
rESIWKGctdNj7cLyrm8QLMyBAVTwJuJQhvbAAw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e1KYv813kenm5ggS9+C8Kx/Uhbu05ocVcsDBE0RdcS7FQ0IEwiBSW+djBiINubQFO53JMM9f4l53
LBhrpApMBwzD5TaiXksN8hOUXAfIFnygHAftsJQop+rKxwGae9hxfU4/ux5mMO0sfeJr3f4ovODx
2wEZO74s/us57Gx7p5I=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RA4XmB9hm4049EmVNgz0AZh30NFgURwVqeKEIUL13sBA+J1xz+pOMSaKnqnhfzPaQvcesw8+v4z6
UKo7O9Ct72FTX51PHi3Za6DnYnpsya1I8gwGPQQ8975LAXAU+SK/voZZkI2EUI88ZylTZsPTnSE/
MIAUf8d/neDBnilxMfBYdLuqSMLI/dNuihLwjoECNTqxgNF2zMYN/EymjX3ff5Tdr63RdltlPpjp
0zCJLN3tqAk5bqJV0ysVbMVJV8em20CSdyGFVod9KozpbXw/XIbc6aroDHLrMnTeNv7KqG4WKbNs
DFLfWbg9KC3c/0weKk+P2TVbMHk0A0aM56IJeQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 681296)
`protect data_block
XoYAu+Du9ilYpKMZHT5GqWZKVs9xzbK+ylrYNI8TbTvJMOFShxYQ8opCxssUxUQwejHLFcb/yMJ0
lRsU8eFraV1we8beBVlSTDBD7PW0eX8S0Q9KbdWbATnwCJwbp6qyT197G51VFsudF0uslkw/tBYQ
rubaPq8kQ9GZ++3Hw+MMODxiCtyL1p1nHvZfXWJo/PuqHmTfHK3cTMYFhMZu3St0Bm4q8Vo14/Lb
n9UQElt1LLkJ4p7QLwa4KyqJTx1qz3JLovmM1+hms138cOtFsElLjX47xY4cyU1kAVxDRSHHsUGi
UX0yCmSAS/0StE8ZWtFCLzCOvjA/o3fCfmDwzS0mmjweKZbl1/i0drpDNM7yAJ/Z/Cx3tCrwIcLP
nWPviySQsaOCKaj0yr6A8tCZ0pWbF1Q3e3bsymoZ/XGsXjbQvPOhP0K0d/juPknB3u9ko82sOGLp
g7FHlyZb2CNT3VbROusGMPn6zUnSBb94G+wkL0VKJgEn3VWgZ0Un9lsEEkZHa/XR6ZreZah6VjV7
8ZfFKFgZP7iwdozDA5NdHy2unZwe58ynAvHdqZoBeeV3M7qEgBDZd7UQkXP1Afw1mkPdneSUQ7jK
5z+k07y9aRNkhFH6WuHFrLBp0zjz+XmEj6QP93ThN6Z1U7bq20dPXgFayXAw80n95u46QVJxttv0
ghofYWvpLkocD68VaSKPUGENwTxBIL0NeO27GXFFRhSr9U3WSHb6NbEASNNlwqyX99etZ2ib8lGU
2iVBbcTsKxo/OIF1wtrQnQ+RorLFMsOpsMHncRIsSjnwEkOUnC0dnHeXc3IEKCQVLZn8GPqqINyY
eHUbIwE6CYr50EzUHoEn4B9MffEbpPXWS8G47wkQRJ2FT0ztiJ8wFib+68740hKrzpmzD1G7cf4F
s7h1J9aHofSyNS6FepJzwZYPgDxZu3h9ZgiH+FSjytIzjgMa/F4GCFfKvJxp3Cs5Q5a01OeY4ZXa
xjNLT8nbEbJfcjJd06BQDuvvpxZJJCZUfVN2ejhMBK1MCNrosCYFtYLYbWdMphClf9+Rtk3zl0NL
gZXXus2qZ/ISMp3jLscckCZ+cX+LgKpxipdUv/N1k3NtH3I1Aoi9thvp7oFSgvlK3tDglIP6Kp+6
1wVO42KfXrz5kRtytOW28xuGKzb3raXjNk+ZuJ8tCtDyme4T5udfsq3Biu6fNlTkuZLqHe1i39kC
qoyZQ+0rSBJWwUnktPx2AwLw4cWuDcJg33a95vH6xJobtfinZWw+pHQyyuxLK8n+x2ZSQnHgp/A8
Sxlk9HHHZgqngHxkjaaZWQMmuasu+7FpOjfRQXJXcSALArO0JNUJSHiPHi/EwS07I4m9jNSIDCfR
oVSN/MsGHtinju7o/rOWYt7KuNwamvy5WBvUj1NhWgE/5kCQ8XKODCBH0+tTsgc5M+9fPzIrMWfR
pibnTfs+NK4H5t+03/yZ2P0KwTX0zejVF3SGnrdx83wahdHV5lcTIC1/OQXOooYdMXZw0Obj2VFW
t4SiEOCvVkjlLdgf68yS6ptOd1Q2EL4pLW40X+sjnzBJ7OKRhW4qtXbznkMywkfBmjY81ZCErtjk
qWLYYYJindr2qSydeu7ZaYuCvnAKwt5GvblWdeyfoSfbd0yk7iWbUOYIkxdq9V6lvEBUKa2jZ3dz
JMyug2WSRE1F7e5c+tFYzP7+LJr7OAIgOhOH/xph+I67amM8g6bdojKG8zZujoFesrKx7UYp95cz
475syXxt8I30u2e7v9dXODeBiYQu3xH2gvsHRQxVbIuWSBbsEumx7q1kVzYoyosHgCtKCSBB82Go
um9C+y2WfV9Zf+F8K30VvMzcMnv2d0TgpIrmB6vsE3hKSPfV0fgJ2gSfstykjAEMM/F0xKtJom6W
TRc81Zlj4cy9j4gBimhI1TRihiBji6ArhkQgAn65CKLh4Tq2ERMSrfMrpXzNAbWWtkjTath32F1r
F40bmAMvwf0A9LwYK62Lme6b0q8RQCypsJH34z2YfX9vMCX8A1g8FwUPKoDZ7CSJf/q8iewK8ryz
p3sSuvx23Z1bHhgjHMJ8ihjwWOMqZ+YccLOPpolKdnKlp8UY9nKPdm7blzUnzncmLe1t9UJPizNn
64XNb79Xn/CMNDf6vkfdLYCcsmZtRPB0PezmC6bUU7xqzzNB4gbJxkWnhTMuK4a7G9/vi4H8Sc6n
Si/LIB5EAlqXR8yj3GKF0Lz0M1oCxFxJQlH5gXtfTiOWzWt3Pr6261Mw3hOgFkS9IhA9hJi1z62X
Gamzafl5XosFAANcYTYEk+/vCR64zVGAqq/X7bfYD4Z4m05meVMcKQ+nrV/6+23JfSPZZWCvtl9p
BI37QCW2OyECogRnRb3N8d4WJZAes+3grmSc+mH8jiXLybP65z0olvEa8ox45RTKuK39+okqGyuc
GL2/XTEzxk19Xfp06xi6HQcuAyqZpekMnqF+TnimBKYoUMa8TTg1gFY60lKyELmeIjVV2n84BfKX
/LbBHzEuoqNKxh76swl6zYxzyDUeDnzDX1N/yXMWwhC0RiAN+jZ1oncUbJSvJ8AOpdkEaWMcIRCw
8xPU8Wm1SYKv1y+lnDpeWK0X5KYwsBWjMsxpVmfiVR0CV8ggrBsgNImcYOVlEg9KE8wjV2Ph8gwL
CP2ZrGc0UUnEwX+iK6EPAkVpXwY5tnuIen2EmV1MwpjMO+PFMGvI4iuGB22noIBt1NLFvRVd9gay
Mg4GaMUF/PHCmEPYKIwWStCPU93drzkClt0XFCJaLsuzl7oHl8xMNA9mnp9v2EoxKZRGkMFLSOqE
qjkuZy5w/b1+7zBVKBcv68vZ+U4WO+WCiZOit+VYdmFcsUs6Stnv+VS8R8O0Mbk9II0D8i/jUfBQ
wPUoHJ/5ZmurQLgRTZSQRWgOOwKEB63B7iiRWYRiFgeaSXRlo7Um+Tsy1EQc3EO4dSzthf4ffAnl
6wNkGH/lm+VI603zzz+U/GhefDvQWyTUhp6pY4y5z/SBS1IVukKNsOCBJOG8PstOH/LNeUoXKa0L
RIykm4Vu0vN5EyDYFxra+uTyEPuSV37vsgGiQBggqil9u+8Dn/98wo40kPKybZlWOexjJAv6Z2n1
uMSwgWJSoWK9qrL03pofz6CdEQ3uzINhOq95oH7EmlZ8PHrPWlY1MlcU9xZmS19/MPXpWoN97dyo
Af3+akHgXoeeYMbPJYco6yeSRqA2i2Ltp9rbiF0C5WlJxxPw1UIjkpxp8ZFotzWg1ksWzRCfpyxH
F0qDy5KMWnRPZ3dztByBl3++EisnAwwlSgEFJOtbZEXBsoeBo/cUlR3/EpYjRmBMsgbuTXSSE/D7
v+CHcuBxu6S+ZGPFfi0TynJFxM2Hx7pe98QZMUWU2B88b4/Rtvy6mAn8O8XU5Rn0hVeOT47pP+OM
lhfqPm7lse9uRpn6LKJzmBxjFg4tz3VMEzAKYl2x9ZCif6pL9W6W/PoZ2MXc5pfiZRM4UdonnlAf
vq94AqESrJrdNWzWCf7U6wfzHCm8F8Oigq8ZqvwR0XSqXOghavupVtJWY0NDcj4zV3JDdyq9YkvA
33ckLybgzzLTvy9lEHtrmYNdkaPW6nks4s9NqXtNf68hu0Sit5w42XYs6yMDBubfle3I+PYNTOIp
1LNIpcd+fJm6kQNzExzHnPN1AmFlSkliUC4r0CmCRmc1rE2y7emU2DtJVNQfFcUfy7q2CKZJeo9L
K/j6rnehDoB34cU2EPYAaGvLd/qolzgVlq3nx5AUxvErxoDz48lk+7ci79+X8UXlDN6DAMqFvviG
puL/khZruHbNudbmpN7R8PcLSLzXLGDMt1FUxHx9SWMTRLPqS/i3ex9K6obNxyV0tG1N35zdFeaQ
GqqmUQypPDGHPfgYYP+bf9I1tuZmFOXlCjgndrqig+GHBoj9nc7+AD5ss21hqHCwegYSnPRh8cfi
Lwbh3d6V3KN18EutM15Pvdg6dR6s+Q9JPxaND2SxP0Hs0HeiDwf1eZb4sRKIBtX+Zt2ReTvbCtvM
fYEtbO0M8OVqJFSUPqnX3M2jagdB3rTTL9kVwz5Uk3teNHG9bB0LFqvMyI1jh9gHRhNvh5Scr1Tv
PXtS8VYzqf/GwJbu+VLw74HhUbX7DqOdbcj8bEl6iZoNkWibaD99GL5GY5eJIRMz+lZv3H3czr9W
qzRH452wolIJBIePBYSNtPMPVG3h8G7mY7lLfVL5XdVdVNNF47vPkfTiEsy8WrHVhR7dDlgUqWXq
p4G6ndpB93kRN8zb7VxsRNYUqtqdm25Q6Hgt/NBc4BCSLifMtj6aQN98e+vIuKTs7nQt5QnD9Y5m
YyHT6Ylp52JpY6p72AFfCtoEkh7rxZcXlhAIAyDCnKOgYJ7/MYOhyg6WmzvfSwuAWrs407oK6qtg
vRmNDNNir2n1niYiw5K5+vWhCkMjBfJ2WcQUKTRWG86w2kGq9Uqa8Zpn3DYfHnJUQ22rpSKUXpzX
ih5rKb8ZidQpMBhCiFtGSjS4jDk0S5WFyHCITHvxFO/9v2dlBUsODnij8agIwawcgZk6EdFNMLEV
YTjGwlo86ckeBH0DulrmqVxI7xoizhc99y3vrxqTqrZ4N1AC+2/hb9CMhmETGAegQIWu3x5t2UR3
/7gN9lEdk8ooEMPpkE0RD0JsKF908YrSegVpNkDzX1ak/0CF6Jb6/RgTZ7ciT4SoTuZl3dDByj59
hOfe85KMI07vyjwbTl1Owr+OI7CqXeB3uM2DhkchPXWtBUQdCHu7oDmlYy/xmtSOhBOOs9f4G0tE
bxqclk5xlAh1co2hg3g9q4G40yI+ebSInIpe74L0QZ9n0QRySwGQJoGXACtclQC7tLq1ltDSd+DY
Mjq6Ug16MAT6FoxwDDNb2dEZSK3WdKA5iLm5uA2FyJDmzfVVQW8LEQLgI2cz0Shl4nqIeEKClrUM
AILOdHKDVpDVYvASPPKMT2XSi6fJK3GMOVHA/dFd0o1qX2oYqBPdRPWOTtnzwYY5CbrrlN9ih0Kp
8UnnLQDowfMfQ5YH2IIaRxROB4NWg+zk62eKVKEbGYzIPjeq/EA4WRJOHfxOGXcTLt7z+QJfo3FP
8od/ngHHRFuGZ6lMRMxvyVdAZAy+aobOManI/yiUPREGGEZNDAzTbdT0EQCJQlnIUKCzEUo5P22Q
bfDhKD/AmSDmN+VNLz0KuWvN1SgDu5ElklJCR8r6LvJJDpes4XuWMiUzniWEjNPSzEoujygvUCvg
W5aFI2WEjtD2GYk+Z+hvVdhSDP/N0qH5wuXoYhTouDjiSDnS1+eC5bnXXPHyUkH/k1GNe45ZxVcY
9tdeG/kq12KxL2rIQgm1yoM4uvlHQiQ/QoAd9YUeMKQnzqoMEcbdqkr4/ApkzoXjP2uwaHns9xIy
REyr/J2i25lbO5Sqx+hsq5fD9laFoHeV1EnSTfPIeQ+3jQ+eyur8GeP29gDyvD1hmEITUBUmB1Tc
VsBGjOl/f/DwLhcc92XJHFWZRuB1cx2uXFx68HbVX0rLPkpDtaYvr6Ad0FO5OUI3RYdHaGWCRqAF
f3z1u+Jrc2Hq607xLLP+n+RABajYbR2VpF32zJCmUacUU/NqM2c5sMXNGX8PlZpUxnz7Gjg3VrKS
ZbS2LuEU/KfQeTsWwcyN+K0YLbsd0NRg0HaOM0HF180JqpuPnY197/GRg1wj1Bww01x73FksUssA
Ng+s9Ul9wHNuNH5FwXLQ146cdgw9MYcT9DnQwYOUiSXrEEXcEjMTB63y9tyUJ8L9HQM2wM8v58RT
G7Gt14u55cdJNZTY3NWuO3VOKLN6x8TaGHr7MD+0P2USeHfpTMRXROGhgSFPqNqNPqzyH9dVyYAP
+spzD2qOYwg8wLTm3b1JUUAFKLUnI/VrQNe+aN9h5yxT1iplAtz6zKbd0zj1OOouKo8GRQ0+TYRd
/Qx/zIiXrwXTyKRpFDNNzU3ukFb2m3YoZv8+1C3yYpDjkh5wIGyhp4DSa29tA+6oVTVDQ4elI/b0
PEroNMi3nv6xZMahMuJ7uGCMlCw9hkBMd5ucnwCRWBVS1Xbq+3VFwG4mqAUK5QPkNRnnvCjKwf1C
JTWBHhsXFsWnFBv92wq52VND/5rCmw+xSk6F+bsnsWEg1Dw3t25mgiBSk2jO0B3xritPyoxm7Orx
juCsaIGpKNFM/SATulH/ljQdunY+5jk5dsz/OIv39Km4tXIiTxE25I0MINvpco57/BnTsPU+iQEi
y3ovkzp/gVwwPey84oYQzO+yE+H9VnUYhpga1204VUqZJX3BAme3Pgj3tk0hk27S4OJVMdVlyymw
Ejw/+LU5Zj8gyiO/3Iw5cx5/YadQtOb6oHzhPHcbkhErqyiKS6tVN/9ldFyA7bov6mnqDN6gC3bS
//aOFtvb+hoQwa7FZAWlJYk0Hywe+4fJCOGx3trZh1rQqSaLX3nm81wyZtopwyXIPJwb2EYHSG76
RB2Lo0u7pLEuRDEJVMLYEdor6HzWN1ccpvmzyKtK0Lomgts1sO9lWla7O0q9fyWZ/s79Qdx5n+sV
arnxL0gDOKE3LtN1FfZNRCIiu0ARXO9ZfEqf5wU2eDwkgVHB9U+wkjcYvXmLomkm9Cda5e9EvSEg
ce91AD/P3SMGd3MJECerMVOcny8phjCGOnahuEoc0y++l50clhionKjj0BzapLD0fFPV7DFrsY1n
poydKz9aUJBf4Q/HgUKI2kzyL2TWqtRYclIIAHZzlWq+FnrvgPcTS2NHjiS83bRtLl7mz6HmYMi6
L0+t92qWMQVrVml8NFo9Go+oN10KGxbTPF7ybhe6l531li4cdfqkJCE5gdv3m25OAgs3I0pUZHPN
wIKNYl2w8jQE5UtW4EfE37sT3wcsae8FTrgdB9n4uGdqDd7G5tpq5u4tMrEEtxEoz1/1o5B9EHAp
f0llIDndzEKoqLKFQ1W3WdYEDNm9HGvqjwZAqROwW843C3+7htpN+rxenpVwuV7j0sfRZWR2ff1v
cSbHHuyfzxik4V6kuAhiNZGQzZ2BiaAS5xwEVdSNf78ZK/r7OuqVZBZXEIWEuUIC9cv1rTYmSdqh
buIiD/9eTDnuH6uKln7ps0uoA7woIFcyLYfEROiuxa1b8zD/EPrjN+gbvqdQOQ+Z4RgQAEzjt6TT
L9k/ibm1MdgIDr19WCCQ6yVAdPdjDXULY2aZETSO7lrp40ss8s1Cma39I0gbZ44YU+e5o5ppY9Ep
BM0+ifGdYoxJckguQ6bLmygDDl7632hwItF7UOsx3fjrls5jtsaG5b67b00VRONMOgj/VIJ4al87
WcdWq3tzCptP1+zIkplJ1ISDtgb3J/rEkDQCCf6J/3tarfUuU3nfU3nydr3YIHdePVhM+V56xukI
pegCWUORZjcLVMvTo33KcSCmd6nJoD3kZUQA4jrKHFBmhd3r8a1HO6PDw8GKO8I6R7CEb1gEQ6fg
D2x3wfre9FqQY6U3y+Q0zIbhMOtETciTWs4yxKScJdcJcf+NDe1cEvJMPQN7EnD1AXnpUIEHyYlo
PeONL5lIuPvFKla0ynFv6rF/NFnO+3JZEuHAPeZv+lUr0VteQToYgwdlAlxmfc/heFRWHIVFDpf0
erfF4l0K5mK4RcpZ8IDZLIyD8lWSUtxa08AzT7uZW6pXsgOZ6R7JG5yinf7NDDu/vJ7B/9ll1PF6
hTJ8TY9+f9GOi1MLn60Mbzoy3DFel7AXXFkRwdWr/yDWE4hSCZ7TYhVLPRblj+aVb0lO6OuQnOLK
9vsPtVZwP0yo6HWm0AfgUtLH2xunEGKpBpS3HT8k4hO3dBVvOSByq/faXDdhPWnwNpvtiJ6WPLnX
QLCyJY0vSLORhs23E/lDWTKr7+Z0JmpXQlzD+5Snz1/JfWxMw9GPlW9hQRqmDenOoFUdthDgF/DZ
scbGf7TPMiX2hOa/qw5GWh5QUDuGzpLfoN4cDbdcIRnaNJMt8GwJQTrPOrQ6u20v5TYQQaGE6kGY
khBToRpALEe+++7tO1/fpHA1Sdx/y8TElzKlAk5FyyEJX88S2H0e7nNAB0/10KdhWyOkd8nbx4FZ
RlU25eNjV/0hgNDsQ8l2tCm7uwpRXWkW+B00b9NoPpfuXqlQ6Zz7SfR7T8ucd19nNnE2LLppNnt3
5w/bVzBnM+ZIrBKE3jxZiDWZUA+J9pO+DBcm1uVHEk8wR+J3BhLyXWeW14VGVKejmr4/MDgKSuI6
EUVpIzT1D1HERiZ3IUE3jqcrYWPW0oZWrxV5rH1z6Utg4emwdFZbS7wHVn9t3iaEDK9UevSKqXON
lLARtuy/23ZE/X2w3QuU2wIOyrpPZVPAebWMAyPHg9QGJzUu7HR3X1/Y3bb9mX4Wla4ZtKL/jvDL
EC3qRMNwr2+ypuhEY3clevXFDeUTC7tW3+MPxdHYWCqnfOeTB0hJct8NmOuwOOLG/ygKWaDiEuZG
tOg6HaZxPeZFe8IapogjKLuHzyqF5edkGRA/QL1YjoH3xNOl40qM/Mh+NgcN40GhN5n27Iqoq3jX
7QR6GGKmcOkiVGd1NmQmXWk166NlQE2QUbsW+Ac6IcruzSVXK8KUMi3skhnC9t0tstdix2/4tVFP
rMM+P6XYytrDDZvnnpqSarzYtNXw0vsg3p+j1fFz8Zg4w0kqmlbqAnZc3yFoq7sKEB55KuxhSR43
Hx2zSIaFj8phOQCkMrYUwmPPCcavfjle2yzjSsF9TRqwZGoZRFtOgb/cRLGnf4plIyxbmbKK4Che
u7Zv94gbl/s6y0+XVcw2Mc5iRy65fzNm/mkMxWqlXUrQDyTQC+H8N1QgrJXKgUCAP/Rn/3JELgWq
TuPaTfEppLHJMKaX4dnyyte3fIB1hya9cnL1hzLFE4D66FTba7xT3Aknow1lLdNHj8Vx5FCpXZnj
mQWokchdvUaMfom1cp/J4QKTh/ky1OmpF8nMuncJDG/jhXSsE8p5YlkIoAXMqMkgNqzfSTP1IHqU
LqWteTGDPh17An488Hf9wrTGtq4zrK3Rd4kc8Fj9uMa7PjtnnAxEwfH41835ZtDgbL9u02GJ+hAi
nvQubvKGDUFXg5D9l/zkfosRckjr6bpACUadVxX1mG7S8/NHbG7rYiS29qMbvLIk5A1Lzc+7h2b7
FP7fQOfRgLLpyfy2ItdelFKfBqkEzva4PU2Cg+QyD/66+MOeCk7d8kLubur0FZ2FDKZyfGwKu9LI
Jx9PP6tteQTDd9KPlJqT/79BS81SqndGyyP2UcrGXTKi6BRUQjpoN2wwTIQxK6dY9q42cXo1gHJP
bvxD/322Zrn65nkR/QkdFRF1NOvBUvQUQW3O1lJdE84oCTG/MQzDCCRcI1ZyA2G2XTvibjKyGbMB
NaE96ZnfacabKhTVCrgjReKoP2wX5+/Mcq3IfcWunzKpegWmWybnPHrq0bHrPsOadt95upli3t9c
9c3HIyKEZouj9yA79osYDgjyapRM3Lm8toGqHlRyKPJhRr7KPJFQH+IEmclQ6Jm18/6UZIplY/MP
HlgxVVnTUJDfKxyPFAKklJlhlgemFduR27qrJEDqyAuU8LXGo9l4utXmNRu2N14XeHVnmq6y/yjR
1Qe8LZorkxZqM8itW2f21iKJQ8Rz0VSLVkTJiFcNZF2s14UxawBsV+d3H5V8Qior0li5JKlJ2otu
nlleJuda05p3eIyJWGYuwzEuufNg7pvpU0pTH4H2ng7vGiVKmfDURb/e9wM07jRhhXsuqZJuV9qD
ttgbvK0d3fZxgYXPK/ffkQNJrNwxNrum65XSgekeKyVe8qApZ7KYQGJiv8bX2AYihueML5N7/4P+
0P2hFXb26jmpCIiOsJJMoYwLr+0cz/qgH6NOEgoL8+7WwPxxgXFYRW5wYFWCp0+HRDnIpSv25prO
WOA7E0axmCTJQbFJo/lQESzPmIYW9lM8lDs84woa1UO++Vw2CKwyxQlSbbMnJTnHtzBSdqSU9jJX
qFOBwV/ewIL2MP+O7o0y4mwYTEkOk5uriH2vtbjBRNe2PoUZTeryJezei6TXA6H7BJiTEG7ITuto
Js6CLaRJeXcfg3Y5X9Qx/7E1a4EpnzgAt8NZBsTZnrSO5v6/2drUC360YKE49a3IgWefZTdgQvza
i7gEkOyzKVk6i4U+x+LGyX55PFpokhBp4TdlSNDBRxUCmBAZyLscxS3WeU5tGDrrNNQ22Ig69v7u
brtwfaYb2rWyh2/XXYr8BnLVSOMO1/dE9OGstQfNSYzQSTvhk6BP3jfk/EWi9aJojdeK8ggZpPJl
i8IrQdH2gstpQha45meJw5I7r6FPjzxzPYFEieE21QUFCX6fam8aBqDLDeUULSa8kTOBmRWnAPL7
tE+ZfxfLjg1X1yaDT4TgKBJPQ5tQhiWpdNEcK9JKmRDBaspBC64crR+kxt5QIG91PDfbq5IsHtH/
OC0DbuRtu/ZRxvRjiYfypyDLzpjIaZpZNm95Pf//Vr4tI0CtLn4p8z8YefLsF3RA+E18vjI46LVi
Wp7a4aAHgDapfRz9+xwlqaJVJsWXw4KXj9GqC6Z2mgEUJpBNIh+CHgxWlcjKwpcDZ4uirDHHC236
RsUnWona3ecWEvjQ5nToooK/GNj29l2hUnuKBSNVmqu3hXpa7pSQayKT6O+CO5Ch9oXQVriT4Wbm
Hadidk0lgH/zL+AWM7U6mo+k1YX0rxU4mvuqiMapL8mS+o7Qzom7o0YDMsCPoCElzqAu/yjuVN38
ip/IJzjcE+vdVPXiG8gN3K5XZ8wIaUQ8PIy4JAExaluNvMntROV7RDsusj8SpXJa9rHuY3wO8hD6
vzXp39SV3zQcWTpxo3M8zx3sqkjBGEEh9w+3ks1+kICcHxl7I+Nso5vL2q8CxuIpSnacJ4ehogiv
WyQa8KGvpXOsQ6T+/ie7uG7VgD38VVXsyNadb8S8YO4bDIGy2ELi+o5lFMHcVx9EZB0Apo+eYs+v
+SVQod0udtxh3NgInxO/pUUTeWNzerRvLfDzoHyiK7E8tDyMfKLgV3NuHI9Hm5U85upDsoMHreF5
lgVAGVYYv5xbB+ivfXCZmLpv5PILJWSRCFH5CY5MPQ8pc5NMBMSVf5mWV7FqT5Twt2J55/mSsQRB
AbvUqfsIz/lsgYuq867Ivt07IK9PkEzU3j14rSb92+qLCT5joVRKfqFjVvvN/0UGEO7MVhduyaAu
YXBeLgPewDD03PtSPMhCXCgQVaVMPSY7xa7S3o/NuL/vnSDemWWBmIFyBevVfheif7MoPicWleyy
4a/Eg5omwFSSWojSc7dGl+qU0nm6Ovhyb3oo7UEmA5oht65V1pEUr5y6uefevuEF1eZQEkT+ui/j
VziwNZ3DGGw9xGVASGxdDADEAVHEM/a2+SEXbboy7scBaeFdJSAXqHmcY4MYJriDgWqm34IskpLo
rabZStc9LTaFK/7gMNb7zhBN0itj06fbg9LEHrJl+0qslmNBYI2g9uxfqQE0PDn53bek4h4fjK3G
KPJ4AZKhPDlR/igsY2bm/MH4lIcbF3zeQr2l5Ats8owbwQgnJrSDyM5vhDO/P0RsFd/8Qj8AV9fI
6HCJ9W5e1dq8sr760AB7iNPAFXzW+5uVCCwNSyAofGWD5j8zIsgzBp/mboX1A5C/G6WbfSw9r0/5
fMsEMaDSSB5KjFL5rKLcy7KFUatqXcBZdl8edNrTKHVcPyHoUhAoLKUDnWJ6rkPX9IhTsY/zAtrq
nqlBYnfTA20MT8WUvxgkjMLf/T0iZERX3JBjdtatJIh01t/LV4qK57xMskkFg4vp55eVyZEz9lqE
F8iWDvMokjofYGG1qcTloQ4YF5X0+SAhTHXLY5q+cc/FLJ0M9zo5uxiLiS9MF8V28zN/dHxUXq7p
r7WoDmKXCrPTz5Nn3ypuGOCQ1m8Q2CT4kZUVRPllNCQLn8/DMdASs9kiMlhetMUjgPsVjGgGB/t/
OkJ3iurPrBgMTM8Df74psLjQRAnJqZRMT97O6pZFSN9VzB4FGbv/YM00RNi/I/clsifgKWsr1Apb
J6dMljq4Fn251Rif4J8rthiQvt34Q4poRdv436szTwL3n0P5O8Xs6xZEIip0z6BSyUyp5yNcjI5y
HH2NZlJbXYWM3go7WiXLsUm5PXb5w6TbDS3MiDuAG0jVWjSEjam0TiqbJw6bW7EZvLVrOqpyytJn
9HoEmfpYyd2M+sq3LJVocR/OctA4vQbKQUMMWfhVVRlT0QKVm+eh0qXRGKzeO8JTKyT2Gwp5kyQp
cNPKjWWXNA+tEixS+dmqj2ktJjsMHnd8jMPcUvgWhI8ChwDVqJi6o8cR7xrc5GeZxI1gseTjeRmi
yzSpJBPq7NpWbGw6NlVeGd2d3ewEUYTRqSHF85sZiGmcdmHOU20P35Tl//KbU4TRKILpMKLbnNcV
ptYuyuGdpA2ozJubyjjYt0C5R1n42w59+7/CTtFTvZJrbkQ5pkVmf5jbiXUVX5AGYWyUwZHjv0AC
aUwR1J2liu/EBGGJ7wxfsDsZQL5qMs6kEDNBYclGy8D+WrytKzKP1RszI21tKXzRcctkTKUn9eQN
otNw+e6TYZ3cKFjNUyLb4l6s6DoQdtoT1Ts3mYe36dz+r7xKm2rG5q47A+LnqhBBBSNWeMjcmUox
dfmnfmV7Zdt2QT0LXqVQsw3wD9q7vBtPTQVKmwSaAhEjiuMDjkyLG1UYf/bqCGoCDxoD140LpnyX
SBZclJntYrgpWYsJJlmmVRV5t7ZyPTLw6fGXgL21rCFj8woYFtuRrrkLSQwmlPr1X18iS1QjPFHH
0mi/ZRUlqczVUadNK8QPb28hebLOqWYRCEAuoVlfRK7R3kYGESkVBpycoM9d6JopRzb4rG1zYD/W
6b/g5WgkaxskSU65RHwQmBDjrC7otmaMOSY9y79+Buaftor9RvNySgv5QEf1MB9lWDerDnYp3v5Q
GRaN47fL/iyZN6dxgMswKDizCynECmrN1ldSO0X+RUpeopI5zG8fWlLZUvP3z6J4Ve7LljIxvuQB
DDhiy1p6Rg6Jl3vOgevXac0wlbh/B+1jhWrhXP0mlBCZpg4ADBSi2nLRQEVfLbvGPaRchDVvQTGW
9dg6HYaZXe0Th+VJHQ4c6V1e/nCGSZ8YE3CFosoktPwbusU90v9YZvhqU/htqQ3vydbjteAse4Hk
ELe5DhVmnVwlxY02RTM3IUTwDw97goeoz5kxM9UdEd449e9P3mhJZCRzlJb9dmZfJzRQWUM/WHgo
+9sFppjLsvPY3E4A5r9Tl5ZnAnR/p2U0/oLcI9Rh+aZhqcXSwwmTZd5uP1Jl4/6P5IEB6HBhijeI
aABRlFPaHqAdVI9RfHF2sDfhbm6LIQW38/2GqahujDTtj7kq7h9ToKligKj66x4dFzbNolG17KOc
61twvwFZaY3fxEZPW8ivE/kLc9kPDBC9hfWE5uJn2d0ThUp9IXT664eWW46JspX116OZm+sM2FFr
pgjbjzDEfXdIJVDzTWCuxiMb7FXyyI7j8QyPjLGwdb9a4skD5UYOnRpBgZaOPU3nXZLa4eHcnYIt
QXoH59yXAGX8bwrJPbWpufd+pjmk2ZhIjf8XvWnH85CoNvZSmohaqJoSOYIpA/i8q0iJKo8t3Oiz
J+4ihvbkcWnmqTusY8rX9RsDAwWCqaf4APk7o1fv8VabSszdqlDFXzF8rUY3/DmEacwnI9h7Vrqo
cYkUef5YzZKn+H6iBd2VGUUixRBbGyGe4LwQ79kMsvlTylXuXjPxh0VISN/359MIIoLkm4179pQc
v/4EGAjkunOASVOfxjZj+ghrGauCLCoMJJcSc7Y/b7GuxBPK+/yrca1/B9AfMRHEovNivxLMb61d
/hVWRUsvIsnrm5FxicPbLBg092mf642qi+Bp2UbafdufsfSH8EIGjrKlJ0r4pi55lq5YrEmgAv9x
YGKWonkwjhggAc2X/TomAn4GGBtdLPknHMtl2GvE/RQZT21hKuZ98K2uGXoI5eYmt7MgDQO1M6SS
YvKEyhYEL7IwxF4fqmTMPqu43n6yCsLl5iK2RHWYaPPuvErANc8BsxrHPFxsMQtI5XSqRtk7SB+y
seF9m+RLn+TNjStKWItcBcmIXsjfLq4aS6Gnh0vwG9plymxRBRy/UJwKSsD/mgzOjb1xTk2nsiHv
QEzKOHVQTJ+N+QSSpUsc7zc64miSg+4cOIbwLbEFH60ZpPbxBEZshMDNaXt45WCwRQp7bczc6vAe
Z2x2nTEzMOFBoOXG/J/vkNWmzo2OCVrVkdSvjvJOB0uf8I1Yo5qgUJ+9Io3272S8+lSjP+SgsY/4
x9UycgeF4EonxhfLOYP8o1hqlv373vaRSiS7cPBPucRuaXI/Y9h/VBWeNWuFAOLGtzPPO6N+t4LK
VwNkyWmaWQXrQyN2szqfZCBIhrYKnM5zadintc0lyF5+AG21jAuKcVeTdrFvBszYDUmNTIdxDLyL
ODLBcCmy5hPBzd7/MVReWMsxeC+hsp9N8wZNBwE3bKd5yyn3Lfij3Njd5VNSIg9DZUCdrWimlJ/D
plQcgKQXTnj56cq1Ngq/beFp+/Ln5XiOlOuNprovOD8TQTmweJFFA/9xKH21DRXyzVVo8k0ZkPm2
hhjmu1X3wzSlfZZOs+peIHFZ2YWyiTKsjwEFZ7LE5qSjmcfAqMsT1SzTMDa2SREGhZrg8gGJ1daW
vUICJAbrpJ4o8EqbZhhuApSugknYcmSySAVo/3C54o7sVmQv57lBKzK4MXI09wCkT3ZBnS5Lingn
zL+wmK8WLYZ1NulwPYFFkaqq1K86p9iTHc3yxa6uogiWRYjiYOQN2+troi0hftFXRP2Qub3oz5PY
Gk5puunjwRjAzBkvgKcjJ3I3KQ9IHj+Nfl6QT/jI1YEBxDWKowkMFyScRRdmdIH8ocPSkTLAmnjv
BLQl9iNdCU4MFbwWBitfHniyb2NB1jkVSE1ZUkDnGz46MA40Z9vz7JyQdnMZWZEm4HFpGqSAJHPy
lmm6zSj/Ed06AcImDaFj5LBFlt95TSFFO3VHljoz28h6K9V1vmGDrDtS3Lum2Ctj3Vnz9Tu+Qtve
vg+vBzeoY0yVlIoV+z2k/E6zZqDqJZ4VOQJPUY531Qz6R9SFw4mBrbXroZNgx+YIB4pVsbkk2PmC
fUpsCF4CIc65Sxr7S/jeZakWiSs8nK0Yg4v0QPCCy1VxIq9PXKmAMGKFPH+7xeiLsMrRNQ8BY54m
sx96qhOmMbn6zxHOmmba1ifbv7qwD6N+vgOJdV66vDzE3tLIYX8k2zCdSdgcO2rR3ihhAMKr404r
O9MJkKZ3uW0C04yEoq/3f59/LqSGMxNka1xGfzjivFbMdMtucqNM6olMInfjsJ7Pz6ZbKd/Wfd50
kh6d7gmjDeTSgmSlviFr7Jv/rusttSf8LUEdKL1YS9ybP6rGTZLi3mjX619GlXJXUyS/L92fv5of
V+MvGnkBcuSWF3TPYEKS7wETEQJzSlLvGzwTSWg27dYajCufptzmj2LxYoNNC/1TwFptHTTJHJXR
ymHH1BWXMMeYZSzvmbIJUBm+eOqus4c4CJ6J/Y8ZJ4SgkAS9ARFs+VNNSYzqAKKm8m/IQxdydj8u
7w9S9eSBaEano4ddsEE8J2IBXJj6A1T1Lzuvo4tHpvsmU7zL7ntxvsr9iXfSp1g0enOxsDNGy/TX
FCvsXxNoz4PhGtniQi6Z2xhtnPFDxq91kzXW09F8KJK5YV91d+zy3xUKrUBtWVWWokZWNH/Wnx+t
jQmWnLTotcmhbprwJDd6/aC4dtSiK3wC/Y0RuCA0nNuR7XouBsF9q7zOc2JYI1y/I53diV+rP8QE
+rUBqu+fFPWkddUQ4K5ANuiYWMUhRNKGg8RflqO97An+CXKykKCPdqpXUlaEZUWqniAdXE5pFHxP
P1JIrqotbVAvR8AGBF6Ah4xgbncn3gda1+GK1WSqrRa9X7dnJr47l/eDQ7nnAP966Py3G44L2W6Y
W0TGSM658AAHHUr2fkhGccix+RX/Qi+aIl2LAMwul9ltAXswrRP+lLVJsPsZFinRbkEkAV4SyfhZ
SwDbw4NcwmpIPniGo/5EcczxiDtc8xHcqAFCkXRJIdDL+4/HFlBhKtRoRbvBbFeB+M4b204MfN8V
TAIkOmeMzuOU0zLu1kzqDATaIA+VkpYvjGIBDaffjA2WUV4mNljcWiDPUfG1XuJ4WTHtG7qxE4jL
epRVua7O9Srs1GrBySjv1YuY5mZ0v4Fx5G9JJOi1uTWYSgSTsaUnJPDAlfxw/S+CncsbCFPgbTbG
2bV6PDghtr3pMcHFeDgK0ElmpNOfxMou5lzzkjYqUPKOePyzUOjO4R6/N6alG1NbhPcrb5lFUyk/
QUPJ5c4RcuakWSV2HUaAHopDX2S/K7d2tnhAh97bmrrWGeen09nmLanYrbnieYIatBjhyzJUgVPU
GzkBxNh2glKrEWKJJXAzcoC6dxrR384zL4dyjlbMmMXqbVxYjmIIvk95GbmnnhrokISR1kb+Bj9M
AKb+YjmcgGsq2bJm5E7Yjw0ZlJox4vIs5tX7dOv/h1XOEu5BzzEX92YbCQnIQt1Q5csEgRBVY6G5
JbazW/Y6c96hrs/PZgxx0zndQvKJmvppCpZ9n7Xss4AxirGr9T5B51UdNuyz0nrcJbEMcJRsXUIA
NrcYdaDD1knjc70YpMcdHOOkTdpednTByizArzU3uykD+HQKnIocYlm7kyeobD2Om8lrv48v75qq
fx5XOza3T+5+5xxWsoibht1dzsqbgTKf8jQVnARGFV3r6RpUPGS2QZB/lVy2qb2lhGGPDflQOU2s
lPCMHNMFl3HESSUAm8Uc3sNoV0ol8HOFnovS7ERdWgv2CJuM2VVXwBS4qLYcNTftARavTAvoCfoK
W0e7plL8FO4xLZyo70+bLyOPPTxeED46dTdXqdgoucaoifdw5xilVNBkneXD8YuJPBrZojjHNb74
ZinIl5S8MIf7kzj6ghLAk57Uw2fzpI7RDfvqPyhg54QzbclMs0pFbrDFGM11197Do94ybgQ8dVND
NmtFC0HUxMa6OHMYj791+dzlZnmBy0aqQ/KCZa3ncZ06pYWhZCUk/qVk49crO7IH5F8XSUKOcH9w
mjpaZipMoV2CtEKx73sSFR11EUFhnSS7HahiGWB0FUnDfu15B6Tv4+DxGfEY2MRw2SSUvemInhaB
c80w0ysfv0YbYcNBanrUR+/WwPC2PlApI4S3l5YkgM8q0N8QhWhYxRNSQLNp2u8dOVLVFgeg16Vz
gFLoFs9W7gFi4A2qxbYX01jqvPkIlok2Z1AIYh1URanfNvImR0nLUZZ/+5HXJMrcExFp8OwH4QBU
q7CymxaDrPVCXG2vG5QGycLcF8PxeiklQ4W4zsD4Of/h/6OwqSAZiYeebfA8PKk0UKO12K/8eeDw
PsvQ/nbxs+KtaIngTANFEDiGFzpBDIxD/vR4EzaMohGOGw9Mu0PEv6bhcFWw+M1GEERfLBvrX3ex
n3qPuXkqbWT+P5MvyLgBcUkTd5SUGgJXvb+nNJMZMeNJBWRLB9T1OFSOcC4om0wfBD3dUBRWzn/B
G0XyPcUBn9iKYR1im2BXh8lLld9/GcbKnGu3QIEz4GK0cWQgxeFAzxHzsdnduyqCQfPx9TTBUck1
m7UdD5xQG/SSY339onMPCszKkd9HRhSCErnfQ+ZPruBVKZg77oTt+G7ATZtGKplQmUYFD8AT17D5
KWnLcCejFK/FfvfNn6gQsskO40Yk9cEixDgaBNTAFNlWutIt0xn1XJjip9kgVxZAoJ7gz2xIXHad
0DPiA5DCMOJhZxnrva78MzVG6SEAM1/7sbIxeRjqG89eQfIgdaMZqK57+qAYRmyaiTc24768Eeum
0GOwXYIHmkIxnhJoHUGPEyw56eIW8woadZakVWQAJZgrU00xRwIBU71myu+RW28gbG9J7zjX3czS
FeJnTY8CfV75S36I7lxAMmOkALR0AirlKLl2jwRu6kccRTfTnsePoXzU7OXrmJ2wk8CZlBxn/VGu
CWqtr4RwBn2Jfc0A10kRtRabN9v89MyGKffUSqR5wiZDhqUexzlBmtd6OQEc/ONNhbbv4EfcDeka
hpqI+nMcU35eN81we7dW5OZZO0diMjM6GcPqAf2dcnvz2lUcIAcBNexxXPaPTezeDZoc/q+ldxRB
fAPVNeeVYv5hYfnW+0l/9pUmr6hhmQsMqKpS+PDeNgrZG5Wty1HlQipNrJpottHy/z2VIs1hiWZS
WtOtiAhBWIY94gS1q6iAkeVRaCTViXcTdGB2AjUwGw62UUSmJv8FJ5B8e0/NhSpPgR7/PHAmK+Ik
zVLZMRMhA17J1q1+qBfGQDkNfIDZfHpzYW7u83QlNlAoh/hm+RjZZ86v1rqxA4857GmXpZgpzHWx
/GXCjg0TN7g1RkiIfvSrM9GLXX4x6fAUHaEVLJ5mxJqq40vH9w3pAxo+C6WVFtflA0YLd8gzNBgm
jAk9eEQGPEhjYd+tQiQAng7mT7/4oOwn3KXgCYQjlUYqisyA0d89ITwRvC/ZhEVI8BcYYsPqHaAw
uBWTzsJcvz5jID2IAnUo6k4CQyik73BU3lQXag51J9p4nPVpGHSRfEuJkORvAL25WFXepe7t9rq/
H2w6YuZa56x27lHkquMrtXGQJvRuLKtvT5ml6T69uO9Ns3oJmfn8HhTQeAER6avNeR9BEoGXfRkM
fUtNz+OtlXHVOFTk7eX2bwY1nLblRcruJSWJrxF2yNAfW/Qpkncl8kgLtrp/Oaj4cvcEBCyfBo6j
6xxswPCpbPJ7b3gz87boy+2NbMfoFFoN9BvMfCQzkLz7ko7uBI3uASGpdIR9A25PMVuY0n42jNQk
A/XDei+w8Mp/J7NewPa+r+5RTH9JVc71DaSMGLmMftxMMRZUlHyNgrvN7VHeSaFMj8p4d3H/uYCx
0pew3BdpJ7rYr3I0I7764WHOueJqGtkIVPp1wnZaL1J8C7/T9GdTfLCx3xfs+Tg98pMEDxoxaFMr
5svUB1uNZAo923t6zCJxIQcqG7Tl0p9F4U7Mxxh/ii+DmxIblkDna+X0jheRam5UeLfSpTxRJeXj
SmQj+Zc6g2AUYSx7fBKCU+xoTrxQqYW3x+wiVO2/bfLZS46zLx6s28YqX3loAJZeBc3QfUz+b/MZ
JziI2/ArpLOwnyumO7q7gNF3/mDJ6tz8EDqi7Vb1jvRNrewvGjvXs44LVEmniZsmj0edzXfekRk2
DH7vyaIRlMIWHA+nM6yrta/pWFodMjCYzeQJuzjvSSv4xhGOx4hUyLZfo6banyLMC5/PQQtmxSZl
ckWCt7WxABAztOFu7ECnfbg6nOFEA8iHN0JrOwiL3R407EsJo5Ha9RkkRmkOmAYch/W6MKy+MZmN
Y5Y9QtvXpOzX5TuzOVjJ3LZtp2AdwU8F8kL5kPWqV03sZ0+2DcaFCF0CRXFJhtdTN4xtE9P6IxpK
1BaepO0Qp7qskrA6Zh9BeiSQRhBHxUVYsGPnSGYYo8vPd4e8EueXLtHb4RZJL8CUfvukhREGMmbK
IIXJixQ4f1HZcKBV9EvuWHAjHXcMIASA8/hvxVKZYNWBFuQhHzghnwFjIZDwjWYWD18oxsxIUjFb
aOLnoYyixGaoOosojXboIOyfIa0Xv6a29SMhwpktTMVcpHCo6AqCiKeHc2gKJ/jxP75wrgVlcnBX
DkOedVP9GmVLiEWhk6tOqIUdVOKQFYcLKzMocXXItBHeFmI4O9wEGpJmF0sikkt9pxhjFmCR6Yy6
clVg32BOcYzF6mWuM1vC89i6OYQ7fTC2C3RqAoNyIHYLJ8H4p8dQsZEc9VDmpd9248+iYY7Qvn0N
EyM1SvWUIuQ6a6Is6ana6y0qhjIFnBBLNNL3m+xRJ8BTQVXI/6X3HkNv/LCLIP/1CvX7a0WxG96I
S34MXPN1BIcS33t4MQtbAq4ljuBjglJtKQMbut5h7A/Qa8eHeiNs3Noetd5pAs1G4L7hbu5WmNU2
TSBaWEmCRvM4o5GJgJxELGt5/M9s7Je6oRQc+l/iNORkiGBP1CeUq9ZngRhTbBJdC0dI+Ro1O+0D
Ph70YvyRloosimVvcMaT0oOjF3JozlpSTHyCnXWdLExlYhq+41tV/XFjmca7pR85UIGi0YMjOfi+
A+890hTmDQUJS8O8xHNTu45WqDqix7q0Zc4KEGvsNH5GcTIj6dzORvBi82WeSlQaLGkH4K6KLtDm
xb0lpJK5abePUlF4I4LMC0ERi6xDN6FNTlaoOMeQcnetESP4fjnHl7cMfZpi7bmzg2YywGdhJ8ba
brXrTNNkC7vn3b+MrMAYod0Je5NsgUck0l6mVploRLAJiyeKtNl2IXymwyZL5/PCnxtj2feVqfkA
ooJA+UoAslUIfBgGNe2wL1HYBE0mjsfB1N7lhygHcpeaNagopXW6V4s0MRAFmB5nr4jtBqmQ7p6R
QK0a1YFj9J42qGotKC1BSu2EjW4xhwdIwvmcK14Mp1j36OHAKFzsqgnX6+1zwQqXp5wnjGZHPVlV
8gmhwzIfgVRQlfWKx5xNvLbD6t+5bqKWRpLTUrmbvYCKuMy2GE2dkO3hkiOiidjzpH2kSF4jCB0J
v3iQX59BB9yERk7oz6VDqb36Nk5ftVd1hrH3CBe1IKx+GpZ4GIaElOwF/0egrGIQ/Z8GFJhdpgoR
OCJOHVVY/VTCRV53hNUe0ovr6PIAGmPQ/V+9+5o1qShYrhQKLai5AwoPdQKQjaBUmiMQrR3LdKY3
2EgEIdk6Jy1ksADN339nGsjgX35Ao79r7q7jTJEGAosomGaatEEJmdXO5cl2PyggjuBHb5m9nLTB
qv5uyTuH9PJ9bILTyarWlnXVnlV5FQkZBgKrgp6nM49HoTIt9mErgfQewuNYb7eHiViSCQpUWN4Z
4waD5vQjhaSLZyau4dFqsW5t7+/nU9HpbKWK2JvypNgK6dvqDGWJClF8l8IEGeCiwEH5WyWMtG2J
ckHUgrPdC8Qmvye7do+ErKqgtSdOg86mZrKjZtc2N6IoO8gPaxAoYOoksP3hhtqEcOdAH9+70uvK
V91SBSkpT2OKHiks1uhIGBvFvg0tQp2x5rhlUrdtPzfWQJAmwyltz6pEmTNrEOQRrbOR1hb4c0G5
4+5w0eHCZfINxpMjIkrTzQBGVhCBy58XC/s2+BLAbVyHEp8eRDlS+UQi+HBlIWfTxP7Zn9egdNHm
sKwkk33+7vy1K8FL3NV2kw05izbqKiU+yR1mqMVu4OUYvbFC7kIq2H1kGrbOIUse74Y+kJkO0y6m
YdQcAuecxVQHXMHnsb8+lT9vThEVTFezBat7X9EibscmLDpilibttgtZnilXHDlFtm2TIm4ZzKSl
7UzWTu4jBaQgpypnN60QzTPBKgXOQyPTLJWDJzWVDxyhG7a9Eer2OkB4+ydM2P14WULTKfwBFK7l
R+AoLKpQ+Ol2rYQzXz3ynkxvHJBlYfRvjXL0vlMIb6oGexxJiLU7ZGVjixvqlhVcjNRae7fRm67d
i8LfcC9KvZH17NxdNF3tM2xN1Eoptk7muGshtg9/N2s1GE582/H+Njp5tnbyHkfT/phCHiBg3y3J
vBh80Rz+It2x28gaR7Inks59IJ5lSkQTuZJUPySqgtQY96EcDxU1DO1lskrZKsJX7z69R+L3IlGL
JjXrjzdOZhJeUIxneebklgkZ8LpS5LH2aiXbeBLQ6IK0SO0t8SzStowl7MwCy0YH2B+KZH7l3sTT
iApBO0OniGBREr7OnIoHPWtbvS5hzcINTyXatOrqlkp3jtimcrHRt+AUcYVFe03evMKI6akjbOib
dK9Wf510Q/WESokcYT6sdlYmGcBP0+3feRSEULphlNVX+tT8k7JFFnHm6u6CjJ58QYvSCMHtK37k
efbHvxKdZ4ytlA/Bq+s9rJ1Cl0Tvu5F2hFcLvaeR4mIFpT5kcEeuafhXULiriROiYVBImIQnkUYG
GWQ8HFufQB78W2+tfPAAnEpIqWZGO6u3SNXbhNs+QCv7QfFvbW+nyMxI3SSimmsaD8+B+jJXflIP
I4BZ7vdc6dz/NthpA9BRt78jTLYr+62x+d4Ke5BiDxrB2BNKpxnOtVCw1zxauWwJpPkjGZO3Qypu
d2WWWzvF09BWMzfqQSrQbiY6bNrUZO2Q6vEcIf2fkEWDoRr5vvBHqZmcxkBRETcS2N56Pe7vli9Y
kYpj+aUkkiiqnXVGmzANmYKxBThiO35VTa7w+4R3spglKaapbyOwMGo8koMEkIT4Qfmyqog/GDXw
Je+21l5aJi/X6nkbA2jlormuCfavl5bOXXTCTvHVe+z+A6vwmiL1cvUInjsTjz1MdEGdCN/gFFre
KjehNn5sIlwnhkDzZ41QCQOByaiXWR8JtJUnKa6gy9t3jSwFqccL3cfpPrvt/nPs03EsiedFtbtd
OIQpvKBopRy08wvxL9fHVCuz+J6fvopJAHRbDWLJaFOMFnRS6Z20S68Q5nUiJJUX5W2pWg4ZNtL3
eXB1ZekKMfdxh87J7m3xlmqDjjkeUHXc0ZN/voNdx8gPq6cH4/ftCY9HgEZB4qodlIi1xF2Hsjd3
qwuVsRPJ7/AczNdgzrbd5WJSD6aDQPUQ7RRqZX097SOVzQry/QBMSA4DFu5Ve2egTae1YtMDwuZr
tGnVj8Pa9MkiG69YQND5NFVNb5GHgdPTbqy4nQXSvAaiX72zhRIzTqTqOJvIq/7FMfyGXol+GGm/
1a1lpQbNUueJqvNoqLQts/giE+C639Wku5qofLxG3tDFv7QPMXXgJDqu7UcD3gNWb8O4PU7Kh7oN
D+vViUJ9Gdxq/cgPgKML6LZBS2GKv4ghM+UgOlwkpsrNdlmEdvQu5ndLs/MMndiAQa9azLusLzOB
S2y8KQTgenV/Fuk4BOgaaOME/sq0vLrzN6bQS/hjEJPLwazGdyjORzpCG30StnFBlzTY8bZ7031M
jonDTzU6MJ18AYfK6jTm3abK04NcrtWbNjjBl3rVHzqFGm3C4iOP7qW2d9Ej9Ry+GzmjMR1DXeK6
BIcRvHK+d7CBfXrJhSgjByXGVxwq8jPoegg3x4M+ueHWlgk5gLFnTp2OQ1ZVYHi2A1mITnC7E3Ck
u1bn1+5sleTn5dzlA5OfvkiRgQpmf6ZCaZKkJZwKnhH61jHxr3n6McxPCwBSy1UWd8DIPKffni8t
8m1owSrN+7NZQ32WdyTctJ0XU+/aKiOlGPD2UjE6gw3+c9dyHXyepgDtFiZfgDURYUlq+GyovBFU
oPISB0Yw9KglWOssbF9HPHiKUBoEUJqA1/THJ5atI15euB54ooQfA/U2y/G/fryD1Reb61ZTM6Sc
W/d7/Tx9GCEZgQLHIbS34NqHvlBGFyD7L/8iERbkqfIW2aR3/BZWVst8VC6HDMhF4ccVlx/+RSrU
GcDmjlTgHqF7JdDa7EFzFHEd4mYidmOSFIkZe/aK47AQ0PBzEBeR68Z9qcbO44oLBiSn/voJBTSX
ZCpU+SvVqchJoxIm2L64fovYlpDxyRyCuNN4gUxLoWeAb9mP8RBVGe1qRB57bbwSf7gEy0qOXWHK
B5kfxiCyLO59GLjMI0I351T9WYaDTBXNJQ9DI/I/l/BT9zkRCOxYrRssfmDu8KiAW9ke8rUGILdB
fJ2Yyp5BYIoNuvd0t34BvetQpDIa8D50+ADB+LN02u4gvLH8XVl9vO9Y6frWkAezpriLnwubxcrj
7byi+GtxHWB106Mx5fbQy0VLSp1ExzaEErrUajxuuLzqWiQyHCG4VmD/iebM2Axlmw6mNOdJy8YV
w0Y20mVC4Ms53JUIV5EQpNMKZGI3UA6NLZFYjiVfBQiXtsRoGS9AoSI1EQJY79+6D/E6v1V9TOTx
8/CziR7Qrng/Ozj+Ce6SIeEcr5469GdpsCoSm1RxaT7zpOgqHzif/nsb7Hh5sEKDLI9CUw8jsjKH
/tM92s8E1wyvpAFBIGiGgH212EQjQbKiqjBZVZoXgNs4OvFVhSyAsOWLwyoZNeIAP+VR+hXxKWYd
7jSsTwPBwaTnhz2JUfCcdjCmfIeLEtCZ/H8pxg9y7UsbrVNHEEQjqzUxHDbdOmOWK6KjjvoZlKq0
RlqSNS/picxpHBgNxGtEOQQI1OpRvmsoM4RslRrXOm12W3nSEDIopKd8FRo3w09nDnJF6Axphmq9
cZFh8+v7GnQedSyxRPwDnb9OWjTTu9KNuFGI7Tza29EHbnuJNJktAeG5F8uyr5CrfihZH498w2ce
O/EmlH2roEoBcQ+YGGtKlpFcOthDaKb03vaNYOX3oOU9It4crzGNZQEguDABB+wiXuZxvP8H69K9
jCxsoMUrWx50EuQNH8afoWj9H1saAb8AcKKROCvQy4dFUdwj0kZL/7f7og12sbVK901yOxBK5/lj
5F1WsNdK8hKUQAStSECpasdwCVwXJj0g2fQpEmst5rwc5FwjDvSRGmjAvb9SILy3BOonV9a7jEtT
UYhxmuVcICkCEN1GIeraFDugeG8wI4Nb0WylVrsy4GYVUSzSM1lBwtbNN1rVE29sUbvxwSpS+GtJ
embKng28K38NYNRq8YViCAE3EyIE32eBjl3XDnZddTtwZWzEOlmrDVyvyArJdC3WYKvXRinINx3C
A2dHJUU4vbo7JY5mTl+Of5ScFS48JMScyZ6yj2zvX2yqD7MAOctGJCZV+zh3blqhZTXHdkkfzYk5
4RaSD7MQLUzCdQVKaQDTAzKrX5qHF/dj7+i2+fgVOD279rMHIuA93agds6yy//rCfKkQZmiKOyoK
M7R6RFsOn4Sej0MRaapxeX/M+Lko4lqBkdawwjQiBI9+YYHkzl+lTbAnJz65YmHgE5AVR4GR32ui
HdnTih9AUruuKSISlVVIGxE9RfWiGzIlA7V3il7413xO/FTv5mcR0rlbTQtPY4KTZbIWOS+TLi0l
X8v6MoA6V9Um0AcqNrs+/wApV/l36jo2TEE11vKjdYofpcG1uXsaJhjzbv9HOWuetlCuW8SPRu/7
c5w0HAH0lRsFIlzqO6EHzGClfP1fKjdqA+kfAweQ7BCXszZ/2kyunnB9PO+KDdbq3yJaFyFAkl0i
CVhj0o4xpT9eZ3SGqjt1tz1hFasfKhiTmgDQAnC6apKQeeB5LMNEip2LXahQD3T6wJ4M/4k3N7qV
WyZ68dQQM0/5g2NPkGwE/d1ZB7aKinkFbfRSRUyCcPqcpGDhvP0afZR7D3MuQBqJCEDwHHwVJRMC
MLRhH2FRf7KE0wJNxyYPGX6SVJxXXP79khKRuJs9jtvCz/WW1Xf60UXYN1tgWkuTh2eaDlE46Vrq
lj2XARCBGC7rVvcQ5Q9obEh2Z86nnBlZnzfXaLx+guBKtY2+4I63qcx4RnyEPT54cnDuzN/uOvWX
Hges4ml1VUoqoLzzfDGoDuNkD6mDL49HNJ4pcH36bmg4co1Dw2ylOvstLoZJJl4N/QPbxaJaCCjQ
tFGSVcJTrMVqYapxZ+bMhN10Zyvup7SQMLn2CdvjhGZujl9J12BFNoQlvQNGcMvPG3YH3TPEp+2S
azuU+fFEpM5MLba1bI0FCvHt1hO+qhySLRcb1CvHhhMW59vqUL2ELuQ+npvlvIvaAJq2QFdQuSP6
IHVaEEfkDJUu0gql7D+JaOL2ktXLIqb2Xy0RB7iPp12q/hdxrrojiytrm7QsyJl1CvNjsNLVGmiT
sovWbydRe9ZLuU0CBKJnq7NEk9XtXM9ElBw4+OssUPkVMc8YOu8/neJooqRxkUiJASTG3d7Ci5TZ
KR33aMZO0ff3YSGAmn8z2WF9c4MWxdxiCUdXipWxQgCLvEiK1Sd8e7UW6AUBpdJs0X+WFKrk6s+G
NLdsSh3OvXwl53Qjcm5y5pOaZefERL2VOR9RJgnOPG1f+tfYj25K9NQ632RJOf7oU53Ztiq7Qo95
rFqW09dwAx32/X5UHoOKjZxJVUNL75uAC9bHMIQlC1sJw/YA7cbALkZmnB3u0kP1n5v8YWPNn1dz
UJqCQc8JdEMS+I9LhLGY3wyWPQYiOfZPxVSorg4J1u4ydh0rLed2hfhofr74a4ojtjb9mEhJTiKy
nECKgu+8Chp44L0aLVxbsih+wgx2I6zrkssi697562z+iPmR1WcvIYqdG5yeQDloBujhtPYAL/d1
t5qqzid/5z3WjyjJxTJnE3ND+vgYmrfF+vZjVneJYPnGwKUydtiCpbKu8qayZWlO839UmGClG2Wm
Gnl/8fBnKCaOQn20afSV/V3+mqCfxq2lhXr1mi611FYYBSUu3J6YrUyQquDJLrbhZrFnx/18WqL+
NuGWP8yv4qqbeNubSyQTnPmIMGO2kFFIaYV+fnL7lDD9HoPsqiNlg80RZijQuCQcsn76JyGPO9XZ
rPj4D6JgRM0GXVYBYFi20G0/Plz2cHpKon+HLFXFpi1BTdwJna5tnRY0VUAvlMLSsWXwhB8Wvbo6
GaK6wV/rZUsNZns5G4GbjJQ2vNeOculFdB2iVE174iUvcGNiAOcGr0gZbgJhj1UdIAsb5bLIZE/B
lSiKoInJBvUxIA1+lhbDApW5XhuCW2GZIbSn0cCrpCUhdnyi416kwYL1p6FIaptr4ZKbQz+Eea1f
1L4GIbTnnO/hNMlPuVhBurXBmKl6DPCCMTKB/ptXMu//yvo3V9t+7KiNaAi0SnqWEVPFt4/6aycS
AlrCpIxFbaOeQGxEXFc+ZeCWZUx+EAr6v2hlD+MuNnd8/aU20yLqau0PJCyJl0enyZgw3euXrjyw
KTlxet7Mh3fUmRWGIC7u9nRnZekF0QEz+FeNzlHJAlBlWLecdImTL7q2IV4DC7gICslQa/gn217r
eoEeeBr9o0Rg9iHp86GEBiVvEQVRuAmfV3m+Y96HsRJ8J6hpTlLO5f4gik6dKJ3kj0c4Zc8BMjJp
ck4yB1kvWkQMQla1Ex2f901C6XbrTQnUZY2q62p0e+PZZnMcK1KjIGnaJYD3ub1GjVIpZU73BpWI
bDGStXR1v3NorUt2T/JXqrP6ku97utY3rwrxsKAcTmJDYX+RkI+tfZtisF2p66XxezCzscCJeh4a
ffR9a4VwmzKP+i6DL6Bt+45JOlO7K+XXmuPpo5/Xn34CQ/l12on6dOVvF/DceWelwHStRZ01qDpD
E4eSVL5WUxiLKMyYEnvD6V1ZgrVxl00OFy0+xvbLebbdZjCkBiLZXywX0zswRRHwZaiGL++bQOkp
XO7KkhI2kvKzw3IpY6FKDw25qGf3RUwvkNtFceOnaxF1uH1/WelYE4RiiS/HjWnm8KbRXDPvgq5i
y/U5sOyyxTP2w+zLY2ecb8SwDT+AD4nKGUUDpHDdwZv8Fh+/j5Zl1uSSzph84Mb4wrFBeFPhCGr5
+drG9y68aHx5hlTg1ozz/Q0uKGAbj9WnrF5V9fYS9X1cIvIod1CUnrxVaL8WBp2F3eMiJU9xiWvS
JvXLnAUXaPIcqYW6RNQpQ0S0+4OhnHtkpE5h9VsWxFermO9LIYZGrrzn7qd+vQJI+i9dXZiT2k+/
bvqzV7mUuROUJDoMdP4xvQ2e94zUGPNu6KFwzjPlE1tbV86FRJemDkvK3RZPXinihr3vSVEKqEjn
//hI775DnufRWWglwWeoJdHtNsRnL6e2Nmdxa3WkeRl9Rn1qdufPsVdZV5BkQY/gmt49TnB1ZQ6o
Z1RtEi5vB+a2WtJtulgkIhhy7NBT+KeCMe/DgfZzTHhYa313EUAR3CgSiIREi6eoSDBvKQfj8UT0
kratQonUxlhFs7Womi6njg/BiGkSGq7x/ygXN6tChrophu8Syk6h2+VWvpwLOuninR0ESLvEKTyM
/d1MsdqlhvM+5HcPPN4cLO4o1OB5ZUqbO4+TZ+zGOnklRUJF1ImJKY1oJ+Rwfdd5Y3JkzbJ9aYnj
eYvypU8vFZEwbTWqiIB3U2wsMBAYEZLsPzyR9cd0asZMrba50xB9CFn0mfPoZjXwN60zacgda6H7
FkuFRlKLzqAHZ8cSM18bqdVxe4D7X3J/6NUogyz5PZvIOZ2Q8EbR+ItCHWaBy+phw2XMhBReriC/
TRw4o2DHTJTy5g6+kBCaHFF/nAam0ae25/G7iP72LglkY6U66Hd9JyW9fgpw29NE+ju4Z5feCn1A
ItEqDJYRVlaDuK0sXFVTAdm3pu8cF3Xjf9FhBxYtv38m38SxgUBmKo8+bd5PT1j8uULTEoHs5BGU
fbD1L7q/P6BlY+f3qVwDWMUrBZ0MJitYItiC9xTPoN/qhJAA9Tr6nQPOpxSmymjTKUyJKkgfArS6
HvJl6dXXkn7ZbYS54KNclbumoBo3Hwi1Syfstlu36/DsjbZP1DSsWzrve9OQQ0vkzCsN54EGe0ew
EoLhf3zUNp5ijWxLCYDUHlpPB3S06iBN+kG7HdJEUpRXuHLlVGuEKBzVqE4GLKLfNE0WNOsJ6C6f
gnxNewMKV0x0i3KXTZvm29SSPBqMe/WwG93ZQWuDeqAsOAwXtubfOTeKyjy4Pj2zDhqr3CWAUqed
epJf/tc+nLtpnjJSoV9p4PpbhdWZ2WyFq1OBlt4E9+FufS+n5d6LQei+3yTu/SuT7th42ZbKWCHS
Ajg78hAU4B/DRSR9RfeGLT2fsqKMkHZknWclMBtpU9GP8CIQdiffhgucY6DFrnqqyN005GKLvnQZ
AqgQ97Pfi/rhl6nfgyMdLn8d97OgWUqpgK1ymmJ3RMP/lenpZ1nt1zmMvRZ1H3OKM6CXY2dWnHbl
MwvoWJVtrfat9WjlnGSneNjAaRVigAIsgG9Gb+EtvR0wL8F+IzUjNESiPKwfZFDaeCI1gC0bwC75
dQYvfETYrNfjAdiYFLG608RSScEEVAWcQ/Cb2aiby8Aya+NGLC6a3WoY/WDngnvnMcV5M6R1dbyi
CO/fCbC1tLYAKez9NxfUtmKlPWxR5MjPicmMvzZGJ60Jy9G4DXEE2uIj3iP8VWsFZ/uaEV6AxT6A
AL4oqSBQ5IxNhwTIPll5B/bOYdu0Vl1dr1oZ+gUd40b5y8L1IhagGPtb2AiZY6DTSDCk30p9qFDB
eKKXPEnXLbkoCeiu8k5UHbKPgf6NNQ91bqa8mCKOoeS1gA1gQAic3Ptp7q71wgkh7ojFLeepbfZt
nq8AY0tqtfjrOpNf6KEQzTJuJVckWiXEsg1cDrEBTy9Ep+UY4iLt4jYyqh4qONu/6QeQmDRYKqv/
ZX1/Npc92wO3ncNhWhaszqqbQwSfN2Wd5b6/SDPZPRbEJzRBEkr4SL2DQ8NmYhs92L6uG2P/VPbo
lTzhIihKq1Kk206eBZ1QDUItRgBZN98HKoc2elouaOvEkR44UPtidmiEMAO02e6zqVie336RjJbN
HEHpQIF3dUMy4Jn5XRSjNPU/1gNp6XT/fxCOD/m6Iei5LTEWmsOUikrrHo9I5q/RBIJbq63zEVuQ
ohVF7KqVX1/8h6JOSYWbtiJKEmb01/0SgIwISxMY0YII84a3PE54Gyt7RoWBqHNZb8Ky3bVkxMAv
c4x3HBfXgxuN9eFik1R/+UZJvbgcQ/DrJ2Mlw0iyr+zCyA/OHiXrXV9xgPq94sLjyA2V6tFwr6lc
D5SBc6Vo3FJlkPQijXUQPwIJNqFhpaAR/MlMRbhVmRsosQby1jsEiunvkeq5ZjlwCWyUA/epDzws
Ryxw0aVEvOjWx8MnDrnUEGF4ota4qmFA9/BxX35FcBs80GgfMIgKgmko1oiCOOCk/VdKpsVVAvrh
pvKgt+gApcmgZhwXRozLRxWbXNzzE89lEGjtwRpxvqoqDz7NuvBasY4+eSyMHlJiz2rAKED2rSOF
AyRvVI35BswoYndgFmQjx/BoDoS8y8RqesusYmeMASwpbZJiKaaq//pWqWNref2duTo8DX0BHNq3
JiB4uQYk9gDvPCqhkw2RFPj0xeKg0UlgmeC9eNS2v3lB8JIDmUOxhQPy9UV7WDHuHHaSrCg3EUch
/WUcStcw2/HRH+4KoVZZcCD6q9iA4vCUIcSpCXQI4y/w6wYuThs5e5Ea1goM/Plikx9AFKT3/9xT
9Br4nikXNPDXLghF0gDAvUFFxPeGqNM66h9wo8RJLfdc88pXTSu06NGOOGqs7wKuML9M9yYW0Pmw
ZLoaAltmFxZEUgc1IhbjGgXezn7A3yZ9O84fQmQPC5wbb5iP4u7o2Wx2RN1zpdmLOzfLMz+5u7fi
C0E+dsnV7vT5NpqgF6AuS52q/N19cRYRfBRDMmUM1spfpxAHRa1gLsXaYSbRm5bn7oMFQowNwG3T
JNtAeQ6m8PFeu6cb6/bDQTAhsx9Qou0spXIt9ibHIBTA6WHkwCukodqlktfZqR17MjDStPGLtA0/
90YrIagMVGw5qQAxg5ksJ3xVUDlPS4oF2aom8/3ot+smNcMQNvJS3iFvCSDQVAXgOdzMihWffZDm
g8K0smbd057M057QdosP0w9QgqZDrHyqA37O0yTCV1Xl7oomno1swxC7INjMQsWq4NC+gw2VenWP
XENcFCK6yep8lNkJuEz2liE2TYqhnfawgN+dJMJExUAmQPFUj0qBZ4KvS/iRIREAA6OMmxHYsIeC
gWN6pnF6Fb0Q4iiRqdVucoFVeoouswGoZiHAYQrxz+DhbwzmuTOHOm0YeLCLiqiLD1XiROU8Ze7l
HA1BcuIkjzzFypxW7rPXcQtcfwnt8BRcQfIWlXzbWJ0+XgTNpKYUavEzITG4krBGS3YJ/QsNkPG0
yiQ8o4ZztSGMEPp9TjUjmkPBZ06z0fAaVSEqiYAtievabLY6iqRYVBVMhmZpMJGCtNZn/3NxWHHE
lsoKKlGfNLQdc7bAsemsi2VDTpqXK13ttC0D+OFoiQnHc8AAQ/7Z4zlXvZXPJZjmP1ayVSH9wMkz
pa5Zavzc3pxqnsIZs0IHUx8RtXbGM/7PDu2WNedcYyuqzaEVv25EZ0ysdcKJtla9Q5Sw4INtSQiz
y6K3oNd4UfxPHt59fCRKe5XFeBP1Vb4Xi6BlpyNYyRI6+LUuBgTIa3D6U3/W9HiOLdBw61DQ15f6
lIWEV/kUVsaUXEoQ3Bf68oUTAgfyQVQqvTx4V1llyxxB+0hBQ9iaFZZ5dy3E8Ch2Dku4y6Qe8q3d
hEoG7f0xyD/c2gbjY4wSUIsWE8LWgtrOaSwO5647EZDJqS7gOT6doyA3VtFHeJAxL+yloCrtsRzE
U90HcvLcp/WVLYQvjVe2qTfd1mKrBTlFLNn87WzkDuqRIqyoJW5zId4+8mnvdRJv4U4hWKQIfLHi
rlMDiiJMw89CAdFcOPhk5FWA/t3Y7+8bB2wjy5InOId9CK0KMCDaaj5pAI/PTnFLBUipwYzPF7nZ
4PX2pTgqoqtJPxXei+LdDInKO9isnBtw2N3+gqjFidqGMoOyoeamMpODE5IyluzyTY04/MDjVRQR
LaJCxF3lmb2XBztLdYtA/BPTpuY8JoMVF5sfsMqHLS4UWTf7ptUGi6JIkUzpoWoUCD5pfnmsfPgM
KHqZpBq8vkSnMnz2MTHEFFYjHxaqBeqfzKqxVFWOH6PHM2Q6Vj3xYqGzjBo2EkZG/Ee2RI9bJTTT
hwGhGTJKgA2Wykod12ViYZiRil4Zy/+JSsgn4QuYiqQffGDDR2vVmIT+tMY+MHmR7donzEWgrXW/
wPNiHLSruAEgayLfCMNUHZMNfu1xuqcFQtjgasfYQyiDFQYtNSQ3cooUpIPOIqcSliaofO8V+FoX
lTP7/H2Lbm5wKYFbJtJy89+IFJUlUTHjpEpqpnuvf4qHQ2UqjiYj3wbIq0pPrBhoDaw1ZcON9cnz
+zjrdNqj3PMrlBsBXMD6lVeSGhrdjx52W7+fa0cAiM5dckTDGpxICHU/pjQPtJtpdgOJZjn49Cvh
NasOPd8Vc1OnNuxunCFiuEqWTsuD9tOswnka1RSNU69fG/t630sFbGp6YR1vNl5Cc0Kis0J0DtTx
1KMdP3r8wAbKlPhogYzRBIDdhVpOwJPzwrDd/7iMQEvSG8ztwQMZWE/L/k5XE+EQsLawXdmXr6qI
CzG3ZWs/pUsUgfVUbR516/FrrztcvBzzu6KarjPlRAjKsZUh50DLKZHsBTp2NtUyQ9mURk8Etjgj
b2h7etcWHdlwwyKl4mQ4JfqFahKq6yj7i2o2/dKNqFsNOUaQNiPi3mDPXHC/R2hlJGsTV5O2OIqc
UL7IxsN67aqULXOcAW79q4kdgYjrI8ckLYrwmfnMZkadDYxrxVyZCYLHjsFIgQxlIN8Ete4kapYr
Q0y5IdAvHK4DV72eMOw8rKRIeeaZylJU/pJtnl7wSJaQ74Jh1+uTetWOqSIJwObdMy7P1dYkD1eX
KKwRivSgB4MtMgovpBJhO8hxDlNsafI5ZUuWqNrRsuMwV9AIJH43s8Yvsksuyh8JghsfeJY423Ij
E7wsc2PWI8GN4A32020BfzXOaRDWw73lslkZF6QK4UxFrD/2Tf1X2xiMv/7jtag4VSfvdkbYhYZZ
IXU2fd6MTtcQJfj+/B8P5FoPM4KAIm0aXeAvib3F/K/AcCoE5y6nCwZaYhugZNGi4+Ft+91de7Zq
6Lnk825fJ8NqjD4nTRDPkObGhdaCq8NbTVvmI912VQmEa1qZtDBbQ0IkFzFWsU1EcODnQxz3bwWE
jsdaGPUAdV6iH9rEXK1bwgpVR1NzACoxk0qdcgEIZKH/cn+4A7ptvPLodR3zHO6Dw9XVnvnVsyF4
cyIOf+wdt24g1xkTDgOjykImuy6aYIs23cyFlJHIpo4r7ES7Wm5SLzoLHhkeV1aib93392Eduhf1
3XmvA2rL/YchiP5xOWEusdZuPr0MQLVMINfAeLGKC2qC8K2CSUgKO2ZfORc1kxsj5uvk64Uu8kvZ
9DBoGKyVS6MG6KxHKqgsPFNwG1vnaBx3K1y7swd9VT4zz7t3k1UUnYZHuWxyVHTuzFdmTSfxJLPx
0f1Z2Dn9qHzxjP9rqsq4NxXnDWvxCiZvqAZtUmVbheEHbmmFAHL1azVwFtpyaSw6V+40GDjA4zoI
1uFv00ueIDvlJgrMpQ78BfKiud+SN0fTxkNEFUxh9ywBTAcupBvRii7aRjtV5rFZ5wC8cJaQsDFD
Zu6R1S54KePkkL1V2uwZPrkfVrwg8tkxkAYCggEUTshIK3a7s103R4XrH66xVbSWDTmO8MIHV2uc
E0A9d3IKLfFPAQ1P2eRsGC7g/Gxb5lTlX9g5t/YaW6up6NdvZ12cDxW+pT4AngpRNT6YTPnBiNtX
evUDNRsJC9YbAVVYX8lv8LIpWkiY0N9CEnBaMFVLFF7d8dPMl3su6qfmdfAUces3cKm/UdN/P3fJ
HBuKXTgp9YNlqMZfVjcqWXg2T8qb/GxuYMl6s8ldhZ7zIW9DAK6rHasXSfJ3bShJ0HHLHZN6r9Wk
7z0vmMBkFDKIhO72p07tNVw6TnTTav6pKO3hFAUV7pCSNNW+TeMXgtSWT/UGby+bQjKL0LMV90Jw
YhO4xHTsLGJf57JufZzNvMjtgBkVcl6fPnwLR2Ypn7LlEGk0cFVE1/FC1d30pkPoLo9Uc79ixPGw
m/3nPVObo1NofzbrJAlG49BRNx4E7o0pqSTz+PjeSDAh0Dyjcpr2yErDsJOjP6tmoSDLOMwdI6w3
gFQBarzo+Mdep9Angx9iYGhyDt+VgrSXHIdg7rJm3nSHdvadrkaQxyK7gI21PeI4WSB27Os+E9ip
pwkv78Qxe168u7jYWb6UEHFxRlvnSbJ1huXLsgRGfrJAB/QtA9Tl4E1UXm07byFF3KEkkn9FInFL
GV1hHgGb7knZQbg17xhVGuuiB+0nPSYKCAzbhLJUSN5ZJoX90t+gCBesAjdhakZgDdK2uVXtM5na
epYaGs6JAaI08CrwIh9KCEFW4XlaPTS1nsn8PGizPiuIZ8wQOn1VvJwotkaFIFY9aY8K2KtEwAmC
La/HetgoAlggvp1/q03yMxoPNJx8+28n16mJvL9Pk2jPR86MRgka7fhz04MlOsD9J8/ufkbGJByX
r/xmvKoj53/TCnGl23BD7kIPvPOD7cfWQVj4sFV8wAsL0R/87FGJxPMGlR5CdHQVWpEqI7o2mWAw
bHWAyg53zLTB2KTRnqvRpDHDnK2i6qQIjU3lti14e4jcu57miWW/fE48akQY3+wIPfB+0COMKXVv
IuMDstxrF4yJnzjpSRVyxjP0h4JHm7J5hvF4Z9Uu2W9/Fe+cWnjwLCo/mznEcCWqi8LeeAodFJXB
nFN4WrQWRQ1g6LaFx5zXGppHkifc6Wk08vUP2rBMre1M1bRi+RbADTUd2AkecqkLR8QrhbaIFmYu
8Mx19VmHgtMsYqe0+J0oGYAYRexS7kKsjP6sVxp9aU1djiAttjtZvytxfs9FMsjOgHwb0k+B/dSD
QNu8dvlcNJ5LJD1fhI/6YZ3CU+ejadG25Zj+9PUvL7pNAekeDAD2KbqHrtUn1Z3NpJikA9II+Hvc
CzJ2pW7WKbtAHIbkkfhsgs1DeT36QiRJs2xsXv6usj+cyLonrQmN65KIfviijHR+LByDvOdmJ+Fm
XqQj+Nt8AopxEuSogwU6SRGuAAdZ0GMwypUz6IS6ytnrpvhEGoWdDH9GNXoG1//AojMWPB1Zn9y0
fPn2uMhByhnsXnM8cChtXeQqjbnsyAIRHK1lYttQn4CFqYGXV9vCgnal34ZDhEs1UqftT6bgH6JB
3kEHm5wgXTIOnoNW+tcEeLcZm2rJ3z8RUvSEM3VHueySXNNaHnscLdLH/xQvf/HRLSxh9+snyjyf
r0DepTGWOgs09gSUFyfZys7xizgaWPBCvGWbpfmjyHMn+SJmcV267jGzBP/xkgdt2Xjm9DDBrWPu
iRq28WCQS1tpJKXl4oo8bQjhzzRpyDVAPe3vJcQXuv007eP44qghnQ0ozwU1tz3FkH4nPpntLDHu
GZNMVBSdgc7t0qPJQDaPuDrAUw9bnHidNQLZpjzfoI3zCkPz1c4CQtsWK3b0q3ZxKiv4bvJVfDJu
WBQTGvJBqOqpJHLU624HHxtt5nIwzzNgo9thsbOqfE9onICgXyH+V17Jrh5GZJgjGgYK6VlpKswz
sWpFDt9yWOpC4FgKOSNRT5XNkqpBO3bJ2vP1cPI11vIcaASf4ATLXzzrR089yp77oSHsAASbqi1X
3/YApjdktSGv63pjGLbUWnA7BlOoZeGcCbYL4+6PMaYhAc8kX0Ns6WbtWAvynrd1RkDIYnABYrqB
FScCW2FS9b+KrRH/b++Vvkocf49i1MCuH+of0rFsWVWvtYaEatO5ZJ+ie3mnAsaifRTemFVaCLGm
aWwoBmbF7QC0Dd8wSezQ3hJA83oYT3LKbO+K1cwcMjbalCLEIVvNsn0Q81JmanEUIXUqE9yIC3/p
rAVlzsl4/H5ua9lvEAgD8PDiPifUsOan0iVJqRVQe2dv8/suDP4LtVnS0huiWCaSW1zXoJpbtmh+
YmLwPeCVE4qqNmEM4b77K7ltU+3wwlscf5qnekLVXKZrLJxN9EjTBDAjg46JaVF2ftvAs91IzpYY
Bcb01wpeeTyd88CkwMOl2NBDhYMeGF+VcH6w8cJU9GcBUCXWBKrprySGKgXtCC/9dUG9xr4UIBoB
S9adQoCZt7UuYiNfMNUBb3pUB28Rk0GuxGv887lJRFFE9g8mHBjHfHbWPbxMoMDK+V3tRaqqYUvw
j5B3/6B9e/Xo7SrQnQ1cPHq/2QDy6zNoA4u7JLjJLOBQLRI8RNpxbCZs0srkmoUlkG0SB8PAkBXW
3HCxzpiQgfbLxYdVbA69xzbuLm6u/H8zALztoM4RDeapgJ5QqptEzOqEru3HjsCRCLY3GygbkrXk
cNUjjK6yhZwoXtdwG+aLVZ+c8PkcCNJTENBrBY3PKyAYg65XkF6DLnHGFtBRidQ9UJmsW1c96JcQ
nWv0m0gi5s8fc5ylLkoctGPK/Ht+sglJpAAUu0YZZo0tWdEUyLrnZED8x30Xv592K1mWri3fbCoY
EpbiMp+HSg5Cd1zVMfb7kVy4Pdne8FZ3yM5HUIqnwQ1HNEb1Y+/2I7OC81yTTDuYBGPmJrkvK7aq
bVEoYMLjglyXIufWtt2tv+boHy6ABPfldxAdXOoqGG0WO8tiKp7MipSzwcVozZ2SU8meaNk93YTq
NgMaP4STm9Duf5hbdluUAnLnAcFEgT9wKRtPhSdMF5v0Ek9IEkOWgmkuH3kbjOTnkbhMNkGYX4Yf
hT6kbtdiSgJuNTFPU6dAXFnn1hfgTtP35lCNFZ7Vr+n50J9nvTbkK4SI7siZDWTgpmbGEhNOKo1r
tppWSPxPIMknuS+/fU3ta5TMMZ6FJqcpZa2MYK18E/IethcXK87oEB5/Z+MpeXcTzajiwVcvO7Nt
FjmIjHCJDlxSmAJ9ivL9xbArHjwfsbDBaI+1/eFJ9Wc5VHREyN+iNg35IHEqcbJK7ZqB8Doow95P
Q1kStRZm0ODDXZqC8qtVJf6kIbCJw+oQbjRxm3NbOnCer9l6+mf7vS+AM3YRLbLW6yMhRLmj5ylq
gWKRvWCyIeBY9TR+QtDCPvnyOOZKKEZVlNovUllWgR42E8TBrLgJGg6OqngWCnZZe/CWXfwvK/ys
qJixF2El/vJadkWKvLUQusdi8iVcy9bl6+0r7IgfBU4hlkkzsS58r/tSnJXQHH8eulFeRwCG/Apw
fsoJVyUNfIeF8Ssx0P4HnH6devvd9D11AnV4TCWO0ocB8BVMDXkupjSdnxzn//PSOLC6RLuVngke
9VbPlykh9lCOHuccG2USNw/cw7owIDCC2dYFj+gg8Bmyr6IOjstI9Co7nsrHSbr6FNbPklcqQdIP
7PND3riFQQqXpEcs8QYitNfuLV4pFQe34myWCWE8bnfoYDfxAzOpUIVPNbHkZcBLAcRS22V0ewpM
gLY2Rd+GYPWVYvkZU4CcSy9wi6bObTwfYwf5IDbdGYthZ+4OwvsqmYohmPkjz96WOQhUpNtqG5uR
oD2GIOOlQciOdZlYumBkHsDytQkUWo8koDcWzPAQeUptWtQETUI/LOrq4CHiN4Lj7t9/+e45fkDs
gnBDwHCYqG5JNor9T+Rc/eciy/rcxZyJiaPcnC2XunhsSzV22z5MHT5IL3325gY6VGe3K4GD6B2q
k15XQmTkPdh790DQyqidlf0fW/lB8bLVOy4K8pRAh9FVbpR8sISJmNdnKxGU1RCVnUr6DIw44Rd+
+ZeuiE7EqaDBIvAtGd6jB+GgHZrMIJmUWUnaljAt1+qXa8/RDrLET6SxmKlMgmC1asjkBi5FEJzS
3gMKKYKhjloattzDfqtxABv9MOJ7zjWOsAN1ksOb4DWJ6iIIO+exQDBi2Fno0e2oE0PoQ2E/zYxG
oqagz8+tBhgrmcZnGLjXS8yJUzRP8DkBSmPY3lKyfYQFNfKpNL7ZaZEeiU68zzj98XtstIlZjT+W
HfEekyDdS3OH7gejRQC0U3DAiheuJEQRD8Ui5QeF+1D34cjuzEwS8ngerEEOAcvVg1AKxLg9Mvf5
oypKK3D7sgcHdPybNEzTMzWuL8tNNqoN2kfsogDBi6VGfj9az6nYMDWBG6BePPs+pe2i0uuRoZQy
Y6tQKJSJ2l3FwRchsP5kIuSfaQfV7gqHlZnYZDlJwCA2s8h7NszEfQrEjqVxCrQuD9vc/erhV+FI
DsEqQreanzMFdm7Ikg9A5OuOWyHfMPC7e6kWEDAXaJumV7KVSitXwU37FfRusPCrg3zU4Iwr8+qQ
0eodFSCzUUhEY6ZiD8mhzUoxwxw6WC2HAXY89YFSjxdvbIdz6Sk/d/DOksGvkw95Sz2eKgsXsqs2
hT4DOpo89Ma9C2WQ61hpGSfjsqNI60W8ozS5m09Jk7Gzz4dKPCdDoNxylK4Bj+lGzSbCdZoPmF/i
ZCleWFcOa0xdeKvSWWTTc/vgGOQqjfIR7poLYVDwOYJ3LazMDb4JyswYqmbVVTpMafMDFBla28/n
Oqrn399SGyFiWaYWysXBNjhncQlS4SqW5+osXw0y9xaxCJVwSZUhYsWX8dpvzzAtyahUJJSqBifQ
5/MfzKp7Vchzn1VXM5c1fZ8BRhU1RI6zGlJahhf2XEZ75M7crgr8pDO3nlDQgbwu7VMw5G7igcqb
1r0CtecpYFCEe4nCynNt9H0RkJc1701fSDXup5sHB3/mpUXkYHTm7BiBZ0RXp/odb1xr0NQIpyX8
SgrQKKGagrB+jnOdodQ4MNMEAYWwzakzDHSx2eNkcR+B6a1lbXCpzI/ocgW5p+7IhkTrqxyajPh/
K57LHIkZgfIP95jPsiF7cbeR/S1qLG2e9YrEXM8MlGQAPs9kg2iLY6hQYO/yD1xF2cL7GCGk24s2
udSKAoo5OaM6zSby3SWaSz4EEITj5VQBHKwcK6pU2aKoKS9pjWemQZupR+WSBFGvvEaAwEFfXEg+
Jfnau8n1TgN0undGqerovBHyMgAGdCXg6NILum5NBxM+pJMNHwaeASl6ICfdECvTlTcMzjB51XJ+
FzzAWsJAsubF68PjTl+RnNnYdwrBnJCpa81lw6fQjjoA8Ahxyul5iWRiZV/RQy9MOrEnKrG5AUnc
VqC9tbf9+P3PylvzfO9ADE74/GUvY/qp2OLqyaNhCQYVVlGdRa4CIbc6so4+UedXwaC8tGCWYP43
0f68bWtQk+0WhPq+8aJEbwpTiF8X/kwX5Z6TLNwLm6vifv3UPnhGYAZ9CDHzQYPC0D0npBXrIEqI
ZZcSMqNMhmrFXT+5Nw3JLHha0jcEd/fO6p82XxL83N0Mlpa7eeu1eN6dIinoNP64MV3ZP2UTiRp0
Veu8dRS7pRVbsIwS1iTOvVKmy4dfuAAlzt597fuWIGvr1J6MrRYve5zW2C0HAlQPJKY9rqJ3RC+d
RXQQK+VvDYjPsuIat81yuko/w7uan0Q+e0TXLikwjcPWdtr4QDBOrvlMd8Hy+BCOmyhuXzJ3k10z
TmWWwc6QWeOnAVsM2wgj7aAUB/hfH3Pxnqy5nZiVd04zAfEXVNl+qZWo8P1iGz97cueEhqJq+fJ4
bxVcYSYhZdbyYTHTqAyV6SL/MQKrIjvqwBQpGtdXqjk0KQECh+CchOUnXNi/ajbTKlVLohsXwYxP
Mn2YgtqXTjv1Eyug9JVVMpqj8uHID7HjLmq2TyxEtUNjIrPy7AsKVWglyIV+1W5qHIdL1lrJ+mIA
TrL/S3SnZpgEqfDtyXfmlmhFykpPqmOWRpooUccE53+wqOUmNunL8e49dof0M5cwbRDAUif3tEs1
PL8MLxh55tb0mlS8VnEO8RCFWyFssPDJ/voixPH+QAzsOAI1BDoErx4Vvt86PrFuCX5KYY5pPvBV
loV/650g/jqd+GupeTL38pJDPRz1wWEqPWFhWp62/zekC6nBJlm73gy/Ymi5WidcKfAOwrZ3YDrx
uoC9W8ZIYhcwUdhg2kW7NoWf1KinL6a8FIgm4iqNns29tghkZz4H4WMEZX4rCfjA0Dfkfz4JM/FT
94KhWe29J8/v2/U8/KQZ4FZ+Qq+c8wFvFXCaII/mS/sYLTjcky9z3x9xuEALYzkmSetqc5uWNg0a
YaJ0am0IeIAiTqeUKvqxiFYycVf2LE0WBs0RuUC3PKhktwh/m4MBHIdLFqzsrEXy2UBS/FRdkUPk
jx5/+2gIc5pGCSzk+gduYBLWKmhWAaHEjqBJLQi2sWQcT+44NdJWJrkKipTDq9kpZ7dsa2el1vMw
c8mV/ufyrDB0dSTZE+RGijazjI8LrLXg3DwbVcwCrLYrPBTLLc1XPqIl6uSrXNRobmgqfAV/8faD
lJPbsgUV+6GDBCmRDq3YrVvbB937OfGg45a+DERWj3mDPKH/7DIwL2l7Qd4oiLWXBJ5I7zxoC2qn
hudIBCYj+3Rd0qC3i1e9M2RWqYlYrYnSto7VEe6JzCj6/YnrNHeVKlFfVCKaQa+rnn3QUrn8oeJJ
tMLd4Rd/+aaP5HfDX9YOOXlYC/zwLEAOyYVNc+LmQIygLppxACqCliIJ1ul7KnFlhQMAO3p5zty0
TRQ0786Fvq5GIaf/l/rpM83Ym2VkpqzfNof3hfuV/CjjGUwy35c8hTcK3pcozdb8WOjQik9bySyN
nftFJuX6rQWj/HiV+JR1LSoUa2JzNz1jW1D1GB9JT5unBwyjHr75r1NEQZjyQWLhg0i5SMNGtw41
IL5W0id97qbpdCcCmuloDwktaKTcTArj7QQyC1WCd1AWZ0W1cLYu5tuPehQuh4C8d8sCrdKGFq51
PGUBFFxCcqY0LOy4UVJ6GGkAkFbu+QUozr90cNSfOO1CR2N10SYuk6ETai3XW8mZqE2mphY/ye4s
VCzL7uRUQLqFgm5fccWoDKJExCt1xDWaB+RBVhjdrlMpi444VmjyuIHTo9Od1/CmxARt+X/hD6LQ
fE106X8x84uHVXvZJY9GrenyxK7m2mbM0rzTz/xGxa4kpwLVHwH42OqAdOqtSQ0AK6AHv5od9w8P
Ybnz1vSwQy5N9BbwYHSmuBgbB+5ZhXmvOfZEXsqP/eDqTeYEYU/i5joJm+CbTTvWV7L91dYh79PQ
lQ+91QMDVYLPiFN3J3QIphNUq1J4Q3oUw9GMh9A0HapkZdnRTmk0qzHbtBbZNUcr+du/Ve1J+sap
eVF3mqVqU+GWTPNLy0tiYNN+TJnBHGTSIkUfNdeVNOMBEKCUFIeiWT2fLOCoZ1EuIg9f2fLYKLrL
EicztVpvo2blzujYixM7hqMTxvHAMTtti0DKkMXtOvYRH093OCxJO4fn6vsgPfqfrygGybj/zEhS
T+V0RCVGor4T3fN7TasMaTBx3JBNwk3/zu2taokbifaCLCZJ98hUZVqOiNyM18KoxqNZC8P2BeUp
11hwf3XZILhmvHPJrd59o25IGYIrEXcfpi12UXsK2M6WFfXz5IsljV/keZxkMCQm6kEqx+CumXHZ
l685L6A7YYe/gOg4iwKM8+3PyIPcwtY8xE98TqIPMhi59tnlb3CjpwBAyXieiGugLGO6TIh6EJX5
NraGbQ+poeIrN8VznoMHbE98tFG1kQH1HUUN9dRkJ65aEQfk58GBelJ+j+0PqpioqtgZYeywXJTW
uHqM/JHex09v/FYjudxdxBCMucEfI7ZLQnf9VWfHTZ9Ts8bDchmGDopc8u7A4J6eKj4VHxMCQbvT
qHQWwwawl7+RKP2HaR/t8U/6hqnftJr/vRr8SEyQ4Oq62kn/xSkbDAYhZhRStmnmF1ugs1PF75nv
+aRT0aEcatfzjgfdYMVFIuqUOaVDgxs2yqBFhygYP8AYPhGPp6rScIzUAjgapBXLLJaAo/n7AHYU
IQyu2ag1IBvz3o+AJ59a2ygXGSyFC8tl+erQN/nSb3008S8SI+YJHVqchm7th5OqjuI569qsqvrt
SGDCZv12nUlkegVgOP6UhVXxl5kXdDfOr64Hu667GD44IHWewU06DZ9Dp1l8kqvrUTRRdWriN9g0
PO1mXayn+43xpNk/DuT84X8150mRoprFEC0QI6U29JRloIK/PZJEbZJ14d3lZ11Dyh0wEnjbFRt7
LjE/ATi8hV4rjZDg6gvPVtyhspPnuNGomgRqZfG/J3bkPGS+10uQWvbZI/QF6qaEhmJug43PseJl
0pJBlZprbvD9BAlGVC8HWuPEDkeNjY6QkttiJKil9d9H+vVcxdc1zsoIIM+6YW8ijNz7IyRkk0dq
iPnTlXWwn1F0k8VLIBMO5FSxg33ywf8owSMlITH2GwsdC29yDDcF6Po6Rn3xfurC6arfe6ztMi/P
o7aV/K8Md3Zc+R1jP4A679uN0R9pbRJDlZYtXLrCwC2/fd59JHW9hp666aPdgyzPDaZR8KtJwC82
sqMXXj1lf7LcDfXSQkcbacQU/j8fyKxfu50tB6Azm65CopPamHF20m/2yVDvtCxTSb4Io5VZk6ta
dWX0lGfXfw8XAycr7FQ4vRwa5ivor1XEWzsTG6UGDvNZhV9b0UEQfvblmf8mfkNYq7PfPvmiNkVz
bHudPtFtVEhoxYmDLPh5A5/VwHSaThykvxbdxgzgylOKEFgwDSgxle9Kacfnc/Bf6vphTCG/jhc4
e7Yz3OKI8OieFyzGUU8uq3pjv0JO683FIya8/9U3MPznIkDWhphEh9vjtL+biG3V8Ko4aGFQQekc
9hFoa1NvYVPA5ifKp0/2M2sTT1GhURVwIHBLbsfNEcM2OgyCPeKfO0IEBM7uFGr3OFV3dKMhxaaj
XpsjDs4nbSR11iyh4zFOQhMnqkjiLf7ZK4a7eYptru74c1uFi9zyxSLkYNhdeMpyZHIvSdThstri
1JLtncV9vp3XYfjbWRA1PSOsih7iR0rv4QYkz098YQLe0WDtt5cTB0TdkQB3xmHd3B1Ccp4ul369
LblhhgpGE+DO5lYIoUyRgWuYX/jb9XlNppkWoV8gDi4jKlHbUoUePwskNzo6lkx3VyQiAktQH6ga
m8fRgXWSdaJFbLflQnl+/bu/MsmtChVD4weDY31UJUuoheX9iRFNRWPJMOiLhTEr1MN5yAKyEDBi
JISAJL5wp4WuKnDpCl9+o/Tj9wktlXep+Ow1ajNWIZmF+9wu6A7pZKRfo4N6umwJLeB1Bb+2ImwA
8/7h4VgFnSW4MQi0orNr9jhtCldUUbm5+UWUzu00BkUhqVBVrkuEIUGaDsMSs/LvF82uVioHh+fK
HcvH7j27UWTfsycJWXMS5ukdbdgmZVwsLIi77K53jA21TQx5zG2pq8+PZunHvbCs3tZjunx64+Op
8aWnkcGjnMyPS0BOfgEjWBQUUcIJ3LW3knOGs4UyeTDYHgcmiVojLxAbW2NXRN/N/zhp9FOQbhKW
wP9rSbrNoWt2Dw3nadzbZHdQ+/WDg/ei1H9z3V/O3N2XkQah3OXtWi7VC5cs61YU78IfhygsLyAi
45cDvB9q/jbXXUb+ILier353Tx+2tBAlgmMxH403c9+X0Sg1CLuaiioCcf2gYmEJmn+D+cb3hbDz
TM19GZSr/y+V2e6xnCycIGoAHM32tD1m2a6To2H87xoBnwnCEuSJJTRHnoJi22sMEgisSHSgmbdh
ahmXXPtvwiCAj18LXmENGP8ki56L3g13hlisg5qegH/h8WV//XuOYQElVF3mQ/KIoBsZ4Uf/CQqz
p3zyOsPzKjF/222kZUu6MsVf7PLozCsmj8j0LYKaMug3jR4gHmBenBKAKgImxgxJcBjc4uzybpww
/LLcSNsmB8ItRwEYA9AAF+cgYkZE5JpyALZO3GxJ+p2DQOQiOPJuAUnBVVArADLj6xUHqIoyOv+P
4zUqlPJFcoSfYgpOn4M0Z+6YbdBHtk9Diiv7oJTgaBfY0BkpXQlHbpgQ5xIbBvliUI1LYAIPZZJf
b3unknxeUIvJBN3k3tnAZQsg+gvgfrbN4wv0c5cH2Mu97CjdS3M04ThMqQu2jslaT+YkMAajbjdG
VQ5JdCG9va6v2SGCTb1WUxaLkzw3oguP2D8HEPvIOtzQD/bRGJcURv0ZdsVnwvDMAi3nEsltc85k
auSyUm3Pe3R4fpj8hHUu/PnJLmReNPrGnZWPeA42hcbxltfFNJAW62zghDbcCl26lZCmKmJWQ5DD
v0695HWJ90RSDZelrieyLhJhaLDvuo/ScTnKp2Q/fuOIhw1HIRdIQCay6KMiLQLrIOghnh3/urbG
0Kix+JSWyIzovAe24xkByvY0ieIXfYCGO9Fv6RiFKnVOQ4FRBGGeTkdcYIZLp8iOUBi/dpL44a3r
MqUe/jrRgCsCXhYNA+0WY5ivbjcljZPiKMSkDMJKnva0+agVn4eAPM0+74NKzB64B7gP45zuCINO
/pzUEkFGxT/k5wkDHj/AOCs9gcFYU9tVLYUHZd3n9sKYhJMUUNceTTYQm9m+uSFH4V2nvb79yxuI
X0N3+sj5maGExcXnN5zcHxuSNJnhoqKeP2JETo6xchdlwXmIenTUZHA9xfFLKt4Xqoeb0+HAIcbG
as7NdK90XdlRD7OpBQXLdsRavRXj+es2cziJeoZBdV08QLV+LPiUdIpJwljbR3bLba3JIsNuXWr7
foJKtv+jsNArMqva97Hj3iQRGssTzgaVxUYq3wjDhGYov2nPntbMRcNMbkFLT6uIZPeJpSgdKpIo
O0lsySVPOsRY80D0lji4r/cZT9XikbrZ77M2NHJ5EBd+VISIZVFFz6i5C5hFNIexPYluW2uTGAEk
aZoB6isBrW++FeQnFAgSFh1kJZevL73zMa7p4DMkr9Jpb899RTC//w46fNKp030MgAAQVYqlMBBY
FQaswS86+p6pB8wtdvVVES1bzFlO6k85OnMaAQ5DVGTqdvdyeXyYs+hyeML/9FVXCqesg+n8GBfW
WBxiqyF1pX76lwc/8f5XhYCS9O2+1txjRdMnMDFstlbV1Fq29fUlr4T53+7YxCXwqwgCC9CYHDrm
THrx48atzBXiQ6xTi8wkZKY4WkthVMeo9S4UCHjKZ1AdRVNVQ9F5KQIvoSFT6K047Q7BmUfeiGSY
skVQc7uT8turBCxKE70/02u/tIFEtJS6SMVWv628J5KQMYE+4l348iD3Ohkj5ACbRK6sTnSYBtqS
t65+eBJRX5GrMbYQdY81q/mJOqkzHGeOfoq1V2+5dDQGpipzsy+QSTB0uIDxxcc4HvUWvBjzRhJo
3JBQKkld2JG3DxacqsYCsJYCx0spxYrCOJAnoKMPpJoRgAuZhR1/fRC+bLTV/XVb9zluQrIfRUey
j+sBgVX9diVTTQyskWJD8ceWOGxcA1mFT17RrYmkJuoucCzPp7sRY/8FeH7pgjytaFaWsT2lbKgu
OwmrhVpj3uZn3QJ8BfaX067qg2gEDBQg+BYfoUUTdpr3teOpY/ytuar1EczomBFSSrrHLyq2yMAm
OAgy1AiY38FSxyut2XFuDVz4eatO2+0aMxi0RkecY4sMGhprXlVCJZYyCAoKVelILp+SzTynWE+z
yyy691je3MF3/h2GBHa8PuL0Cln5eVDTVKK4xxNy9zACwZpgz/A6ApIg304+8J6KFP21uhVPVcwq
Rmx3kSfAL+DzSbeSBiLv3kYjJymP+eF0GJZwz1kFVmzMyszjoSCO89Y8IDAuZ1/Ob3Bud4WLT6WJ
P+ndEuxrIOC2hucSX6lG2sOAOhm1MF324Kt4kq7ovjL70x5+TOVFrGZx5k/I2rXZRquAaQt5Om8t
2BewDsR3txkGRohGTL2uXtabzdk2M2M117LknqXHUqHIBhujrI+ltY9uwyjnNrE3n2CHkaFif4hr
3H9jnWdnPJ5pQj3y+hB5pPJbrelKsNkLUkPyf3AQiYfnQLaM0dT5OE+bpOzJhbdN8YHagThLNUva
y5TdPnh6QW6Z6zTIhheZ3EHe3gadsZLVjEvvdWFP1GJE0YAtFt1gPX0sulCjIOhZ7g7rq5NS1UwL
oc7bJc3ointWiag2pMDCDfHN0/+thd40MQhufvvSix28sBm9xA4Aq6ZxRpCXDtHG2AA/N4GcBRvf
4LObnfyjxY434ww54aKpn5oB5oJZg1BIYBFoE3mwM7U//ts0dV4DpV8+MRtSWkEZtiaP3U13mxyW
c/daMCHoZJtZiLXPP+3f5tfRvgcJy4Y2KwCVMETahT3AXTEwjutOJ4LaEXgZrIBZ4sA0dtvZ/ZWt
4ImyXijsDe0QmXnDd57RgjUoMz9UH5RqSWDCn3SosyaDHXSLmcauAhc/LJYQ2hvjxvWmEtUSM+wz
GuqJaChqGBLMeFee80EWS5Zj4Qw/yc2JJV4HbQDYP8+MzG4Ekuj+2PSTk3tiGVwuzVi7u7RRJ3ON
5WhtUmV4AwLjUMzYdcI4erhcHPW7xNxU/wPBsz6ej1Hlpwxmo0yulMgXfxuQZ7ohK6bSTmxyLSsQ
kQpzjtY8gO75KEGmt/MMXS3jBlBa53gOJCntLToiVUKhvlyeBfPJd5IkXyEndOYQfTo4xZB6hFOi
ZwtSN5XHRV51AfgrEX1veB9U4UaChl4bcZOPtuR6AR02wn05cUK2i9729LsktGW4ZC6KvTaHh8JZ
SD4tKBkPhousr5s9ZiwN7QQ3R0iTuC2q0vklU7FyECSos37ZgsBZe2Tz2lOuJXh4SwMhT/jklS55
soWrM6poanaWtjpOEavqmVraxbxAwPanPEtGyiDgv8eEj7OP9zvfcs8usNu2gUINcSZPy5H8VP9t
HZTaQAfKajIoSz1QEL2awlzR5o6uHaBitF/gTpfPsDeCA1C7wmQ5OooODUPgen32a+SRo1TaLw2a
S0mpP1YRfnJkoiFrQMvRpENwaA5LAgxO6J7WMEjAy4BUpWIjSkeBQhpZ1sZh5fDNe8n+6coV0zF+
3w/RftH0qm92E+r71Yi5cIioPT0K6RCO0z5jS/HF70nydsL35hKT67NPn/zVcOCL3RFaDlrmEGdu
RlG8V8CJbJqJ90gyTpQWxsj+BlzXakErsToTibJ3w2LG+sdr/+Iu86PT7o9P4n3yooZg9hwjr8Ey
3PncvAxAOJeeoKT3K8ijMrMZ6wmUqRW0kDrKu4Kem1BYnwSTxcWWnkiTeqmHT9QrbAhV+lRAF6+u
tWYylqkVyeUsP1/Ow1cpd92/diTc1I4TInSKT924Ym0lqz1nSX3HtG08lUTR6CyXgplmsjeoe49e
85cNbHSUX9ihe+q8hjLjZ7TIWcO6FAVgY0MuiLYWcn4q5Kuhl9lFDZ9FA3VgW3O2smwh704Yi7e7
iL3JsoZkd30gnQo1ruGYkGsqBTRSNP9aCfM5x8lEXqtXuQW5vEsJPDZKbMm9C5KLPWQH7yQMtVlO
KURtwJOaasaijcY0k+FILiJZNfGzn4o3xbB7MulMapAs6NmEmrrw6CV8eLo9gzuGLGQrpDeX8gvr
5oeBssIhaDqIjxjr89RC4+8sSYhiFiGQA8XLK97vxZMdeSoJAHiGGDykwZdAOR1RqaZesNqNcty+
gj/I6FHSO48UtcqyxAUFGpqIjjGbRTVwIGD57vFcFYmt/jbNJ+SerUTz+vFZ+lY9tz2uNBuzv2Sz
AHJn3KVHEYRmfaZj32QeOgMbWUpYqVmvw10VTeC1kUt+wSHz/BJk0dFxlAynUXlZ5824d07eRuzb
QLbR49azoKnPdXV7KE8oVKlK01nz5QHoVMtjlDBOwK6uuXAj1eVwKLl/TLOIBXCw5edVnN0KaTcG
1Z3SA+vmeOpN62YwrIElOag8YZnxzJDRQHLlFcYEWWf4ZdGwoamQqqjxvKv4Bk51lcGj3ZITIUE1
C7e6FD0PqOuDTYJvBDXBZBIpJ4p6fAmFrTVgGCvN4QCndD2UhDZ50WqUVhW1sEB2zmDPWB8ot1iJ
IRDC8qE2n69NAmZhMPywfW3V2o+ujtAzNWcFZHiEUSlon/y0d2nqSgnzmL/9ZUt+5xTbY//hrRE7
cm5bj8ctJ/mikGA4WEsbsIIiSeMRuiqk1K1YZpFgf8BTOoqntIy8ysBQEmwbJ+YFvBp6DBd33GbR
3U2fmOQDeAWg7SYsHl9womDsQC8HPAdhO3e8n9rgpJGEaAWOD8MoB8n4ofaYDze9XNmqO1tPejKQ
sQ5vE01BxVq67S7wMv+lWHPNpOWGBDBMcRFUnnJrfTksl/gNMNhCy+ErBlBlAMALSCgx0cUDUkKf
nVaO69PARWnUjpO1KzgPYIRX5aOF5p6Vsn8XU058QLi8OZR9V4mPld8JzfTmtPo0KNX/cTaaVlZT
fEZD/YMFqQcBgB4bSJ9pxnqIsQLjxq2exEatlPPs50KTu/PYIs6vqUoUNiUuAltWQl89YpqxELpn
2rU31FlzY+Wt7wu+11hWlj0oGDSDx+ocnJ/ubfsrJcgmn3TTBsJXMFmX0/35Y04h9XGtm9/MMTZP
foIFbc8Z49DNJjcJH20Zi34USRnrB1wARvMdkjywo8+ef5H67GJVTit2COtKIyEF5Asn0Zey1jCL
B+4Yc1FYBaI08rkw68vU+qyviiOOMRHYy8D/xnDZlH/gL/6Bzn0SeBIRGjyH2Ru3h5bO8rSV8Ace
7h7CSoE+ZhmkXolHOefIsPqbkPeubSO3kLqm681AGpTmZsg8ce1tyS62pJwL+PfmXnP/Vbku1jeL
ApKrdxFwB1VgBNKE7m1EIjnK9aeB4F+nI8V2b73jShp4DbpZTeGy5yedyA+dCdDVA1S22X1x0e84
aeArtgmrpFeJgvplCoAHICyu2DzKx0AAcwOYXR/uQdkj50ILdzn9Pr95AloXkq/AaGYI+M7d/dNK
kaTqiBhsfc/bcg25hvaVqXfoZWLx2VfBXwEV4WjWi4NuwBQb9yA5xjrlMeDRjUOr4B6zjQBz8vz/
hVfCNfm8XJr1JGOiEkSGGiVO6MeaqeASISqJQ7BT79jWZ8k4HqLqqhIizQzZiqws4uQO2vZxzNlN
c07aXNqSuAmrSzglLKjtLydmvf+zA7jVcPfTxWfPOEbsCabR1kcW3TS1YMopofy6PJTrqeqsJWpA
Xe2XC9Hgq3OKL5SagOHwiKA/qxoDiDnGFvEXPsR+uya1Tvbn3K0YuhtBAnNmLQbD14/KFsxG0E68
i+y11vY4bPhRbwuT+a5I1P5mnx620gYib5UhVJYfkjnOxsx9m+GW3GB6TllWms8xzOHYexTbXlRg
xaix9dJPzcDmG+oHU7ypUIWqzAI/zUTtGLVra9p2l19SbAP3wou8jKEdmxzKY8/Yf1rNJH3r7mGX
OcRf3qTo/3lK7rOtGDaMsnce/vJrKK53tcWol+qgm+xZCihJG0slMAYW6umz/zefEGhX/VHF4IaF
NnBPxCyIskmPdD9SdiH30sP54FtXk4i10soL86PdjYyhvQHV9/E9BguIJuJR0EQ6kQ4priSOuMsf
c34EgKXTniDbREF8JTjYu2tZsxIUQI1fszh3/uGf9wwPefKNolFaxuf4E/rGtoM5kP24UoUdnQA4
2Z7SAZ1SmLvwMp0KuKww2+JjMG5m/olpmcrBdSGgzNv5F15wrD7IjRFelsZ98kqFVIRVeV02aQ82
LJZR6qmVfn5Ch3ItYv0QwtzvCDxF98iO6F7z6LSN63UsGU0ELsVxzkqtTHoYHuXxgrc/VuVUfslk
iXxz1rhibEaULEGCVkTChh4Ao3IZuQTg7ZzEAajfR2vfGhZe08wB1C50IZmKedtwPPxlM1myzKX1
P0YeVTXtdp3kAbXdH6EyhARTL53C7aRr20qSRVADKs5n6XFLh3tYAOzMSqTwzkPEcM7Xitm9sV7Q
s+47AHaiGmv7LeWXm/SfxTDXi4xTRZR0MpIE6cGMpCXWcyljV2Dmus9TZuaCjh5H6AIWTv2kB5Eq
Ci2BOunzFVrY4gXCyeeDZXqMVbc1mjkmDtD83fF2irWH8TfsWziLn5TPOrQq1mDuVIxiSvz3QavU
qGMnFq0DEJh8SbkRGEfy/BLWOspzdN4BJXNZssc1bK6rTVXoy1JGRDPFPfSxMWT/+PyNa6guPoWR
A8GTJ2q0f3BtPvGIcmH6azP5YpTJzFc2IWyfu9bEd8dpQJ+D1mPSudLbVJ7dh495XGdC/aSjF4jg
cwnCoV1HAwTrbmvhZEl7yioTSznODvJNPw//+KlLnYF+0EX1hPkEgLBp9QIEfr0ZVhdBcxGun1bd
iMvFbyAxr/4k9TcNSGKHGL+x0cJ7WxunUrI2dZArMpobc/4hsedYycAqVPP8GoJqv2FQFajj8hlo
eBU8M3d7gbPvVK/kHbuSkbUtYdj60fc4hc46ROx15y0+66Gt2yBalYGhgrNNsvzW90vC3jzoGLQm
JvGJpY0oR8zTHB1imeTKo35tkGV9BbSiwbSPHK7Xg+eEijDhHkRP/ffC8A+MgH1+p7kVpd0H9tg4
hNMkLROd49UmWKBmIruH1hQb0uYXNYJGWk/0C6pqHGB7s01fvAMUHUheWVrc3zYOjKG8nt18JEWD
/W33iSSHlGqd5xOBA8S3zREfLK1BBWIz3g729P6GYw5xyWZlauest37iggIkGp+tGTmV8kp21rrw
m3J6Jc8y6xRVOIkKmXOTdT4Lnhu/OakGMOmjcP2g3vptivRVlQBpOKDEhfTN1wXOQT/DfZma47Rn
mTm6v9tMpTT0dHZHJ8hlubCDoM9PUqK8nL0900Y1EurItBNde2zDL0cwhv4QX+T1iF+tqtDIshYM
kN4Lc8MMvxa1PqkRcTgNthzcZZfUiVYa8j8s43tFqtzDkiDMux2BC7VYJLviAVhatjueZen53iB7
ADxCF7e1ANFGL2ubwd2Hsl1iZoP60HhffU6Ru8cU3s/QILJp5LzmuQLOrMZVydPswGto3Aqqm/A/
ounXKRlg+c59/blelQn6vhdhhdrReixcnBMvICcoI7/y3qIROQta3ZRqSHWRVBXg6QRtAwE+4Q2S
nOhgG9x5evTfC35JCXF/CcoPV8gXfo7ZG/YiiFSfX1yonxEwxubwiLrLCUK6kw75qH7bUP4rL5GW
DfDLTomJ71LUl0m1yaMuP3K6e+FeO4IqcQrcnn9XxNaL/XllRXbxa1GQtMMxFpkAjvFfZ2KCs6rU
pMU32FtiL7qLwJTXVA//O8sGKJkrYAcrLIsKf27PTrLYHXqSW07Opd23X7uPcpR2M9+fIKmlAf1K
lmTccxaqL9js+6o9Zxua6mn8654bQ7k+AjwN9hemLwLTPxwY6nqo1rUWzU/sAKd1hH8WzkQZSLgP
mSqx8Ac8k9k/anWv0LnGH2ysekhJE51znXaG/N0OYe3D2xyqVpCic84IfXu21RG1gSfUhemcq0w5
FLErT/ixcMEmG3x6nV/vT6OtIKnnMEP9bGf1jFkLN7GAtNIqZ2gQfcGeefHeEcRtHNiLvFrXkBir
cLVy0vwiNDqalQqFuH0/MYpztZ+6ToNipLm+PEg0l5M2AhjziETlxhbt+xo59H9YWDN62mML3+SO
7i3jh3eW3XoM9111Ephx5dpge+WiwTHAO7lLxfIPXdNVuFI1GQN1HxKepuwjIo8VTx8R0UZCccVf
7BDUDO403vRUnTJZ0cd6wh02NtOImFAzR3RezxIMJKn67aqg9UKYrPy54WjGTwQLFH01/tk/EQhi
osdhkSE6vCntviVtfntrSKRWG/DjDgGZak1ICzIZFkAI2+43UX1/ZQm/bUja6UVZLDJGNZA9bXMb
QrBDsCGtIffTd4dF9BDeDJSd7aIX3A4VU/+rDeZuUYc75k4eJHAzX1LY4YvmjKLQ0daSfbz55An4
WtGVXsZjZwAY8hYO83HO5P1wTycsyb/IVSwpm1OwjjIyyiSftN0ZPTvcuo8iFnsOOWK/En99rg1R
6JFPu1BPJCQkVzdLRPFSzeqA4BXRPAZKIQXJ6DehCSGd+Mvf8xVvfGCLSVx2V1dL8rMcT/dT2N8i
UK/BSfDtR5EPLlnjg4B/5ZTIsnhIqgAoEU7YQma9RKZ3AMh48TIitf5WGn7TNGq6jxbGxVXrxYky
ukwGBDrGJEkZldWGeUoAqWuKQ2LjYPv2NLc4oVAbls+r7FWNt4U/GYRdhK4ZDxqN0UQd2I0r/rqa
kijpJPYUKeg/lFzAl7M1F7GJUX0uPOv/YtaGnFicbPsrF5qnvd/uCX25GPEhtHHvH5oF2oruJuGU
wJ9hhcpU5+eON7lSoaGi/3V21ZfMlo0LihbK3m1p+/ByIHtcAnHgw/pEU/Q/Q7vvgQ1AaDV8ugMG
hqxqy3LUujDmliPCrJ3sy4UQfFSwC9L5TOydRn41uE8wcLLZi6jIGTki7Ov4DQZMDeQQzbG/eCgY
pBxO2A9nNRKzvaMPqsByvMz/n9Tsri4TsyULQxVsHfXBztFepGAKuMsIIQuDhVHwBsgZ6YIXf6jF
sIuKzkaAu/u/r5ou5e6nfAfhgtiSHHXgOUTQgXBrU7ii4b8ug5VzNnFlFdKPo5bLorLdF55KUsgD
S05WhTrd0vMnFWGfI1e2X5B9MRJBIoe6Wgy6vqHNH/ynZEbhI7FRLUNjfLJNmirqcoWNU/PLYqj7
4BHMFiFXqhViosMJTMlwRiGmFFRCoP3IL0GYU7QykP+YB4cqO5K2/Yz9TMWrubljvFZsiWhLHB7d
HdOMN2ShsUoXUsxQyxPMJq8dWpqR8/ABOJgxbfK0m30xsM/dQ+v4YDVlMhZaEsCYKBi1fI88jpBu
FY5f+zGgnAKHNhfVwm85yQbT8DcQrKVhAQHvOgWBYMuxVCZn8gijlhx16hATq9I38PaCwNe0K1BG
8JgnX9UZNukqYqSnyQT2B6ju3v56FGivypW8RuXOMJn4aM3eF6kGGaZX6tgUnHnsyxxbxv+GZRRK
13JzilQAKqm7zvpZ7WSkT9GKZ1hodXBkAZxAJuhPPA11cKRza7XFBwtsbm9YhIWaD9rwtDMpF6F5
uiQZrsBi/F24OMAEeXZWdSn28QWsRx9BprxDsgigpYIimJnP9ZkntQTBUGlhRiNrWKm2j4L39mxh
pNX14HemBEwX3CI/AFf6ahWqtsnL+2a/5Oy9EqiPt+UZPg4S23RJ5723yCDB7TrRVOYP3Zmj3W0p
vodPa6Ad9OgAeMO3TNkdfqVQtMtq1sY4+Sv8pe3oMlK14wBwx/IB1E/ogKPLE0A1QbX/hd1MIfmj
xd52gJW+0zKb2Nw7pkPEOzA0lBvfDWKayufAWh7d13T/4cKM777JUs2PbhYHoMs4nnrI3s3femH7
25n8imIcf32Pz6EDkKwayxTnyV+qwlLeM48bNbe48yVfe6lVfCJ0GMrxw7eZUWyMigSeq8NBPxGY
PYXxNIEFXwudWim9+PvBfPawB8Pe5k2oTTQO6QW8RT1R6MNPabuBelyGyNhCjKSO+a6aawffOZcw
6clgSbAga9Zw7QFUdW/VhjMRrRGntt2qziVpOp+/6+lSvoY//uXWoNkYDjy5yGtt7eKVOWmIGCw4
GJ8JkoImHc+WH2VLPGsKAZPgSrw+XWdtP/wnV2hcERng858kILWTmuj3YrxMkutsKFIZIUR8hv8I
bkT3ON19D3qYFHy1ptczPpKOny91fy+UezQvK0t64hp/XUmMCRtKeWJfMNXOC1ElDg1SMakpHFnx
RySej5fxgCPDTgCuF44aeUGGqv1xqaaxWfwiCA5rdQtF7d0ZbQFW22iyCrLsBhWb0ctEKDATVhs4
MnPUkwsmdKR5Yc2yr4m/QYledHLBjhswYO0/OatGxB2w1fj1EuGY/VVYmDstDTLNDSiLYWrW1pLz
J/sqCei7aBCUMFSUoMOpo+dqNBiU6NuRL2oYDrJfKQ75XfXBU+eo1+zYwGouPO7cCwuQBX2/Nybm
zQlgN1uryqqSt3E6s4xpoz/H5KO1WuS2HxkYSEgTH3P1EahgJj7U9dm8UUj6GBkoR3pgyBoZubi7
X7F4+3NYKac1oVv/KfT4grW7PJZsFnCroBZvg5QVtGuAb5YjoVu1gmBaq98kWBFTXTkf7fNLVBS5
C1geS4D5I0/R5bnHzHQ7M7UWZDc12FVe7uf7bIajWl5IkNtkPsXvzybcbWq1BZMCRkCETlHPSOIK
i8ORVxu9R2WYgQa6Ghdh/UfiPU509L0HogC0cohWkKiFeOLE5Bb2Ok2UD7nZeBjJeC7dXNYk1eDq
h2NRCn62mk/yITWTM7HE5XKw0slMgyP+iORe4nWrrxU5K7ec5F+OQBd4CISu8lcbLVLmZ7mLnUhV
6R7ejas1QuSNW2Krch+PI2eDzlDruxCWxGLxdypfwRsGYksDFVdYeF8CRBNDilbQ83HHEAfGvfjc
l621bFJC6XKYWTRyNyx5oxsg61SVhCdS4RfWT/toWKzuEcpzSPPHkCqCMPZt7w0EZj3b1J/FkEXD
/TEWHzPHWuS5o4B1uu0KP6muuwWOsHgUBvD8jYOTJqLtNlpxnPU9fPsfvvnFVH/xyKggv8GblUx0
rYSMWIgmBaR247IQ1LpCLaPctVGf9KVBFKlYfv1SuD4NISdHJoUK3ySiFCeFKpISfAfJEj38HD+r
YkrWnXvnQxr1R+c09Wr8ub3GLVl3hYsmw7lvOXCQhC28WwVGssrngiOijX9fiZebVWrupLfyKy8B
XKhiWoN6BDJgvidGdT440BCoomnUKKtWwbtm4Pr8pl08jFznseG94Mk+slYu+WFl3dlTz4hsaSFt
07pfrX+DhyfgDrqRWv2lYUO+8JYMCgzJsz0ASqylm3nMc2QrnnB53P2NKMwtzGS4i91OTqrXviaz
noXnBuqrAMUzlddq0bwTHqc13m8BoYSZSzTvlXOE6+kiNktleMYFkxiQUPnlZKx1VtNbW8aANeEU
cCA2GbPVEy7GsZ4UNWAnt+ScpFVTtmSst9+GbtFJ4H/No3chbSmOhAZFKaq5//Inb+130/pqRUzi
+6rsMMqx5igqmvdo81yEejsRbIrCIWjVAL136/UoXDBu5be/SYYEkv8Hcux4PMJZZ4AlZFlxDN5U
MldbLOpYGhiBm87qG3Ivi9/CzNWONpSJKQG98hyGkc6rOj24zCleoG8EhZNGQx8jnsIk+71yFYbQ
yBSnHhK8GdTXbGVehUhAGMDyqq0IggSH9hzoaj2ajdGW0Ufd7Cm2rKn5kDqgXrb8xov9qhdezKVG
Ea+MkvdquazXDTkef3+7AhuZZeq2EmwTjjAZN95xmBqZ0j4KEzGCfgxyPMpaN2sb85FOGH6XYz0B
zNhKGIYZeN4jRZ3C5wGR984IpPhm8tLlsmEgWDTWBGrcyTFXWXoF3MuLoCIwBgO5uH904Be9lUUh
LUizyKWtKxs1YInIi7PQmXaFo2cGHa9I3oYISBD2s7mcywCq2o+5SIXmItfBI59ECs3iklbMPD2J
l9VErfjqpcOhm9hrZM8ePhmp2icNNuEyDALIXaTGnv762pku1HksSEYfE8YgCMUSpxKaWjXdwi1H
q/uLBtZfJG7CPShR8mcZKOxe2NQsOhIhg1ri0ydIRc5gzXqkh0+t1gwuorAL644O2FDzbZ/Bzptu
5uBIVq3lb9+SMakKQz5P6FjPvLdOwBnkRz6WpMGtqyqV2EJu6xwKFG/6AVft+xz/CyIy47i6K68V
+pfOaQn9cjlbHHyNaC0gichsyqhLqmNRZgCF0BEE5z24FePz6vZSWqnFvM5UZo+TA/HathU0mfqI
GDGL2VPX/GKcuCUvufyS1nsIDX/PEiPGg5wHu99/x5xsmXnGZOCpIIl651ikkcvxUjsX7h+xeHrC
RH3/xljCE/byy9CrGelVLtNOTPXLLQcQCECEjknletAKr7ruu4ywoBbWHe94o6j/ewVTLXUqxXJ/
BlgtZ0KTe9gGHA6ZJLnFfBVPVbwdO8W2S/UScxYWzH2EQBjGpfEtht2SJ6Be1IVgvdVguDfT7p6+
5vt/Q56J58LfcSi4G8BQq+ndNR2Fm9j4nfMcoblajXOjMNfIDqjlYK95MBpfP7vPHpEmTv/bHsfb
f/ponqLfdmGiC7EA/GQDxvRUHHuHmTzMrIhpjoDa+c/AYEEE5hRLoyIBuYfzrpCajTd4pyvo4L8Z
k6fUcJEyHQu2zNraYKQd+fkuZgrE3M4ANMusLHm7u13KNJcJFeeuwFmj+yABfCdWuPat6t/5dowF
Fw2JQDYadYWBR5EKJgz3VfLhzmSkkFqY3dZSW2f6eoaucW/HUIXbTSbZhsn8aDD61I2wi/Sj/0jv
NYTgUYVB4ophQMV12ksYT7S4DWdLMmqjf/43IN1ocpc5/oYCSo3oHXCBaDrV5Igo23wWqYgWU1OG
okGw8cvWsK7eWhYnp55nbvL1dBMjsaISLX+B2bYrAcZtxJVIz6H70w9iRwQnoF2TaG9n+wCyZrWH
qpt+TG73/cSf8oIV7hIhbZc1UntXx3ejsdxyVhLUTBI1sQ2f3qNh2E+cg/LoiUHprlomLCk8VGJt
3hZiUYRli0QSDuj0KsQpxr4fgvuBIk0JSLmsObK93r7BHmyKpFtepjy44Xdk1QMNOwjj7EpqZJFJ
dwT6aAzeQxSsTRfUrRPibSE7gyN9Pxy//CLp3+BLH8ieqYM8Y32GrfuAGhrusOo9ZJ4oY4LHnpKf
hLny5lYg154l0jsG22iFPttEALwAo3xUHEJB3iUgKdvz36XS8MPSqxfS7QgdOoAnvuKJYcEI8hRF
iB8+DONQQwty9U0IgPWQ1UyGxz5m1nZdvCGkOfSu7yYVRmzX9QsPgXJPUqdVoWDY1Shv3+Vg1DSK
0xA5IU29Ww+onIB8xIQaxnPoPZN6/nIXalaXpCO8L1lmREH9Kjw3yb0wtPYBbRNf3iFfstspDFWj
zBx6iM63omVzLj1aUrk1Ni+DoOZTvzAkmUI3MuLc+Wzg6HMPKXnXO741ea+JNVulmdmmw1S5A2le
LDxYjSTg2wENv3V1p3zkf94UD0yeNX2cnEBFxpY3CF/nqppF1CxrvmmcE5Nwh+dYNIgfOZqqpBFK
alM5uqTyu09LFDUFd3A+KG1SAHmD5nsUj2m9EdS7NoykchXRB6gpjHfNdIH3VH5i7DdI3ZdVCw9/
89SaZNPJC9JDyQe+5PeMZQiYFB5cuxnP5tX5Q197ZO7/Odsw5RoWGRoEB5dUz5juJgyhHWQjffi6
KZ0XtsTOHwqCU/SS/0y38p70+g5mDzvNPYvbVyupkcR/1eYU59pqjIZihMQqiRWqkCq8crOabG4w
LrT5t62ZsU5Fv8+vgHDU6iAaQJ0m71+n5D8MK0jkJbyYaVxa3nb6JPFO8yr4KcGMLM6XQ8mBmhRi
N2CSQ83uFYtG2nGwNSIK+A0DFjBTy7fjh1mP+2Z9ZWAgKlsG5BayBdqG1pemNoJvQ3Ef6NLNqjYR
nv74DHCG0y2yGGIZP4fpJ6jCwjr7vXvympoG3XjarWpzYyHJFxmhrJLTjYS6kDSglwnAmZOctQJf
28Ijr9Skta7KIqNqk4UG7vL3tv4WVyEe20/MYYs1q/ZZgfLjxrHexBtcaGi9vgiTngPeSXmSbjEV
jzrN9qgUv28fFUXiXolVU4qMKjBNTuHHqJa8IgyNxYhQZ29PqFhANdmnJvN5oPEaagiEtABxvnBM
AviXq5uvbg8uR6k0BaUb8lPr/CZG6m51+U3kEZRY9/SwUyA8gLTrP85OJRQrw4AfaCPEB+dRTbsx
Mx0619bhAjxAo21phjUKVf8xgKFOzzN1DcuO/8ZDLNww/p2jZXdOecBCHuItFjSErpGPfNN+BmJc
X6Z3ow+aF8rTcP0zfodIgFp93YWNn2JH+iuAVmz6HvFb2VuiAOX+sh1C6BmAPA4rd/P7zCNdJO81
BDxwO0ICUzKbWkzFo+Ofwj9wqcm7emEdI6yENqqkuFgI6RwGDgrIZgl7iMMLQ1jNPp2/USQgoOEH
nq4NB0nzkNl5TKYnEtNoVQKTruKVFe2Gdh0ZckAG8OoU3tusR8Yw4uxIRAqyf2Hsm1vmDEEiAUDm
mvFEozWOs0QNx75I23PXlRCT+riUIFluDmQJ7PZVlqrrJ6yOc8D01FdYQtxOziuG2oaKV+wH8BDD
Urtc2N9lvXE26l4fsCLB6vijxVNY2zTZGOMlQ7hIaQfzFyfGlHKgiF8r3Km7x/UuqrE1uRvaXE6T
b9jTpdpCRHEX3IzxuY2EDH0GE0VDlY7hhRW8L4MYFJyPKTg0YzaaGhcojJXLOqCs2agyOYlkYIY8
cVFzz2mBIuGdKIjQb3x9gcUa5f9WS+amekjJQ4Rsh2I2LjmWjlRqd8In8YaGce5Px5Vqx5Plu/2e
pYRDatL26TTywRL214qw2DPMC7nd/zv0LzW/tdIqy7Ex/0tWghJv+EjFnFQz+rVBdmVTBJLqY0hi
m/JBhsDV93t5ZmEcLHmApG+TVYGTsIigWUjeuDqMlI09Y/WG8us9F4WHQQ/thlY4ofEGuDdh3BrU
FMbR7BHAZTph6/tgqFauBVIafbJkqSQw4/tcQW4dFWAv3Iskrgi4LskV1VYtmDjPLriu08SuRFg/
gxqsPTn8p1uxbJ21YDdEqjv0arcok3vAh3FsKmGAR7QtRBHg8gIk5dQqpqHK+y5UH4LLCegcUvJB
63jrDLJzT0h4iHM870vAg7XokgDH9y9deYArNCvky5Jr964u8tvR2VVpwT4o10g2Uerz5apvpU+R
yiDefHaKQu3S6Izirv9K1dd3vZOLGhVycIgg0EzK3k9MToLH8BD8kaW38CU7IZhKIVwNXQlkKRNq
fnk6EvdF3roBJ0HYiIadT1IACcttf/gwsa930P7U7ii3mteKHFov99JK/Y+lWjwCXpx0IKilLqPo
Tw5jk+RW9rb8LNIKvh4MA+JUvipV6gF1p7PAQ5M3Jz8BzlCg0/Ed5aPybyOznHOojKtCe1fhoFQK
gnpnQGXWzLP7LnJtxg0SJpaWKr5Z7goXin459ouTSuCqpJtkFzWaOdKSIIjaLGPCn4NnQgglgUGr
V4xJtFu030Z96NZf0pyzc1XX/OM7LCDaS34tN84/vdtvaq4ZMdVZYytktqrApKPkslp34yCYVA18
ogRAAg7EAjlnlVxoyxGyYKFEHSQsAkIsUyTKsRZ+dPBK1EwIebwuMH49y5CRyqlAXsmSHXxOEZJV
3apZRlbPb4gQco1YIaFCiHkgUs3B/pj0sJQb11VnZ6RXsaRIOVCfdDqiI+MDr6eguAD1ZyAOOmRY
M3L7BVPrF9OK0oUgf20t9Y7N2OPurWI35D8EkVVyYirRYyP+ft8t619pHWFvXEcL5QehkLh+bTQN
FGjxge2ulU4b9FC4GrzoPRqlm9ra3wA7OGbzmEky5FX1grP5HUWZWGnHlc0aKp2pA7IBaaHtiBdz
6STGeiA7oWV6nKD/NO6BsCsIKJUKivqNYdy9d4xfOVZiDuOHLd1s0RW5uuJriqRtiog95bEBe4nU
DQzQ74Krc6o7zVcOGDzyOdhkYyYdPNmE5E0d4ADVqhLImh1MW0fC4NorEFS85HmAWdqAVPqDtpa2
6PVpjlCspsPdcRCeS/RXIjJNEI6NJhjpiBY/1DHvkhce4ywfX52ggGVjzZKrk7/Yuz6N8OTpx6z9
iXmp78yaHq5a+Nw57P6yd49PTr5dRNhgC+YydyRmPFdiSWZDogvyTc1PliyGk/qy++Rgc4XEGnay
ZuTmqByDPb3kfkuoJTpY1mhCu+kTaEwF5znd3GHNZjfe908y2iUI+QktA1Q+mCfYW8t9CGGK96vb
EYcxYVbYhMS31ZLk3rD5XB+K+qmESmo4xSPKrjUxVyxBWtXVXgplr/z+VO+JOfBdplTDCx6g06O6
fhdb5QozRPPiQDuBf7s/g0Le8td5IQrNG1+dPWga7WR5WPoGYwj0ZjBuS1fCfoVIKx6+RDfUSUlP
Idow5+1j8KjD9YRTtBD6NgIliu2HlgDZ/t3qygVA635PmzjNxY5ktifcKAx9oLNdSNelcL9BCU3q
5XoZNS/D6+v9ww1oDTsX3Tj9GZkKor9tQeuv7db0cAG/rHjPCHZzjZvUKKmaIK4mX7gkZ8zEemzm
Ry30Zm/qCZXVelX6sfbVq3NhJ83g6zIuIBLiUJJK49iKSEr98pgUgdnFs0giiuRcmOTR7hlKgVqY
kB+I8mX+8H/sNFK23q1ejb1IT7cHZ3DAUBPICd9tL9sRYzgOQ12TIEeR/Iy4Q7JFT76nx6FRTp50
2Y0/8JB7gAU/l9y5VfCIW3Gn/adbOyx/QQjaNnv9MjkBfUAIvTJOJURnp1HVuq7ei33SUMRSAnYj
+VuBp3KkF6EtLIWQVA84TheRhi7IVNC2rvDaj4dvm8PMQ0bIqxPR38PrBJUixpcxUdlAvMXcEk8Q
U6HN5XGsAqYVNCFPqKE3YN7n9akMw6oFIqOGvVKwZdIuV2NPqZDBSWStyFjVr8pCxXn3CnMwufCm
5zh+wgA3/xef6uSINeG8kHUBx3mPNzGY1sQlvuOHOHZhHr4lzXOHH76vyQ3Vo/vn3ymxeafpVE/Z
afwYlAwgytMOADk3lN32OY993amwyT+TSz45Vcr/lhFgZ5SmtF6xqOd5fQUzpdejdQCXpdPStgla
sMGpHtKxDXW1BYQWDMD4PUSEN7WUcgeacOE1+GLMt6ABvTIpvAShc/SrJUgO6nMiz3mPHHPaY8Ef
h2P/KevJki0NVFDhhTLdJa+W74O+Toa6qJs/IND/OC2G4BXvpypa0u0yas1uqZLrOgnWi/1aLY2a
sLJ1ov3nbaSxsD55nLMX8Q/ULQ6zX+s26XkfWQWebxq+yZJTej6RK7pKPTCLaNu+nj0or+0zI2Fx
+vcE8cjsPC0oKB1OB/bEb2r3If7WlLPdZA1oaQJ1G9ToRBs1W5yHhiXwhip+Ar9KZGp0MyBa4FaH
pTGY4JURbzzUeZelE4KIjI9WUMCvZZfX/zQ4kSjxLAqHIxzKfWpXF96mm7D9N+2RmvXF+s3suzek
H8NoDNgMTHymC6s/dCuTCuLr1s/RhG3gnhVQg48wNLa+TmULtD1RHa5aYoF4q34Ru37FuEH1zJJ2
SB5aMOzHIts4Nxgc+XlkfS7sKwcZsdB9MNtEL+zOguxOYYF+iJmo3yyU2qnlAG8As8y/kwmxTP3u
+kF8VsD4yk7WJFceIjuyR3IZ9trLOh7iC+IhpYsX4rLOisM4YizORWv5VcSB9OP6G4RTr4OKzULm
HngvhL1ik1O/EMQD3qns9t44LCADx49X22EfF8ZoFKW7cp5IN0jZkh9ixvBkF9Wm5Iz5QsUEKzVU
UHddHPQrEJGI+6rlN0xmSynHTnGmzakQ7EzOA6nyV2uANaf2yhqFwvbYRaoN12UobINjAHljEkiY
PqaS0hR7YzM7Ud9Tr16Jc18JFFHgm8gt0ODMk1jEC32ZGcx+OZd8coRC3NdigsqA+4M0ydXrXgNr
VCC/LvuYC/Q38/306N9CWlXMp0howLcCM/vsjDhGphCeM733EBmWjTCfznOl4L8jCHTqDqSxaVc3
jzfTmHtppZVRha30eGtqzxlSC8QNkW4s2wk/wZLBud7vCswJffIPsBHsTSk/TYw8/VlkVWD+TZK6
lT1/UPTSPfmsCQSiTeR+joKU7Q48o7PxUHLwowBc5XC2WZBH9ZK/ntV8xkLs2aDwnxV9xhTgpgUw
ggsedwS1nMSSM6DD3jIqobSoKbeML36ieKhD6rZZUDP8guIwFhEkMvrpybUka+NhSJDhTR3r+rvb
c8bn/8mmtaU32TA5uzgNRZ1bGmGLGsTMB05Rvpy1H95mI295Kail0xYY6fcIyEzx6uGvn5PrA11L
HBTRwTQ3lDzB6pO9Ovpt3EvVOMWaKvsP0fZNIWiyjHVOJ9BU9xgzR2hmzJ+z3GsgXw1kW7yD2L7U
Eh9RBEJX1/emprSBlnHRgSl6WbfWR6L//I4BXJBnOGVSo9mevqCGaxlLXRDDZoG/7nMKH8RApexW
NGLrUhtmrAg4rEwWiQ6uZL1hEO++mem0bkMWZ6Ri4eA8oikFkgYgaX1+aglGErw1teQ6Th00BIos
yGrSudpiNN/mDOsqlnMPWkEZp/rI5KtGgMGHGsNP4RfIuqrbEq2w7agUDzmkJmWC1cMFaP6P0TDv
ZTrVgD2qz2fV8xBRNLrELlAengK25Gc+93mGPAB35asBFirW6416hrfTTCHj1fE/raedOOS3SpJU
5C1wwV5PSQ01za72VGFEUBwvr561ja0+WOH9KgdguWEnrh7uC8ntYXV/5K8dNrQOKM1Ytl0ooI8r
VCujvXRL6snFYqWSu/NAqYUyQPpEI0EeHEXtlmLYMSKmz2NZyH3Q5pmeA20aB3sefUv/72SXoeQS
MD3ujqbS016gshTQK+hyzszwMN94FU27q+LUuBbJqlxxGpqH7om662tdGyelMm4/cGhsdqMEAGnE
hyBDLqQnv3ackur9/vxSEIGjTz+QZT4b3TyxecQisRWwqbHO3ghajozQJGlmIZT0+QGyZkPRKdOL
WURnrM2IKQZySe2A4d1MtFYRh6lFVXF7BU549SkKaLhZAfuKGsrugNIqG6w3X9Mk1IDQiUzAYuoD
EzRRy3pgbt81gsiQLYqsBwx7iDYaQIhy6JcAPz1ztjauKldIGE6pcB6bGbiM6lDFHjbnJH/oUwIE
Ldr/u+4/wZtEaUXbnKKYzACwg0N5LN5K/3rhFbkXnpc5S6z2dcROGA8iruIuMzlUUgGuJ2zIvs/B
+IB/OOZVPenA9M9+1aL8uW7aloVHiyuQwBNSYsChuN5HAKYEyEzMoL2xmaTTFwCTPqosTddrYRTH
yq1v67qS+x6QsEHDTQ41PLZnyx8jJoCOsTXV7xyRL//86+aIh/2sIZ/hQGKV+l7ARN/KsXHMQELH
q6RM+PObMi+fyVgxF3hVssxx+w1DX3xiEzpJ/qbYgxQnR7NyjLwPn0KMrobH//FXoXIrGcePe9JO
uFrRc6EkxMimVKy2N6A2hpwwNsuLX1qPc+wertmQjJmrL4/Yr9ycyV8uZ89Uymv4cDfD3TPOGFvC
8/15vd0NNJSZqdfCEEY8ojs5gTpyJnehA53SxDFDlYYBH6iZWtcOOstO0L8r0nls1d5vA/63RMgb
czhFqB5cOeGaWDTlcjH7sWGy7asHHp/SeAwB10Pmdp0UlmWU9g0VoI8+G/fvo1IVjy6p5ze+9CNf
KdFIE+OsiID6P9ZIWqNV0H8ULc8bQbVjaaENiEDeZa6sYBXbXflvX3n9rZK/iLMCqO8x7jUGBT2Q
JTFvAIkhIXuNnuBK9E9nYYeCkpkZ2pIBQiPkkTk7tupGI50DRHGJxduuls6ydXaJQf54o8CsYu1q
kiSIPC/+z5VR415NfCjkSYcGX1cd4hMhUj6PnFexrB/Y/GQVgvOGNogpKU7LPgMfNu2SjZ6yHB3I
L1oGiPV+4hmNf3A7M7FZqHT+EhlGbW0+Zqpl6XQ738/k6pMvOsUYtJ0wrwLl0/FNUNd7d2JdwvdX
jw/MqbfSSIvTNFUKkC9Z5bUDIXTaSiCITN9qTOwb+dOzdFsE2wkRmn/WayMQ7dn3FzvA+G3h9t3M
GHd+1jN87I+KC3213nO8pGg4RTmywDlyV5fr2g43WitLi7sdxYhk+qlgxz7kRUcbl7/T4sZubqkF
WKLJudkvSEKPd9NrkP515EsK/sQJooH6FGkkmNmvI7wn9SeX1vh3cDpuuIJ6fpMU8nkl9J360z6q
aqTk7yJbAy2JrSR/uuqGwpHeMLrdvbG5iG3kRCNQK7RAvpTWaeQJbPjRZzHEBifwNyGb+ZljVtTe
wSos79qUR1w8064aveJOhoSSLJ+8Dj9S7BnY8B963XIOl/Vgc04uJvfir9hcho5Ya2dgZTQBsoUs
oChGV+azZT15BkLueoCUfGAJN+Sz/HR3TC/bXB0leXd1jymxLO1hMzvmS2V7PSQ5XZi7QMlMoIgS
OmmWjtEBW31+p1dhdeGzP+Sy9dQ/32Vora2ToBhC6VkwLYvf+asLGd+cbOa72nqWurH+7bhl4f/9
kD2wncnZrDIcwCBRaz2ZzazqIPLhxu2A12iPmLngyqrV4G/vEEZ1U6a7EYHApezBNzetLHSSkBZc
RtznsOHoBUhZA58mXyy3nQDQSC8Jr4FjbZ8Eexy+frW+HuvH25LN1Gae5DanANWI1raSxaQV9V+o
GHQYi/65w1Wgajv+2X9rfMvpu2UeYcY70pdsqc+jf3CipFObGHFCyv8fVEBd+alI57HNEu35v27L
3Yq+XFP1YV5EO3Ah+zwo+/wfFc7tEDpIOpgyaibi/3WXNtvJYkVGraPVwEUgBd3hYj43QLQPyefb
/JmDqz3IyEitBXb5SdiZMKYwlXAHcuKxq8VNTGJFWlNau5ptdzdDOi0SaHzaeFY31tt3/kLNLXpo
c6Y6XjUJ/TPPHNkn9H6b58EAPRxHhV/oPPmGxEaR6gEUw14nvH3tODo9DTOeVV32dkU2U+7mNlpI
gr02NLZLqRoCKGu3zxlA2hxS/W9c6gVcZFh7IwdRZvkNfX5k+yLg4VuZWfhIm72iB9qCGErkWn6e
/ivKA/Fk41RlSGm90pBVlH7NMr+Mx6t5juF4Sq5YFrOLJmpDdzc0B3tClHCYkXDKP/TG4JqHmvEW
5uaBr+i1BBdzveALh9Fdok4PZF4XjV3mVb0/r/g4O4lCJQNTdgnSHscD7oSaVgVlXo2Ck+KJ88jI
BMVC50/FQ2aXG++Mc+Sa9Pzf+WxsziPek3O6koZOyagmMXrteScO1NgQ6D9Bwpl2Qp9WfV/m0ZXX
WZD0ALC59yZ4+BmPk9CMx9PzzKbj3je7+HvEZ93nhQMoeMCSUynsC3rNBl3KeLxJQTeyfOSQuc7l
5x9cBDIivCrZ6rRWcL+Wquhn/WdPxNj8fci/8l1NymS1llYeIN7gngYAUjbYijtw1ppdlBlXSgSM
GTtnAkmH0JLDnK4WZ7vAIkxeC2fpCFENYu67K6H9veRlqR+THAOu8mquSjCV8RmT3w8IKpk9YtYc
/X9k6vkPaJu8IMBNn2gD9IgjXqLaHHR1zcHBQFhtFvG1udvAZ/EniISLHINDkt8AkNebt9SrAkUr
v79NmYabBZN5sbgqXooLgc/p7PTi0fTXxnFVhzDFeAQkD96YxulYsH7U/B68FzhYA20G+ZuYjnrG
xv1gHS04XVjtzck4exoStIndK+H4gS9aQQLn4ITEeu6ynsVwCflxLktFHo1lj+Wv/hJlYmTiHBHf
LXuKQbMWF080s33XZuBaA6+O9MdjjBBQwSGv446r91tvaQLK8n7xHRFCrVEqB8KJArWBOTKoHKCV
zfl8cQUEU2Lr5g493cz+u/LpO7i+71ZvHY60JzZk2et0nV6AyvEFh/ggHkTFx1XcpC9AvZ6FePvW
bkW8SlK5vmyVXdQPGTq0+Xy6+G1O4shlWHnelll+HZzMxkJEBrnp1K1W6tk4CH24EFzn0/i/aqJD
vmc9IXSSembEdwHqkvCEElveTR4P9Gv9AwbQzVHcEVSXMlnOC3Vsvk/OWf4xlvk9Od1onk0DgXuQ
9j8xqVkRkxrMMb+2PXZyPRbKn3P0UmExgGvacw4+/Okz570YQVVL62GYCwy0AqwumYdZgyHxRFI2
hmNuTQlZ6r1+zUKZ9ErH0Gg7mOTvw1PL01Y2LNuef+yUaO5JqiWL7EuEEUwYVfd4WKTWxL2L+x9M
Q58xrUBGcZV+XzbbvfsRnEjMc/U2ExANquviH9Ei1DUormx7EjqqyqSLYVmlW7X7eOX8+mOdwTCE
RgzHANdDG3+voV3yx1h+4lxj01ksneJduOnR5GmWlwyI5T1Em1eNJZgFqfcwdIKTo6JP/YdVGbb8
HoeseOqLsS6if3y5itTL3Cy+KkwMeEv3NQx0+WbfLq6hPY7OTRYIckRtHwm1umsaxFhOTGrcUKaJ
kx6dY+dH8eSe6JhBPrv1pwWoNF1rk5db03KbLkRQxzinSnecqZAVyDbppOCN+j9UkNdWZrGoz/0q
G3VGKq3SMsERDZio4sqKYn9ENwjabXkcoLbXJgY4TUX83uPoe8Oq3Yv1Jh+OjaeeUGuSTwqFE6/S
91qCy1SFeFtmJs6YrvhozToIb0mNbBde4gxa2xH7okfG0tEbGgvdKdpvc5f6JYM7h88rm30MvyEp
dAT+V8p4HPrvVEjoDJRmehGWBF98CPfnmj53OjvIiASq4GeLSgqNay7fBhbpyU6lmlSwd8aZqoe3
UBHooWobMUhAqUU18O2Xw+4mO1dtBBEK9HeuxWG+cEmPohJbPQEfr3XD9cZmqymHYjoJjg3Aehcl
asUSA9VbV7q6I6lQFxxGkrEVWY6ceXXYQ32Q8v3fi9aVJh52Ez/5Dm6u4GKzirsfvybAUoqu4ptC
0m5iqMTiM6rQ6JbE0p9DOJf+rGSN06i1hTFL/iU3rumrAqOcOtBgqhXZacYyuvt2yjJIFX7ysLcq
hlVEzzyGV1aPrC9cKgDArae5c+cTuCBwOCL0hbBwRR7/LecWzBGB9LtFazaLf25gbjrMlqBolgn1
ToHsneG3nTvuvq7p/Rm1yBSxjp+C6SjDPDAhLl88ENr8RiaOqywweUI3fbTF9kFGjXZGW3Jdhfcr
q6XeTMz9hgel0dLDRNLOZA0Z2ZIlUpMzMicnjYkBo1bXj7QaPuq4mUJfRVrx/thEnZD7L9DWEoF3
Z9xZVF2mgluaEejxxiNNeNLm238iUKOxnbMRLXwqdZzHELQrzaAmVlI5hhHtMjBreAcy1lwFDpuK
XbzTosMAGArtrxTtC+n9RuEAj5EZ+jJLQ1VpRpcUr1OAUZ4+fw9vVqWTw1jBbRbyd4A1yq6lXwiw
FCemXaBL/2tTY8k5LRUZ3g/MMeo9iL80SkDeJxFPhwxkiRzFjk6PSVCtJIX4hvl/FIpj5/l9/MWB
nvMShwlpqky13XHnqkT2DsRF2s7yJRhZzlvOeJ89GfY3S08K6Vyw3tjhNRSSknqt50FPVwpFiViq
sFdKuTYrNtOmC364CaJFDp/jS5s6S1zdZBwbQssvWuVHsQz2z1DZYxMd1vGhqkzW74FnsZpIowh/
lybWzbyiLrbyn+OPF/7ZTXe9WvXCp94As2c3XpbFDcAi8fXG/QXjFUGCxIf3fj1vMm1Yt2Re+eMo
P9GkxVKQsqaMspF/o8xaLyBGMbWKxGDP/nIc0d4JVF1iuwEK+DYYyd56WDpfzYBIEpl+OORNt5Ol
uYSbJosvFaAa4kBh/rrlXC0cdXmfBCPhco7k1mpp1Amcf7axc9uQ2IDgJda+TCNvzXgdOCJFpg/2
5JnBnbcdBkAWptdFdRqBQKkZwZNDhU4sWXZBl8D2tWcvjlzdlxvvCnPXMRiUEIp22BuS+3oNjjDk
d5ytjnb3eA9GssKIOqEjWsV6UsOKJdyFlJ9LPIr/4wf9d8wx5X5QRiyZHxIIftuZZU1S92JDOO5D
1HN/7xqqflOiG/qUjtoyaVzDe4HABaoCEi/4hnlKk80RmTismWsj8+bqaKRzpbQ+srN89hohf1wh
RhXtY6t5tykj7nbCYw+MD3TEJVZspkGcK1ihdZlxOMyU/OKmm9j1yQ6vCZez3wcNpJC2n7jSA5yl
WfJl9jZ6FQk4MmRZht41tbO2y+Q4dMyfO9UW/cwj4AprKkGbQtvwOEJ3xonjgS7x7IEKlk9QQUOL
0KrvfjnGJfz6EZ6Fn5ohS+ws/aS0vDKlMjQ9Q/uA08bhOXNLVggjYUbFq8WJfMhpcEeszKgUbtF0
1ISoNkhb9HuY8T1KN+syvnXAsOaIULOHUCjkKV3lrd3Z3+FhF++Bta/Q/HyYtZF/ORIAYmD2cQDP
JMAuQ1QzJ6zm8ZRuLdNNGAZ+oZ3vmH/crRU2L4L4j1Yh6reUOfiP3cVxikpIYNs1H1gQdk6+rTz5
IX5RBYzrKE7mKU6XGgbyfX/8c3yCpL0vKEIdYtvl6ge89ns8ucxlAwEQdxVIOYMCK6DIfbYsSMqO
GCQGNGcvUFOEvA7WgY/I1KIAtMc5T71eNVpPnM+48V/uEtnDUhvxQNoqbabLCgUdx0y9Tghyvy/v
kAwLATl15yux1cZqWULovFsP9Be7c8WAKs9qrzGzmLpBlku7FYbzWYYbkJDfpwC/nAl5awz0Xi5j
i2Iic6r4ZehGjmmAy2xH3cZzesFw9djwH081E2/byIQEubHdTDSn3rMhpv+P8O5iKfeDWA/DQT8n
mUNQPj9EJFO2oZxwW6HXoLw4wzLttEGcfCX2VM1DQMf8nMWUs2izZggfAYd9FWUDG2eqkj6+NPid
Z9rL94DFYwXbt1iPWkvuF20k40XhSgSc6LOsoioAz2U5Lv1CAp7qxHKkxZfH4hCmbmILkVMkbfOg
dlyh07orQTt/VVcbytoF6sp8xo09Tcr9FBSRfeERJURE1cFp5n29j748eyg5gtgPnqxcrDijxTSp
2ojyFn7EJgy/mABOENxSol/OylLZGRt0m3KfIB11PpxhsChC0p879ow7apIwGnBvuf+yNgognDq9
VgjrWhBN6Tw8MvJVHMz7DjSAg0tcVCowzH4d45/CKWkYQsRKvP2lGw45JyJCwqOgIpP+SqbiTT+m
x0Vq9xr4x5LhiS+3zbD660NoLW2+2pIf3SzDxBI3wWdx36JYGON+0JnxEdpuhFiUVgefQG1ez5r8
zgkaVbjgrbCXMZUHf90vxiYVSTgci9otnLsMqxdH2zATrixttaBx5h0pYcUHiSLV7qyPdTmeW1xg
e48s1OUN5z4fU/2L6KK7YopYUfiGb83WUqtTwy8yMRqaua/KXSDXRC6abKwChZyhoKQa/FYjxRXO
tD6QbvSZRW4Kuj/CLMczWyPU37elktyEhzwuqOJ99kO0Ma3p1ENGOP964FQ6i2QaG3gYVYtIFifg
t+TSMgNDqVlM6EZ5GD8v7txRtpdJPTpYfmxRV+zncvRVL2z0fg8ILgs/64c0vXgtcMpns18lUZ9L
Wi2MlOat4AGUScoKsZx9ddyKukbC4v99C55mP9+7f7Xw2RFUIPYaNnpyEWXVZY1QgSfxHnXrwcRm
JlicoyCnNa3xiF3iwgH8incRQGj03MFVvkty+eAb7JSbwcpkkqLHf+0c2l3MBNF/YvGY4UT+VwZe
i5wipqmXUKxL9a4SdQbRyTVCQcHoRODJzqKXXE8PiLgV+Caw9cjM6AKhj/NVeVYtNZSYKK5oJEhZ
3Fo0jI9CktUAGLQf/mXfANO82kTr2xuUAcJqIZrRR46KssgKkf9C7DQfk864sIl+BW1ygSstyUKB
JD8PIjm0c6HiC3Q2ilvM9mxbUVTENmt0Tkty/ER1C9eDGkRq5yjUlaDL9+hlhsPr7HGyEwdVr4Ul
bhgpS5oWmE5nCrPxegje04TnYlFDWxotGkI2B2gvMK1SZalR/CMvdBwhp+OUlL+qkQs0qzjSH9LN
N+X9PDIRsoU9ldZ1lvFl/8HvZESWN2+6nPU0HzqXR6T3iMxOmnwJxI2RYJ+BlXkvNOVP7RDmd2yy
X1fcH7ZhbVuPa6f/wPCCLovODu+p/UFWSsQwMJ3971SlYaPW/MiTxMTrW3/ZSxQH0+sXDoiyaRFd
GdAyGa5ewQHZZRijyeT0+Zlm7586E0x1IkP6KZ0jMd5jEE+Q2kkk27V4SNwugIQjBMMNOIySta9V
jZS90QHDfUoTLyAi20LPuo1tjn7qfF7kuvhtaIuTFlF9Lz/8vOLHBUpLwyDt9f3xAd2h7RJOL7zd
XFSMTZFpR3rQbGoZURKnGZx5GUT0g9bKE/JJnqCAKdS4oe+d3vDz1HWybRO61r98V9fP8ofDPvxg
6DyFIHYEffjQmKse8L8qteBx78VVqbOQ2hwTmgnngEjpfSocHoZwEV/XPYj0i/+mrOYlvBvxPAvw
cgGn3L+DCF/KWp2HS+eR6Zy3ztcCrX2Jls+wBsgAJA+A2riSk3OlzNdhKLThH1w2pD+edrt8T/mF
8PoC9OAqFDuNcY0nCdjM2QM1asstdz1Ul68H8JZGEo/rVZ/Y9B3gKgLCHLLDK+VdK22VF3DyVgJh
Chd6m8HxqCci2J/zRStohY20E4kTPOiyxG81F95sYv22Hzcr9kjU7s/rJigVodHkkDNRnipv5oV2
T87Dv57oZKFLlXejWSFfPWB6YOyklS4QCL2Q89/CY+Y9XrbMwm/Etp3YHhwUS79BNAVEmjns9uPN
/axfo68Xf0P9yvo4H04nKIyUfr6nPYNYEFFCmCdEyGqbJyBUfgksYT3V+MFb+k1WZPEfa2a237zZ
mDbCMx0WrDzC+9krpN/i9O0EGY0ih36XVBaB6NVye+Zoil+DwP6GpNqbK84I3Hllll2HQR6ni+Gq
xlBUac9RYDmOHTV6cuJvuqvfC7F3pfAYv7JlkYenO6mKMhwcsGed1bkTT5olTHNg9OraaQmiWQdQ
t3THHaP9BzcYDCQUEwmL4QpCZ7p2t/FfiszPnP0ATgF6zNPClB5fnd/Zj2U2tau/UxoYbnAkFRxI
zZmt8jGlR1sCpGIy5K67Y6SN06rBmObJlDJ0MDdKHOZNqX3HbAO7eb4ScHzF3I3s/OlmwziW9nOt
ObapqvCbZl8Tq+Iu8dvoHe4bPndiNyny/LDMC9ZSzPy+cv8/8nB2KIyqOmADVEdXqIu/tNPo3h86
0LGJPo9d4Rrq/i960SWtEMzvI0H5bKCbmAxANt7dmiUhcxzXhp+7CPNdDt8t12j+FLCBnwW3AQom
ePv4EsN85omFQLVPSLRJ0RPNWYBi5+zQxzC6DFw++V1zJbPa/NlanNG0zRY0Y5i5s3j0PeJH7oPD
zoiyPT2PxfPgEJpSf4ZyPjenlfWYDpypGyUV2FSIKqZXYWUm9aU0h13mEfh71sF99tjQrmXfjzNV
1v18UpHMgu4mO3B35OZc9XhA18HwceULyYpYQBKTfOMox0C45jfiViMMRnvGpGw5OSTFATN2pxV2
dXLTeglBm1dWXKchpH6wR2mCpA8ZMiTFt/xbnLIu0hjDWM+n9zTyof/n5/2hUYeoMEzfC/mUdR9j
af/K5YaCxFDHXGS9OKUVvblTeRxSn1mqmJAn5HMTQsYMplUt4V8fPqzb9cn3K0L5jj8jJOtmDl38
PtHz4DJWBhoSqYv6nVxgpKg2rRbw4maWFBGc52YbUfQXeU8+IuWglWPoBBCgia2/c0b/nQEYhaAJ
8IWx+QNUOWb0Q/czah116/sQPcrG1Rla69CcMVouh+PFntiWXMwciEN7yvkR68PzbNwXyhqyTsRL
T3Pp57WYqjGE44tkzcFQ2g+UL5CpIZbY7t4q1NuAH8oTLpku0Z+iiGCAXJAkPqVPo/prcWKDw0pb
aK3C6OIERwPhpJ9MOYzmvmIAOPWpkH7d+/hvMoBpnOCuLKXtVf507mnftWUqXilGV+HksrprwN0T
vdbyuXs9kz0WxG6pFs2EQzErSkkQXjv5yX4RfFlCPHywe+IwQjtbp/pE63qUa9ffg46sQY8L53iQ
YvdcVhCcZZBgNSiSza3ZEUtnYP5zg+VWMCB1CJRKpn4V9Lau3T3MzXCYNES+UQrMRm3zDJL9EBF4
KAh9PwJ7XY2XLwxHkJFk+5Hu9eMEu3GZ/m2OsNtvjB4xpgydbK66PyBF18t5A7jqI5uwoL2t4/RM
WXQFYdE0+F569otUsA5pGFS/QLw5tvY2TEO0HlwYyX/ZZxSipunnXJ+NceMyNgq1KlspzTAa4z+J
kyNWpQrYYCL8xbIgyQm0+CASN5Lv1K2pnpq3sGJgeToTNAE6ochThYIX/LiT06ZCRuJIkNBtQacK
0yhJd+eUvzWbFM5Hm7OX5eeVVnKivnv8rWsJFRSIhV338V2vqJiEJoXYa8W1xHxtL5Gpq9ZeiWDg
ShjFRA4vDa7/gZqv6RhjGYYO3G+AxsnpDD49fmKzkS21ttNXynHJww0wRF/6RrhjLGGs242wyt6C
xXkELKtBx4YdQubcYyjM6K/R0mKYNzVt2WQj1i4o/pMKKLCxf/vQce4Y2P3+zm60L+tHqc0hhLL+
d9PAftcuBWRmfIxyKgQwbI8SA8kauEG9ow5rcEOzRO8uMDgHdw6nIIV8asa7dPOp0At95nMfm03m
UoQx7F/1cY0XHA7v9iMN6c+yUMyFUHWD5+ANioO1zoiki1VS0iEP9By8ZjV3jzyd34GxBLdYX7D3
eLWOn48VvCwz56ikI/0oWsTzoAZnqlYg8PmwvzpngR+gU5DpM5SowPMPJHp3vfy2n/p355GKpXsJ
H3KFNuY+FDnweqmoyF4b4Cy+ltC4dndbg9yIekhkhoEO/Fh5F4OV5XfZappH3j5AeSexKLm4hA0l
yxvi7acu6xMSbLDsPHwwh8arxWjh8PpTcw9xleSPABDcnYsjLMGovTtv+pwAEQwRgAX/YexdDwVd
J/l3IuvOOv82jGr+HPC80ty6R6y40PXptGK/0GqZRRedE547mArUga7JOS6jAVgRrR6NghixrogA
/j7hoUP0iTOX2mbYh5zKAaMwOqXyaTQoWNwsYfe7Ivh5rV0W1ubzgcgyCUDHy+pabHVMVNZCTq8n
SLcCvL69be2hpeMtBwUzsEyuJd3Y+WwNSiQz0a0GuK/AZfJIkq0gG3WsSNZlpA+/XLnyIWBteE2P
m1HkwOaHClEMlKbwcNU2gwJVr6j1yLxGApDFTSWzy+uadksrVg6OiaF5r74N2wneyrWBdoNo89bU
mL77/HqyS+eS/uef/qthjWJPfQGU03M9WaS5T9irTCr4mvLFMm/mYuovlSeeXFbCYtIyUXc8GeD7
BVYXgijdJLXo3fzAK43kzI6VIluBf66R0aYU0t5mc9zGEOan4CiB+GXPELSuQvluNDYI4bZbcyKJ
KxpkeV872P8zUxDB+wBan8d4ZIvHyKi2hTP7ZOBvdVSLtKTbz8L4w/J1VKL3JunGtxXvhkP0upRQ
sKpGBwB27ZHKU5iwTdsvXvqfYKGDIyDK/ELiUwCm+F5ndo4jQZVGAzjAS+aXOr1Biy6PulZ+uxWq
FEJbMHyzz7q8DW5lWlD9TZaSZa1aArXhF/l/17H7RTp/2Tkav37l/gKoz0GjYupSNa2qAp9gFJ/I
JqvHvRyDiPc9ksjwwEF3tCoyqe9hvh5mrgloBzMUUUV7qFViNjO9SpTCcCqSKBeVgV3o/IGiVG6D
itYP4GMJc/ITu9HLIaiQtmlcmmCvQWZetg5YqcvsZiCTy+1zgE6M2pUezGYDy62PQ29AX2Wut+dQ
eJ+UreZF5bkM+8zkOTVHEIu/lgnUkU4eLnMuJHmY+6wTt3EDmaJHfr53e4QYfUEkzYnowb+NP83N
3P/S0xjXKY/9iP4f+e8/1ULYCzcyfPHtrIStjeZq2+Ol6HRvNTvVaXMQjxOGkAJigBdB/ovuWW0e
IWj7Qp52u8Mx+EZF+1xvPhpC2OIbS5e/mxHibqlzMBl3EAGtU01HDXDzi2109mZ0CmsnOCkx0Fpl
PT02jZYl3c4OjlcTr/UXpPlqBjhh6/nd1z9FtjmREfYfjmZn/LPgUlWbU2Rd40mrt+2v1z1q7FQu
6PFWKQG3Y2i1p1RK3PhL4h4l6gZLwMV0KWE4Rs9TAetRoYpUvk194NSGXNt8VxPn1u0Hmo12BjJo
d/9FW8e9GFImiYV6kis5JWX0rD8HNrgxxTDTkPCffA5j2SQy+PS3QdcDX9NNKOfRZDRIqJvgQqOL
U37g6T/5P1Cbdjx9+cYvCGjWm4W3xeP1ZpU9VSfDhbJG2jfflGI7NwbGRvK8SHMzW9U/bKrRFLDo
XJKrsH88RBONTzSTK1s3b2GCsKy3nDnvgQITnxp7UW+bTfiOffYjqfY+gUgk560HEwgqychRk+LI
Mr3aaBHj5SN2PQjs9k44APLRlaXvkVQfmuZABATsnR9OiCtHxk+5tFigF4rgyvkcLOrFSSBoECSo
4aOtn/pVRzFVhzU7XFcVS7m0Z/O6YLRvC7AaDCcx900vx79/Fb72nuDxjhqbPmLjZqWrFK/9r4Ts
Ac1ZhMPDhAYr5bCnAMwaFu87UpdH4MXZmP6brTWgFoIyGQoKYq1CpDnEAiqNoAAW5u54bkh+5ZYC
o1W2B+CXB8tjbxo55Rq7wI7OV3H4IzoosmTkrQ2U+E/eUw2lsDKh7hRN70ZISySV/RcEu2+XgCVY
DoH8dwwWgCsHl2qESZfW8JkGfGDrLexbHWdRCX8IdSqYc63I4ZUxY3/D82NBraPUe33PYIGqEPJ0
/au43szppKPzipupInixweYklrCE6Ckwu4QBM+SD3RBH9S/oivFR/YyPI5senRVOD1ZW+Kz7T+HQ
ZwvEjpos7qGYMAPxSY4BzbPUJZ2xToCljdwftYBY+9GB2hwVo29Rx+RQOEA+2ftClKBokt/zzIe2
a72RaJQarS4H1W3d2j6utWcyXJ02SqOQ6vCD4TFDKJtpkb4AfmQsdmIESKkMbrca9sig/IMjTVG1
ZnDr2djS1RQeya7Iv8xIEbZk8Qo5r8B/Oew2vk7Gt2ibjMHRiw2EfORiQ5BBuc3T1Q7Njxzp3KXl
NNXe48fjN7x+UFkP72XNtZh7VludMQg7hJTdAOiJ/I8AbgUoYbTMpa22PZFN2D4A0H3p8G2+6sCl
TGykD/DtzpFdeJEMmSbkasUIk72Hy6qvmr772YW5yUjtzjr3ArwzdQEFDVSn+J+9lKQq1EclHZbX
ftLnhmqBTJE6aIHWx3vRwryJ1R0vnew+BhMIH5gey0ylzaNkU42DmxI9wdQVWyOOBUhkB9njnROA
3ooWMpXWclQhsrv4Qr89sF/3eykSpbaAKeD4tQeBqmrG2v96LCoNUcqbPX25ULnfmkzp+eA93KZB
Acg3N5Jo2uNBtPtzqPvUJ4IFzqtXwcrrUBOuFL5g4DejjQzRNcwhQayp1npeZ4DPxo0UvPemEz9h
CsjKBVnDyt9UkpFtYGIirn8YgJTfeUABbOdjuJv/muIg4EkKo2lRmxZBMdCfzOPTA3hQQ5T4yed5
falX6I+VR5CQ5dWcbeMYAGzitEr3A3ABbGjz+cl4GKAyJY76DDR0YDzkqZE1HTe8Yb+su65rH8KY
nUIKtdkX5fbk0aNXSzRGb0QtL8UfbI0bDlLB5t6KYRPXRTsYHGIYlvDqAmVCunIY9CHEZIJpfwl1
mBB048Euie8o6YrgxNrttjlB+paCVUARi5Fj7CD1nFiFvqIhhzj8KkGkPSYxy630YMkU4nxJtny1
8iCLn3rnIxovJD7MfMVYeFGNOW5FP44Qm3pR6zbo6VB+IZiH4o+57zEP1zgD9mUSuC7xeYQct31T
IIepxs2bVCdhrN6OLDmJj6KXSfadS7B/HMX6hI9XGXELwWtS5fJAva2k4dzQbbu4YbjSNU8fFmJ6
/b3IzwG8xT5L29ZfJ1Ds4+dGhw0QPy0W6cErm3T3DUBaWT/EkjgsCAMwUrKBdcuC1iYGWlDJDzQ1
T5S1+PkounFX3Br2JLKJ+vX4RtBtoUe7kIzHrA6K3UBgcvpsZbTki0nm2z+PkOFso73lZzmKG1RW
7cj3nyRiaxxie/OxeItdvqDSi/+gRUKjWyqo/KaoMTw6GV5u1lbLODYxWErnRdPg3+X2fRSE5Wpd
Gl06+1oCbc2h3dDQ1Dl2bqsil0HQYwciUZgqhqL9pWcJxYoFFjWLZOCy3LUBHajxisTGkZ0zB+PV
8WSN5xgtf95EfPv9gfBvaPVXVGDvfdodITUkDBNpsI0zx0UjhuEq9h/NNQbrUtcRbC3pK2IgPuI5
BbNheTyvJBiPJRIiIwD2wtmMu3weSLjqdke6ZyNxFKGVAE7+nTIokTPjzUcexU7SXkaUv3bDDGDk
fbZm1T5vgHPcFlGku6jjwo6QKHGgwU0jQo5rSd13/LPl4w0TrgEr2MC6UDweYtVPRieyg7itfxFi
7oYSfdBOl7zkiHv/ijANWbHKk7Hi1XslKqTgKWMpAhNLJhKkgqB5Vu5fzohw3sUPj1upyXoGM6c/
mdKI1ee2n08FtvARaEstF1e/HhH+PiuGciJPjzdVSV4Vqg5HkfhU7KHiEjgEOvWevs0TjsrzJlVw
djau3n0fWzN+6Nuu3ijMOdVSNKiLwEUms9L+GG/My7cdvh1LozyE+L/enFSQ0d7D3XScbC8Vafq8
uFsnE991OenP79d1wYJQI04g9oMDAp73M9909LpOgbZMl750HWJKIiOFdOqpMojASYyf9IZZLxrk
T2T6pl2oCY7hEM7mqB1V2DMgWIyvx5JYNze/sQJVQi/cgNQnwi/ymNPL51gRhio/GlNoLoKt6m52
bq3gzp6w0I4LpQNnb49BwmvKTdyyQ/e1bDvq25ThA9enSy1YbLLjTMuUQ+2sA49nn6tx4uox6uKm
TlzjnTQeX9CS94GdcHN9MpgQMRYYj+IiHhS30KwYxJxa3aEmC0xMaE9SG9zfbk0uDwnQ6YJW6Eqb
QcZ4KAMErFOWA8K8wTTi3RoXqHenIPxZ0JSLdTs9Wy3z2wWI6a4nuhCC4nED19glGeJnVMDH7do8
0UB/6dCkrDTjGkz96imUrbJ6BpvzSfwfHRWEUou6Yp+XAFoxjlYSeN2c6+yq1v22bViJx4oPZMYu
NskfNOR9kiVHpP2PgC83Uo36zDRS09ydyRqbT2jKnwPkNfChFPEeCQV6DUNRmrIPf/i6s4Mi0LJh
qaqR5LUtzq+OotVycK3qgFKqUCeQD4ydBJjWm5cNgE3lU/2oVVHgIqOtoyxop25MzsOnkkltai8r
h+eN3jSB3LkVuAvKNER49OfaaEH+TnE2viZxxJ5Rbhf/1VfsCdCsaauTQRoZ1iUmWlPYnt0XlAyt
VNvXyeIvUTApYVGSM62IqaomPtVd+odVFYmlS2E7EtTZPSVWbTxdGXLOE8YVZOye9I0zUUn8tDAl
r7uGvN+Wp/REjnrMNLnAP0C3/KIawMFN5L1c1nnRaICh2AoXo4FZbHyFrXWOQP+giDrO7Fk8q0vW
ZqENttE1+pgUPpaWEndcRd2YF87mBihCtCziUkukt9YyZpnxKhHWBlKa0vyNPs/zQYg/JX5rUoRh
4Z5t0/YYjZK4kvEAPBqVExPXr80p31Qp8RDTG4FyKWy3FdiAjhNMDZToHAjAXfH14+oibIGcK3kO
053QIUhB2jT/rDiTvEjvC1wW347yoXOEEbnGTUTbdv+ThCyO5c1dzfsxaGxOgr8EQwmYByVWAb8/
3ibKwNJtL5dIIMBi8YXSIiVfeoNvVCuaGpNh/mQjyYxTaqIlqHR5DLMVwy4p1aG8YIoxq2CyWUgg
h0biMUTTj9meCQsEYDIAXx1az+6ewOc3ODUJpTGxI2LWxxtdSNKThXSuz4D0pdt4iSSdfpqG/YO2
rU+HT4GgcBKvmAeVJ7Xcty8/vH+yHk5cHVlDPJqeicoddmEw7oJE5cBlpkQ9+3orBSzSJLVKMFvb
DzD617gjnQN+x22aOMRcrhjJkwwufVAVOu4dMq2IJTWEH0co7klb4yOxjsfLRsOxUGZ41grj+AM/
llFHQsPBmmuhZTG5Z2BzZ/CUgytL4dyeaC1loEQJMhrzaqNvfQYUGrHmNbB6Mwdv7mjfAbIp9t/E
kuGdWmLIWDo4iV41ar5lepddIWUod8QHpXwHxWMmL9JwfPf5dxRKi+DviXRXL6AhfFLOHIjR/2Zb
cYyhtGYPj9ssDV3eEUYuYc6FG2ely7IZdYApBRc0CW2U1i3GDUwAqCLPFZhySdbTAW3DksjDtesx
blr2IA6V583hjPaxbj8jy0NkH25dE8wZbtZTU/BjoCdWnrKEd+4tEzy60AnWBpTe9TSc72ONkQXE
KtaXdT5H3G83n23etcfjNrytKHAe4O25EEuOLym0PJxVNbXyY2hX8OV0PjB79jCIcUZzRbHw5Os/
wpAtN34yTy0dDKD6pz6S8Fhmc5+XBQaFwiHms0HjuLIKpGLDdsVRC3I5rehSEmLA4KnL0tVd0aVx
3+fmd97YrhTu99EFqzoQfilYnCD4Ne+3TQSZswD1rGycQw1OkI1mM+1INfRKFroW3HG4OHdXwMFb
Hxi81VMa0qwmNUt3KaUPsbFPk1EHtdO+Rm+J2FUzrIgKmTuHpg46qxuecz+/cBzbj+jjhKenfFio
N2KxGgmxg+Q4d4IBzq0AtS0ltjIO5D38oS8Mmd8K8imaOpIOLtSr+nGmHhK3RPRVYW+HTFyY/2o9
fnUxZF5Elh5k+lSfY4GOGBX68vtZyWq4JahSF/pPiTJaXdD/eVY2nVzFXZ3VkMB5akD+1WMKaY6u
TRZzrt7HSQmJ1lf+YZLQlH6Unrgqug7p5Rp5KgwLNHLj1ErBNEIFUHVT3MH8UUtZ/cvbb+Lbih3J
g0/kP7wpTbfpbzpBF0oQLRZJHvDom4QaA4qvbmmITMzxxsK/M+LHUcxx9mNfVVE7pOC//kHuMqBq
N3QAJ7zSn5btfJ0mvzMVWE6GpmKGBpG7GiqmOOawvTq1cfFItz2C+1U5DJuFWE6U9Im6hWoCwOf4
6LeW1JPGhder9avaYKDUrV4UMS7/sUCkD4GBzczrCq0lb4JqR4jLIza/soffPiO9yDfaWaklqqfI
aIv1nc2jdczuUVgXtu8uIbPmTsRR5cL03ko8nhk+DKxs8MdPegeK2wZyi9tc4ZGthtjsvueHSXps
CEJMAPxcRjypAbiogjCfdTye9OogAQvrvSkWCLpPn6NfKje86UjM/SXA12JKzDqfavwJNLI8JEAZ
LvTcEEqnM0fd/w2UyPQkudvfHgRpOw/8FfZK2pWeAGrBHlnBKAfim2lXjQg1Re9EyYNK9m/U4Mxj
5CiKJOmDfKPat2yN+wvJNp/dTDY4ox5R6BPmIit6zOamc2p9d2h12B6qDsCu/JFqsN8hkmmfYEUE
s0g/B5esKUifnxKt8XJmOMsbmfuxmkEQc862NDzH+HvzpAATmjgMMleI8RcavazE7M5cB5RWXvBN
vLuB1oUPDIO/S6caKziZ3f7wG33VxU5u4XJXT9/QOg6bBErWMCQ6dcs0bhDyRuyaCJdNTFvkssiQ
r/JPUHh9rDeRzTP/5JDYRjFBMVDeaK5LVWBkmzgFcVRug9ojF2yvaOXwWjudZA5Vd06Y8yRjya8P
xDYVm3SCYEFohrGvtaYtMMSIiK1aVWtmfPG77pq9RjkaKABL4uAlhLHgHCRN+ZUocCE5ugwvCfLi
oYuKIDzUbGxPLNwLBD135Oh9wH+kd3sfnmVEId6TG5fsI5XlYd13dN4EaRAtIt1gBgvMGlcdPqXD
SMIE2L23ArlE2Aeo1yvbYFfkBlUT7xZhhAs+nBT+wH9AWeFE/v37ccrE51YjReVZ7+f1dic+wVkY
lpDmOJ68VwRHhsHprFX5xj3bwBkb1OdqYibVGPFxFXw8BwZZqmrSI5DScWC3qF60LLVPt/SMutJS
i42wafDL8aJlbcQ5MuVTwf8XuX1fIHVgrbYMe8dqGW1Yhpk9dTRnyn/LXGC/hfu7COD9OO2NA6cI
50wqmERSBakuGn5vOBMPjlWFPYe44b20rtNdEBeawIJxyuA1b9zIaqq72LuhUe3s2NEybYEJjwQU
Zowal4YAbarvdJwyHFcy05+WLF5tsAX3SvugcFVHnpFDee24BGivx7ZHAzb9lOvIiKw7MkadcqV5
990wEglWftKtfritzyETKoogVnvDtwY2CUEOaVPKbdxr0zwRM2a+D/3BRFBQtRqib+DMwmh4iX8c
WmCDRswe6pAaiIZezfPFj1xmlCL/DmRaRes9YxHPSjPedXxz21RU/6Xn8fMjWYf8wg83w1XjHagu
CRca9lC89DmsjBZbIycyD0qyJ0peVLiOR6uagOOVL6Clkx6L4O5gdg1cQK+oMSJmJt/+bQxH+VHD
TaOf07mCl/vT6dnecOI8+yPMeb741f8iC5lvAJuSTzA7o9A77VbIOD3WxbrCMyyTxlAWD9MyUtxW
WVLDQjAVmPO+HibyPRYUTA673pWgplQU1T+L7cywTDF3X/8P6gYc9D2HkvQTwgZl8iW0I6euLA0u
aBY+FFL8Z2GAlPbjhTNkkRwTJpGn1AMjftTEHA9gretJ1+0iubpA5zUfw4CHJdqvZihhCgfDUxbI
wq1pYLyrydYXfzQRMQg0QTS+eGn2eG5+a243+RLEXRZX8wUR+RSlNodbJQz5GeevCPe1YupLgmib
f9xoFpgXUj6TrcZLjlZjVNTW5QQ6zNOlM16HU/y/Rp5AQo4tIuPqcF2eJmJb7qcMwkk+23HIN6Gx
Tllq94dNHM+yC32+kr5sdW/Aht6bl4n4nkuPT0y4TuxOG7PgCEGES/NFJzszSSruwRJik9NArLCF
p0MPY/+9EojbxyANqJzUlg61/6MErsp/Ac6tG6HlUlecnsA+3LibAqm+mXLxyy4gLIUhSip2jeft
RTHUDsnKFU1ebUzmZzTWSnpBSByEZ5Fz7Sc3ew55SEjYP8Cgu4l4p7pSqm9gB00YsFqcJx5R/kVr
RNXYdfcR3OHjoUGy9e76kiys34nlpeHVwUk3TY8ovPkFuPxwutSEjNSg0HtQELG+aaqdeaVJtIew
t6b7Ei0Oamkv6nmML9jHBB6TQDzXUJZPqSO2vtYUJdPCEoEODKcSFnFV14Wfa5w75vsGNHMXaHQY
uoCmrlEirEfzE2qYtvCX0eEZ9phkTXcHmrRXEViACkczKZ9LbdQWdV4CZY08iYDWC/h+Ys3UJdTA
dk7Eh3seJdgrzqL06/JKSEVjL2n6GKuGQVxxmmatlawBooCPGDzTAFs8ns86kswo1Xn3p8dMM2EJ
QdbUdBEUTtUSStfFUEz+iz7KobmCC68VAJFKntuLIqGCJunb1e73ItuIYbCRixQJ97fDkbL324x6
PReu+87r5BAV7/ueeKPtbXtN3mfMZnEx1NoTTp4Cxce/gDWAagk8PmyAMJLl8rA7D6+s3W8wEjhW
H8iBcSK+UKdiikk4IdbsMZqmeAoTFt7fBXW0b0VITO0tGDNIU3OsBalY3czz0vJ0HKoQ3t5PGJgz
XI5t60/MKyrG1XaIvY8VM2FFgcvyaZDmlz5KNHlfww3FTSuVoKcPuIeo/spRVVP5SQM3i0SsXdgy
mij/khk01fmt2pzKgBINKyYjr4SBUJCkvh+cJE4wDtnZYNWBE6BVLxQlALdEUoWsc6S0f+Drw4rR
ZdaZoK94z2JUQrWkWR1XdE3xebhgcD/85QoYbegqfYHfgVupYG5LNGidPeSN2V9j7HLz8mibUcG2
jIGWaki+W096gz9M9ZpJtSKY7r2F4JJUa5ERcWZajq3ulZnlSXaDRqD5g0mBw5BQaG/eUgLNRXsU
5xTbcW4AmPnPIohUzMwkoOYUyhLsJMG339GcrlyR938C1PulqcKGJRSIS9ZLJc5DRvu+h0dMcSnQ
kOKintkZ4/jdjEwrSiHUCHGu7CRqZuNbyks7ih++wFNwn8olpKs+Fcvyrv1E22wr8E/P9G6QXnuf
4JO7LM0rn0B60GancJ4f6EtwrSaWrnrpZ39MOeIJ9hBmB/oQboCf/XX3VhjtShqEXmHxqDVSFr30
mpbHLEHmPu+bxsDKDmjTSRqdgNdbTU02/12osF8SbqtcvVJUdNDku9EM5gog71XBR6mnxoElST2P
gaY9YwKcLA+5volpmH2awG28GTM1NBgf1IEZGksHXPGuAgJIrUYrnb26qem3Y9UM4DgKMoad/TkE
/w/QIgcsFxyZVPPGglHpYEReUTQG2pwdI0XFm+34DnXwxd/f7jY0xq/1ubuVQkDPEzD7AyQmDPmw
GOvdP3SP6txCMJ6voUuHuLKprcNFCj5mRA5Y5bV7lTjfvAUkhGsg0Supg6INiPs0OSbNnnFR6VOX
l6cKUZNz+Cg/sTHWq1OfoNIG31Gqwp3iQcDuSkbR0uAfLNPvjgV3ddUiY41w5cJe6bln/rpkT6fO
9Sx0yYOCEYGPyn376nIaYnRP8h00Pk7ImPl75hGjlTKvADlK4b/QyBaFiqzB+nJfAY645v9QFLv7
mz9ryajxMGors8HCPtfeNl9gHLBhjapxeI6PeIHYgSzBacDkeuwfuco7EJalisIedoAWTf6EHLqe
NkijkTAyDo/0nsgKGaVENRXQLhGN/3dR2h7hFbMO1y5NL9LE67HqQN9Vwf7AiLKxi7K+2thmEVaL
b58WchNqnzCYaP3Lk2dTJvAsO0g2LpRmIdjIp3VlNBzjZ1/WU0YFxX0P9XFgbab6ugVk7wFYYCKf
wkbkSBkfILuKjLzouTAexCE8fNClYMjFc5rAMdczGfMopIUrA4Wayl2nYSbKS/q82svnj2rddxVS
smPeQUGpK7NObi+vYevHBJPpN5NSjIfvHU0cvBsm8gpb94BaTe6pKl7VY6/tu55g/KOO80Zl5Pbz
P1HndUIAWehjPKWMQVG/CB/oCDeMUlXQ+In6IhNeeJ+5G171OG08AIWejnGE/cTyjKVLK8M+/n/+
Rp5Z/mwmPTOUDaBBUULY2LyMs0UEkcc8+PyDZ4fAFdTSUCxtAVVle7IMj10zFIQbv0BSS69eB6bE
1u786ypuEVIDDJj3U6rjukzEJ5lPF2vaPbF2XbL0c/zH6qTxA2tK4lDIe377TLle294CKnSy/Znp
8g/Q3AdjBaEbeQQrQUGlCxX4Rc5jDueU2KvkUAgLqmcQvWaSzX7KsKFe2j6wKoNQCOpdapOzjptI
CxlS6TTuuPptiM8kEV4zvUMGsMoNoWNMd5iJi+Ls1kSYHyO1EihVwtwtNIv0wcWbi6bXEm8BCbs4
9rjPxNYExP0XV6bI6PRVaZHZQ6eWamv4n6xx87xtOQ3qLBLubnEgCat+r/mfAsdRrFJ7smWpFno/
59MDPNBYGx86Pcarf1BkGaUO4fXu/wlu/9AY1vwrEwyWpkqt19LcfC9ZnDkCTZtjpnSJG/j4oYPV
LB525mGiu/MIiWwwjW9+oYQ1wM3VhvQpRphVl3Jp2vYbUqn0m8jngeYWlCPlEgwj5mn+ab36U3qK
+Klk1CxoEwRyHMQOpOQYIrlak/oOFTHq0Af7E6qQOTuvhArqQwduvdeH4hPNXX5JNhAw8WzBo7A2
UfGFXtOHMz3cjhVU7GEGvvJgwLW6Q/uMI+jVc43zB6L2CE2jBsB1kElEp4EU4yeDtApI9qN8jNfH
SJrmImoSXUoKJaDWa/f+dNHQbpeSfBd9oASrc7u3+7P6JFsh6Igz9XYNqPpA+JX5VNG3jjsqwvzh
UQ3MFUF6o4Q7jteLfQbCr+iEKcN0IlNvfFaSbqyAFpweDQ88WkhFL3fb9dAmQQpqCfspZKGzJh5l
cRv6rXJ+YDiJItpJkSe/lltJJ210/j0IOt4aA/Mq2T1Qy4Efkvxx9SX67LBq4ca/3TT1OTHA298P
6z3Hd2ZsMullQ93t4e/Pxqb9AgsX5nopGhSz/h9wwLqHwJTYam9mrfEqouELoMGYcvBRLJ3Tboyg
f+mGhPzzUYKE1IA4x+329iXOqZ9PrBhEBSxaIMLMrHQJ8mNX698gPrM/tItLcHI2y3dwOp+mT7N9
zW1hlhMYAQ2sDEELymEdfyAOASk6iQfi5zv34JDNwaoJ5npKVhg+T+nw4JRCnt/KuYEibYDKRWgl
75WW49vy/QfH5pQb6ljQ5Q263mtZLuvcMDkpr0IzyqNXQJAdRMgMdDN2V4PRE6IMXYjSdGY0EWXE
Nd0gaQjLPYiRIuwkqcAlzByyKT58STu8PlYu2yk4WnBOtdCzWkxmcRM4LLb/OcmUD6O3KLlqY/py
sLdaIhNGu4R/SKBRKRAWg0N6W7BVBNPbIOlxP/NlSG99p09fZs4NA72fO+0g64L99eo7ihpldfSt
XjsNsYaQB6VzRq631+S+5LsQiFn10gi/mPLgISmNtsHbQn3A1js1vzdlPyOUL/lB1ahOSrcR7CtR
y6VWmEHPN7d3Olkg3q6JjyYaG7Ka2f0tdNrKMufHZjXDL+2n25ITEPevCy4jpxOgmN2WxZ03NJqo
awR0X/CaOQWN2L7CuQFbKQfOm2Lob0UI9K0FqlPqTDvIcw9yvY6Kcx+0YcdkDAMWPYhuR8yYPCnk
NfOSSIZWAR8BQ3ofTdg0PpPHoaEwUJhJcSNfEpTrZGtGZpjpFyj6lOBNRNKeI7Yls2hb6cX+u0Nt
hpXkNkDxMXxrqn1Y0nGQgYzeRQjOWFU29CzmQlM87tsDElqxJTbDMEKPWx/UG1iROqh+3Azoqw3P
3mmZBED/bz/IqC8FcFyb+ec/Mug5kbnQeoAK/jO6VAEw9T+Q8NYSFg1WshDe/dlIxtUxWZQ4EcDo
canMB1JTDRn/VtjJW4ZIJ7aYYaxwEiN0YYT7fIcdPGizuwHEAyMapv54jFp5r1qZlkDMuvP5BjHf
J5vGjwJBrU/bdSG5l7j1Q1N3XRL5AGkaK5cv50Q2odXadRkQCgRuXFj8nrIn5qpodlcRnNPIwgZT
dm1gpodhZKROejR6YGzOmt44YVPXqAWJpW4tVupPnXo5BaE95PAXfeswFtcBxVmckyWUHa/u8BPr
rzueETsrwAmfqqG2iBwzISdY9zP+5TARpbThvoe6obntlofGL5clBalDKez4PLzeHZjPtSF1nVGv
N9MeAYATn9NtBAIdqnSBndGVRMmEMKPMeU8d0voFmYVFj8tZJ7dgog2FGWr1Dk9ENW5DD//uUU8y
cRdJnD7bT/RxGCjrhG/rMqhYQsO4TH1Cn0EPy+C3dXTnrcxgXnKM72+2vFlIaXlByvZYQG0RDoWP
HYwerKrO+JQzhCMj7EOzL1exDItm4wijifWRl7cElM8G5hPbeKg752xlO/FpitJwonvpTyUGvSq7
k//eL05rTQQyu5+kqD0pB+eYbPNz/jF935iqS8WpA3V1TmfqiTMElSIROMr7uI109wChY6GEafsI
uuqho9eCw4ylEoNfdN/xvypaVt4Hp9L/v4MdeE8Q7zl6uqV233sXGfdsf7eItitRazf9p+iVWWj8
jWye/Vqg+cFZntb0kSs+05jZ7X63P2pr5+NDmD/dp71mgBHnUPcOSODV6vtwYtj5f52jgqu569rA
EcyRsNRfDHLgU90kizIrr2w89JMS8wAdvTYvHTUdvxgrfokRcH4CjloSsdMTiP20GEmbtE7JTbs0
3iPuK9yb5cBM8mLmcHJde/XWIME5FwDD8CBFcGN1rNUfq4efYkKnQ170IuGiRDiWjcWJwBLh/RXE
K0EOSIeLvL3E88Z95AuT64O/DnN9X+LiOWTTOcLblTvepzbSpMQQoUKmL/+wAZn/PUNqSO8QhG1t
cUUVM6KEGC0vU8A30i0iNEkRIGgZIdgVsrCdYpvWlEnzzXsMqsAplApu4n3ruzpnYgLZsEfSuEx/
ypFdjnTaqu75/kphAExBAe8w4wBF7HOdRtyvDLcBeQoYGN1x7pbNbO+wC7PXm8Pc/EHrvdpufr4F
9f2L1IOvfR73XLDL01SMZffv2ixDVTD5zmZ1dfQ1FwVx3qt6IaJKAgeeNSvleGSFKNemJs4egxFm
Ld4v+h3RIiRbonfbGlc4p1qDNctWWhTmjdb+CORMZuBa7LCOPs9WraxnbpAHAq1Eb3/eN3XLJbBQ
2DNsNx4XY1z2aPUWoB31F2t8Fjn4QP8StFtst2Kl0VhQupAUah7ViEneCy+V3AqrqvsXJreb+2Xq
Bc6hfPVftSu83a3j1AJcTfg0KSEa2bvGSTIVSSoeJcXpPeYtIUpt/fUYnoVK/Mv/cskGkviocGDO
4SIJesZgnCfA3bCto2SJbnYrCrbSgsFaevzZL28fxr6Zfj5LJgH8syZBmeQD+4bWnno2Beh29x3P
ZGR2oYbJcG5wKk5dQIDYKyGgPGiqU23yXU5KjEnPxkKkfA4/SurcHKftXTytsbZf5MJVcJ4zjL+L
oDsYyu+RVe510s0+FHCjSTb5dBMW8++idNp1G4hpRdGRCqe+MHJKnk8m2PVYoYJlnhbNHFs7EiGr
x057nS9xMSkkyHWAgHKBIV0brUyQjbrHFjFamRa4JkSlqHWrfBubw+wkFiVmOWxau8n2pRZQ1QbI
dH8Co3IDfYehSxsCDmvq1NCnSXCj2UqCT/O/ljT2e9fG49lfFhhpcmLEOPFeWpSWfCej6Bo0LUZS
RziCuqPlMbK2Zn7eiN/1cRYJEHM5mGRGMouNLq5btgu/yB2Uk86QqI6irwtnKvAVQQvYemVhPv2j
Y5uLPNOmpZXxRWq/skygPBjTofDC8XNThPmS7PQVcfOTrN6te8vIcnyEOPAAq7OK29ILfe69UArd
iYklmFcLsoKXopwoq4rugOPllTppzXwJBVFKQBq5t1IXjaZKRRfeeXv9nAAu84AnKbHjL5SgLdB3
uh1dYqN5ethFtH5SztRr/OwfPPS6nSi/EieynmJuYkwONm8JsHLOmS+qeoO28g5FzsLT3K2zXQrP
R52opwRfSzgKlIrPbqS5ichm7b0dUo4u3mOR6/MhymsLvY/X9G/OZljbNkvMUXaGS1bLxkp5XgjX
fJ+o3E1ZreYNr/L/gcgHkazc/Xtx9kZH28tTGSuwvmOw8VGBWYJ4bOb88YftFRS+BgT7DNSYGiS9
5giLnlOulc5wwvpfrrJ2PNiqf/ItIRDscGLBpKnKE8mqvBO7XyU+oVNBtOu2PLWsFglR2JPOuCtJ
8VKwpB1QZyvvUnU2eOLZBadIpfJGGoFsGpBqebvST8O7UyK6WgPHu/zduJPHw0kz4BlEbj25/CiE
/CuZSu6jDx0OmdqYaGWfo0omjyeSllaYsvlhmLOTAhdkr8iapsjpPSAU88qb5wlQ8JwfV9ui45LP
CI0hZVAYGEKBPPJbc/o58YmsvxEh1VQ8JVUdGkvFMNnj85TBfnx9gAX9vZtLmkblu+sJh651hSIH
oqlrGWLRF2kSC/c4FyzxV9THx2u+g78r72ywvU8uUpzK9hR6S+yrBeLBBnk3TAUpXYU8TII0kbes
wn0Ek/A5cCx0yXQhARlYKgbbHexbeiEtH2hIiGDLTtbvMzKz51kroLLlWTiWPGd3nuMpjojUw5xw
LRdjiXf1TYqwiUmT/Hs4QGBdH0xhMowRkw6OYj8ce5uRw3n8U5qPPfSQI6PB5SfK78Hfi/8Pup5B
3HxgH1loKMMkvtEKuwdM4vIFq26hmyBefkr3ghxdI1J+CkR29YZ2fFppGa0S0MC8DrnIrAxrojfb
gyC90NNpvPf0+7QaTlT3et2qtc+0cVkYAQIMqw8NVPfzYxg0DPnW+2ejrIWkOt/yxYi+tz4foCfV
90h4PheEeo5yOIUCgOiNjl8rG7tUWpp6EZdewpiO5hL1op8+Pg/mURiBo5oi/kjfT/K35SEmnaiy
ACiTwdq7LGaZf9BT8W/wBY7PvWKgm0rc5lPoxXpO0gDaKvlvjj46e4QO21jShPy/DIxEISDiZ4aG
RzrAz8yApJoeTnxJMpHGtx9ia+wz7LnJMhoC8fa9zli009u2pb/Vpf7k3tKBBIFmadYLUUqhsZXH
1+fn0fggwft6KLhTFRPtAbMrAK4RA8atStoGY7gbAeBo7E82fmmyCFJCMi0gf0kKoClXl2NVpPJj
pREKLSs6efAwc5z2hIdhB22BQ3xjDa/myQvGxeX3mFPNq4eY0/3So6/SYHOP1BFgYZZUdMYIDi1n
+GRhpH3hY4LuQJajCkK5Ppahmu28075IhpxZJzTCOyEEKbLyeDf6MTi/qv1BCCKO659OcBlFqC+K
aCoRNqEvFeNELrDSvkuWjrjcqZc0dySsc3JifiMt/6w3VEFrWoKyLPTlCakC06LjsBF5l68LJfK6
/d/Jhz+nErIk+lywSEZNnou8NPcIbxbbPSl1alY06/hg9EjSDy9GbJpPFK3wKccv/NDh1PsPzIoM
h7FO7+QmztMs0Hge52hj5XlzqB41MRuA3m1E6OKdNrTaEAj7sFDuOAYB37anm09s8k0ON8Ktl7cj
0YUpdBprMudyFhGKmmfiVW+Z7Da23fcBTaI36XaUqscZq7PlEbfjpz8KE5ZE+d8NPtoDQu3pUu4p
WbIYT8oK2QKUFsm/9x1wzL8/c9rAgd/Rjayk81PIaU+CgQOZ7FMdJRPz0uNyfxXlcUzvdDovqLiH
HHzqmq15Z9dJQ5fLGoPZBbatJoicOeQHjlY85LgRMdiykSv6CHxhHDiL/+wKZ03p2Gkjiw90gbBI
nFExmFukT/DaNZ88aaJyXj7I7u0EF0zXv5gnxrN3LWGPKefqrzdPdB/pzJ6IkQBtsP0o67d05//R
E47WaUVD0+jiTgEws4eHQStwSF7WYH8n1KItgPvJQfh2cLdPWpjMH/OannDEMQigCPiIs2eB/xeo
Uy/6WnZ4naBwn13nO9W95+17lW95eUxOEtwDFrrJbbUrvHL7m/C+qWDbbb1AR5SMB9YbtqJ9NbjH
OyQ+6mcD11GopFrEy+kCLZEJYm4TEalUU/PKhZ8423A2sHd75W5+J66eWgt6DNuL71ar5DM0+RDU
yPSmMxgao4OQ9hujBLY3dr2mo6dWIkrjnJs87U6NdjXl/y3TwK6J1QCE8ry50C9AAPukLaB7/pub
F9DkXYJdioDNK+0lORVRdwj7I4xomHDAAWfWumHzGnIkIcluQJC2pA9zExBQ3KHMEqze4YTLlBnx
VsdRB1SMcCDAhntfObYnV1amfW1zcJiKXoj1uk6+c4APRKR6m4+tweTtFd0Hn+AxdaScY5FulWKF
4rH+Hpp7pQiRrkytRlEQQTgMwawg6SnpmPjhk6l4J+HEUa6Jm/U9q+zfs72/orZrQfyz2mCEO/gw
sdKIwyvrkdr8PQiCgypJZ582E7T9noVBtb3gcRHWz+FVW99Ep5zAgWDzNDo5xjSc8QpAwSUgjbvu
s+QtEtPp/BiaMipLHNUSq6LVJY+V2U3vNoW1UnxfR8RUz868FLD6n6KkIoFytEX3ZKWtTEk7tpDx
EBrES6v1R4MnZ8KFCCA+m9oA43FyL3FNVyzne0rpC5DRL35U4Dka2UZP7woPXBBgdgMJ9CVShlMz
Fp2IHctzUVzky+m2tGHDtxk83kFKfYkuyWe0QACR0S71453hbnbxKF/FJQqWAWaTBbRu+8DiFDAQ
cJQ0FumHL3LlEOg1oaYorf1ZRpyzeAOYFusZJf2AmHzZAszTy7VgwvmgWazrqHFl8O84SlFwUvJn
dOm4lLBdKUc7hqvA9rHFdCth7FF5tUaf1WTCc99i33b69a+s0X/8+6jT77AcXqRO7KRb49yQQR4J
MdV8zcpAVh8fzGWr/8u7iupdyN/SpjlEFw0W207Qwq/YlV3sbvvL88UN7T+9xlgPP6yemnbhnThX
R1IOrciSFSS6AF9feScDeI9fhQgBWcTnjwXESOE9C5/ILoA6EcNOOFbNN3DyLRtUXNmTbRO93tY2
ABr0WOSGsXYIdDveSSAkZJ3eBEFmqxXc857NPyMXWqpYvqHC12o2N0hYq31fAmZjj7oowKs+m92z
JOHSzv3J9tSpBAFKsSW19ekshBLjnPayF+HFa07EDSJhlsHz2fVHt6JxhSWFMjHuGrwQT2yc8R0y
C+dHRxIjT2kPwFSGK/3wHUhGHusozbfFQ/p9xaoNXTuvMiLs/P64evv9qs2l3JKZkMKOTXQ8ZHUh
r/dtJNj9bNs7BoMQp1sHoeLyz53t1M4nKOe/wIlTrlk7wL4pBOIKrLusW7Qy1l77Y3LE/KVGjMLm
N/dRuQ0hLGFefDRJjI03v2tPdxztcNcjtPQsbIw1+oKOEUW49jcyr7Y0Dm+IBsPktoTkclEO5fjV
9ifw8iss3jcdpoDHa2dFYQqN2/MoMnBnAqzJzE40lTbe8S1DIU0k/eePYmxe+tC1ZqBaoA4Wj0AZ
ZtBnhdOo0lVAk7Rikl4f6BqbROAYEX0G7HOB4o1HQNbfS9aJOPd6zjj2Dvxwlg3wrkSvssvvQfGH
0s6sQzOC+k6nJXJWaUOUTwVOakXk7fr5aPxYJB6ra1n5HzcwmJxAL5I1/sLp+iA8W9dvCvUMxGMR
skBVTtoX6llpCwmP4JF6CgDBCgI3pn369Kopu+VVNHvp+7mwjMC6T93Dt53oBol6+I4APNI37JOO
07mN1h/rZ8RoxFe/6tlIv7o3pxGySzSqdYo+puUmOoD2k20INYgjtH9ouNx8f6rTOGX95ANVOGVF
vUtaHEDl59dIiNOnOb4/5yJGyM/3xyUL16b3UOSquiN8SV+T0FfFRYvy6tdsSDA3AkIpaouGRdhG
WrmwFyglgLveil1RwpP94mdDFAMZo1rY8cnCpn6FdHcl888sXgMq+DwDETfQDQxEtGYPzS6EvG/n
0B/QP+9AgczMKXwh1k77opWXR2pFPBkutPtqNiSF85CB3yYM8+bnVQkg7KTenoZFGFwXmkoe/ZZP
hA8hPhe7Dl98yycxu83PZFPgkz4VrsyP4Uvsy/Q0w5mCYYKYVJ9cSHHP+mJYo3nwIq2krieu3DZ5
M/5HnXwweDHcjC/JSR1eUC7di1MhIEEO884ExwYjEk7bJiWOdu8myZQCP/iYnFLNO3Iaejddc/kc
BfJRTabKcSst4kt8qYSRVX9bjBiPBQ+4cEAsuyo4JbYdRosc2nbURy+6frt7NQxmGOH2OBQ5LY/1
L2TardjasiCNuIPrdY72vS4tBpZGLcXDOUxG5lEtx2ugEowNN0SOP0TEIUHDm1I1DPlfn/bQH0VY
sCLzEaxs4CrlMddPpibu2eu4nmvDa4bG8Lc/39LEk7aSDF5dJvKrr08MVxcaNNLZ/F+99BusR9U6
VOR/VVpXtTqY+bX6FeFIM+6wAJThqe5x3x8w0hvrRJTLRpJK4C89IJWyjMwW85Japxz3S5LGlz/N
VpwAguWfzbC4lUUQVWOAMPgm4nUYKpmP7FPhrGvrbuvUem44CuSsLcMPnmMoLo6INYehx28WKhqc
XQtNB3rp9kN9uMBpoRdy1JBC/hMUrnfwpz7mUj5yj4GTd0PQYd+WGIuPh6RlC1T59RnJfcDSB+1x
OWTnW0YAfFjfIjMZAMhD6f1z4r4hXyQtEM2RAUyBgjrPz9rfhtu0wZD+XradKIaLjesH0H4tHeKD
ZF8MH1A6RL5BUWRRR6Xgf7359Tuh0c4Uq52CpdURxbLcb6hwepYFSNthuOgo0eZFFTBiLr58xyCw
LfC5Gt2Dncny3y82GPZb36rF3B+Rxz076bl/PUPQ6YEABXg0ubVETpOnVCwKgWDJDxeCBM6zFpR+
VzCQh7dIzTVvB8gyDiQFmNlFU5SGpcMtz6JGa5rmWhxNOkxKhHytLEx0jOaz7W/eIxkT5VKbUlk1
G+UNuxLnfCYkipOayEScqtaDXZEay3uHOnGgITmbirbRW2GnI8rnYkkDjE3ujosTbdYzjg7LnBqV
35EXV0ikL/Wq5efLsAHHbGSUhxJJKSp2T/3WUJmY4o4Gd5OwaDHeiC0DQSZCcnVQDzzvBf5rPRDV
y75SttYJw4B3uR/7BPclEcwttZaDDECRGGMyYPeMQsRbr9YZl1N6eJWE2VpH0uT11+E63Nlw6Avz
Tus7devqkaS2oh8DmyNRJevFzswXPxbb5F+uL1oN7uzR2nyBlCI2R2pW3CQESVgtIDFCLGEACHGS
9Mou0/xNTG+IXcV8YChUpI6pXhZZnqPK6k8XEutP31VZ0KtWugCz021MOfZix6cWLoaSGDnX47i8
cM4cU2I7r22KHkqs/a9N0A0BBZXqJPCVB3PYIT2l3szEQTg8PAycJFQgbkw/qQzGlM1/GAMJ3LIs
F8k+V9SdLTBpI2kzkVHrBWb321+LLFxMwziT+mkUQKvK+L2GTR+P9gstdENfM2ro1gk6wANv+6M/
7LFQCAXR8GJqSfuyOmhbDtTWP1oD5FABHTYCCVdgPXCD1WPhd/3KgTSnFdYekCZMtZTK21NfAvQx
rlJE1q+x0L0XnaIMo4I6ANapWlHHudk1nsNe4R9Ajee2FqVmZ3fH6qAnsuqqo8CTKPwxtN845Gy/
C6Ya/XbFVwhCwYQ6pawNgP3CEhgIdgPgbbSkEW+r75km1G7Jys+6RpD5UrgSWJuT57pnjh9uYJEe
FNDxxaVqidk/zYHWOdgeR37Ct5MGHgicehKbId2y6odV57c3dGoSPdGWfcdpeknOmE7VQ8UGbNz/
If0iBrOgiuVhOnp3uFmV9Fq5CLnmpnxC6Z/aWiiFkckZHXMp24shztCDTEnv7p5ubPa+d3zQAcmR
UT59vN7vFkGIlTC8eCGq5a4i88jRFIe6eC5F3KCBK0aHKGAXcs0HEV/SAhDlT6NbwdkY4ui9GFEF
xsrI2qskOZkwivQY5npsb/yo7OQo3C/r5hW3MqXHN+NHJS0eBqkWm8HaGT5nXiDHOLXVoFBS97tT
7dyVOtVdkv4E/ALJF0ZAAyiKHQ7a+/9TKTZdNXvEJJksHrgL0aGrX0hMhVTv7H6RstXlxQGWHeSL
HrAZbG2Y8bB0eMVuc2fie/EQHXecNWSH6Gbc/GpE6ud6VkmSrawNfKBIS9O5baF+5BDigq2UkSkf
jvE/bdL/ebwXQ30Bhw6xBSUN9bg3URzKWjL9Cy3r9acLLMmG67ZYesOdlzbd38eJ/Rk92fv/eQVr
M7SAaUbEfWvR+6/7HYQjjU1hZpLwzOAAnR9A3KFNqeXq0OfrQsxysOMGweOK4ARq4E2r7UT3oSF3
XCnu2TB+qARR21jZYBT9mpovKRkA7QX/iYMKK2xd73jWAR6hzR5ySg9opC8Je/y9/Amtl39S41lt
drywpanNjZWH2lkhU2x7Fl2YE9wlEgLBzdhOJT9P02w1XPB8Qhzum4Ed7zVFdsAM6Qyqz3LuuaxN
IfROtLqL7ntUJn6N4sVL+okkffzNNl8AFxdUUuTsWWmgts7kS1YfikooMw4gfZWKcT0M7ZF1eM/1
CV+/iF3FBs4wTZ+4mPntR6Ge0zBsLwA+FFg3RnNnopkp7k44g5vHD2DBF/T3jgoMZbeFtexEZYgP
zK+UGQeCfRZonknlidmE5RV9ud9q3kPEyM/rNu12BkfoHEtIYN+YjYw9vMnq7isFWsO4FYAUAuOL
eBneHQFT4ZEmDeBFPwE9xn8kwkTkAZ/b6oxdlhBc+3UyXnAucXlaS4OGXIICAgu22jcSeencEPsv
nmKfEom0zMpx8RAVQtg9tAtw8CF0olVUenKS8lG6xeX6M5NVMZYJqemExw8OZ3GndFARt/6eALUy
AnOJX9ZXuXi/lKS1H4QNT2UCEa8Rrq4P820vGpRDYSox2O5o+0cCdZrSzCynPb0iIpObWtvtQRrC
BzwGj9FSBUTFYkB+WLgkQUqAFeWIPETUBGnqUwEkMo6wdnScbN4bf3qaa9zQbWutz7Nfy+R8DyJi
cxeSDmjL2/N0GuhyoNlbOdQ1s+KUJIhnvTPJnJqvNDoGw613fQuqgcTdgWophhK6AkPEgv1ZI4fR
xfbc7gibvsqE9MUqB7iRueZqEQQKvY7uwzFUgx2QbeJBAT+xgCksf5aPkgWyMjAGdXYg+NgllyGQ
sSf5nUsOQD/yJoOXUryliroZomPMCrTBBVGPOFfQ5rE2RRA554f2Mq033M4d4Q7zaWCHcwFAIQ9e
jUUXrhKxhLf9FDGZCnU0mMg+us4cKzp6fsizfFHIR1BAUnsB2d397TcPCY27/Til9Q/4RlDB01wW
g9VZlgWay6JHffbTnOdtFZxzpjYsebKgoLjW1Cjs9j7E7VDNHQcy1aySal/1w/3ybTzKDK44TK+5
RoTSvATWxlSOHEyW/wzlj/JDlPaN0Rjk63yuLgI6YDcK0WmON3ijaUdlIJZIenVKcdOChoypk5P3
zcXPh7AxIUv8bxefXYglu7TLIRg9FJ1GCIV2oy2srruMIyOtfOM4KkivPImYVbQaThhHoV1LWhKk
mLo2hTVmfXxFJrneqqtDujSRZfRD5oIp+z6M9w6qv6Bh4xZwvnbehVAtei96GQ6txTdQsBxNHFGP
riWISxM3xQp/CNydCfeYJzIBPSwhj6mRGlharQxf+Q/c0Zj18IUr6Uc3KFxBp97BdG2sXVE/3Thh
ltOmOmMy4myKqMRILZccxy9AfkZCsd+teFC42R+LDMdQfUDwL6/xVWSBlVh47eMRGZXLy5R78yhY
/cMZUD7tel4ut4Hy7IIJ+X8IvMjvdm/bNmBS5LMpj4nl4wVRzhFRyX8QCfzQNcC1AQSwkDnaXXAB
9S/0Xn1iUuu/vbx0gou3DizJMhFL3A/VTHJFAdlZLj/FYDrMrLKHPlY6Tv9FG9JTHeNnu5c/Bry/
E7LhvIUNaZ5XmHXAPOdM6XY74teVjNdAerDiKgg3Dltfk/vS4hhdzPVFMWr0hJkQYFlYdkQWwXRv
ikKkLT1kWQ9CdaNdEyoue0p/oM1uAEI3eiRr27w7eTZsnLHC2kwDJJ22jJY/W58MIDF2OddtKYaz
jtEPcFU/ktw2nidO8JhEUHEAJMwXr0c++oAzv3wUB7MdZrA5lLXpCrSpfeLl26pPYkv+i0kpyW0o
Lxnj8e80r0ROUmEMhnGai+P3yWiHVDd5Nv/ocCHNrDr7QMsI1ayOONUTIc2Y2dMriCV0HQa9fkEF
TKl2VnocNK6ANlhxamhBG4l2Vbt8v6QckBZNcXRxbh5WFb6MdLlEplB/mM5pZFadbg5H+x1np5b3
GejgKludA/FlBGmaM+sANFovH9HNWBiVLM/TfBKLcamBG1flCPoYXWVQHS8atTXwm2EKJBmf/6/c
86ggjuCBa2NpH4vOVnECW/7YsgEA8LVzxZBKNzTeG04+DcJaCpb0Yqs2f/MyIYDtnNkT/s+OxpEd
uWPyQAK2QiiPCEINPoNMKkQytM6HsK1hn51rDLZQ7l/gUpfff8yfkIv1VWYtCSH0qwqmK3ad3Fpb
4PLxi7FHJ9JTjwRuDMLEFxsWx3gM30l1AKotoyXMm6YH0c4dPJ+cC2/NNjGSs9AgbaNf9WkdmzaS
9o955ZxbeAA+zY83sm9zWA20HlZuG1Rr4a3Le7z/D1Kry3zamnc0L6NNxdYaaYymcvbWBK62lPiR
1MY0QXtfyxrH4X64gC8+p3IeAzYVm1z5fKD1Nx3xhG8Vj7Tw3fbjzIvuLWAaDRWAGrcFuUQLKZQX
Aax1GjrFbAWKyfflBqTJzRtHoofpVqlv1f97tt3thFT3HbPMqfKiOIU1nrmDvPq1MvkLtYdEypFe
zf3M2Pc8qjn2FW4I6xKG5yKrzcBlgjbZpDlspnWGSgMv8jFt8aPaep9/zFnu2l1PK8sGfZFXvt+V
saz7tzgGM+T3As2BstPCGtSWx2YvwhUhcQmjfnDoXfCrhoBWv1NNZ9jRsPI9WsV9jInFU3BI6Ja4
DxLxo1uH0DR3CYeeEX/ZYj4fqNeStsMobnWcMkOvEM6xEc838Ba17VPilWPKf3q9bvCNBGyuVV3N
+/crBE0ypPcKvoUnk6MSJfV7lXkDN4YkiBFSRBfWQ2mzlxmKuCJjHG2O0p4sD1hmMYmKcoDmuH74
uxyjOn6rHrmNlBYYBtygaJfkJB6roo3/5NZWjL9BofKuYOiFKQZ3rLW+rAB6kC19EjsMeAyHtDSo
N65GeqmNEC1i4eZ+MAUhZWXEI85rqMJXPnfxlbhCU1jBDnAAGaFhE5N9yhvVzbL1J7u1zsfclNro
QDrn5SABRnAO1Tolt9VxckiVw4cm2N8jtqZn13eVcOtFLvQ71SCwsiK3EyhKbUHBQDZ0vbmbTWw1
lYe1bQpvD+VRby/4WntLSTbQbEwznwYsguXkt9VotELSva1jfv9L8nd/afMPQIZZvCDDOEEPCAcw
C0SUCIphXvDDUP/rw3f+8SGvVSeWsns+j+WrG/Z1vvF6CR1BjKrFU+x/u/nYfGXguDwURxN8+AIR
dlRiY4/S9SmiKV9dANpV4OhHSWxb3TW0SHCSCeqk23leunr9FjXiL49cytqllTSsm9J08VjR2T98
+2qxM1viMyTVtxY9NLXRFKYHSFlA5btZsNLQEp0hAlXJXcZOfLJqYx0ObHL/Hdg/L4ecQkbKhtyz
8ZjEqkHPkqcuNZyMTWgoWZlL/3PGsh/c9YkUHTxlM2icdhXwbODLer3Dh4O2MstPtEga5kpltY6a
kF/wtloeT6MvKCs3b+RHPZOfmctU2GUNfyquW1g+0INnPyino92QoeHRzCfSwCrTWR3CzbTYo2CU
nTpk0+CJvl3115UoJuDll0sctpM/hJKMRZCZRGTZbH6yxDCnybEr817tXJkERS4lQez67EAMlwL8
sXAkFNX8D+8DNWNsIgnQFimfg1MWJQLo0vXzlgUEEhCoMhXwPfyYuO+3KwZg6MrR0LxO3uwqneCR
Z0qnwImcYrrYYjgSwrx2Png9yP7dGzXXlDndE13CyrK9fBysQIPKS+ima1P1R2Ko4g9bw/QYRzV4
AbXZLNSl/17rVu++VFEovGLhcGNpKPYTSVce1VdgDV7oFACogDw9TyGDE/A0BHfvDn2GQTQTht/n
BeEXMoxAZmCf/r1c7war4Rq4ZCBvW/mr0NJd4sKLjDtZ6PT21GQlm651p5hinfv48YFk/S9Ummm4
QtTOHJIs5gxWK2S5UGTlDgd9lC8dfRXKYN2ohpK2f9o875iaWv0yyq20xYCWJ8CuiUt57fKuc4Og
ZZXNiQFJjj2b4j1Y3S4NljIPQW8w1QU21CExzeHxtTYVJ9bOZv94F6R6Jml2hYkccKJG5mmsIp+b
8n5p9UHUl2EXgDnLeSGY+2snCYhw8kqUlof6V1Wou4BvmAMqtGDpRLNjSmLGouX+r3/llVCgIczQ
vf0PLpCqi7ZE/stFT/++tFMwObBfxTes7oCllZF9L/UnfB1nu4dEeBsVUQrR7/ZLUrfuJozvlQDK
PQbEG+uWBYe7WyBfHt5Xa8IctVDlVdpBaVVFWbaoQGe80Y0So7c6nnDNoHu+9ma8romstnlAqcKp
LJb606yWmSm4o2ZCTKU3sGZVyLSXX4Ok2F8DnStxOBtw8csO0WCjuoHFv85XAqK+1UFO92YHdspk
UbqQUYM7iM3m7QgeH/DRhyqXeOkS3HWvbMVW1SQg8GHouhL5rdy/S+Yu6gvJwDyZDHfDWKqiGYNE
tOye05U6cxA5RCUF37VV4HfSmWluRVBIrvcj2cauZXjo044joljAFaF8do79gcHR5Zvtln+ADAgc
IIhSLLm/5XOFo0OFqYpqlAvU1nxAo3p+Da/M6Xij6sk+NcHtPu2iNeMDOPQnXzc26nWnBpAGRCMj
s2PyDmEiXAFallYapudnH73C/OFcrzbb8boZrr1k87F6EsmuC8iQiv/NxC1z1tzlFnkTOPoMwMee
MbI7owIRD2G0LSUQcyG3I03WSN4JmwcHFR7qRsTtjw1Y0rxFZhXwl7KH9B3bi2UzPDZGyMOtBt6N
OgL+D5jN12e2HyNbyn3xpHLAlj6yqS/R8FB/6WE+xGQx/XalSG71SEJzhCELV5pr4raVqgDZkjhE
n4qyb/oX+RCZ9nGKGykgSR7FqM7RpWz6ht45V8xfe5FzA/37ebTnuursuZrNriyjGik0aavnlQve
qrWxcje5yW+M0xvufbzj1OGJtQXO5DfmBk7i81F66tTDPtuMXtDpajr79+RD+Cvc0+ZHSFn68Pko
ELcA9OuZWhTKsvfIY9ljwkeZ20w1106eLDHeefTYnyBcKzAYY7MsedsIh0zMmUjUzEBxz87UijGj
pG/JtIecjVSztfQ9NwCs25fQjqStAZ0ZWPlKv1Y+CngxVzR/oOrHwZLhz2EIgKtx+HnukOaoDI5s
x6TIjNushiksI+LhCMKVuLXAyzajJjRu/aMht4rFkUy8tFVUuwcomwwM6zWqdzrSk49WOS8Cw5a9
TyqHMXDTjDoGjEZ32W5CG62V+W1bxNk8p6Cm+03ZkwtCLezJNvEbLJEoVcWMYNp7jE5enDmi3/bG
bWXzYcbYu0UMUigaUllM/OJ7pO/sWlS1NR1Wymx9OloLEhvqD/nwgDZXJNiJMQlYyxtYMPkxqtpY
ZLpIoMXRIi2Yy0Ht2C83MlTBu/mJW57IuwjvMSrm60rWtqapeHKNWsNvd2EHXRX5orCjJO3QFn5I
I+BL1xkNK2u4YSXhSrlyU/uKjo6/Cb5jiSUWt9gsKfYd0Bs2xldsgWMbERuagllVYngDCn3Lpy30
ERPLeTv2/nbvpEGd3nzfXcz3BnbQVQ4Sq+NnvIPpM93j6BPNa3vv2tPzymVMSqFixF7X8g/mXwkr
oIgVuxrkYHP1tn9WP4Xrd/RW5Sy9vtbaryjQa7h8ncJV/0jGveef7GCdzujKOul1fKQ7XPQH8ZEe
5GG3x5pWDjqo8IcyHasa+aZfgsNrJh3HfvmUP5rSLV1QZo83g4lmdRw4gfBsmcXFaFeTZesKMlFB
wR4dLqKUOOPhPmuVEO3JaOngPb7jjLDTzZedb2lq4fVf1k5f8Bl1lR+peSnToe4/cf+0V0xIwXGJ
TPE3BKilc+WYzvYbo4oIL9v0yDB2fDbIZzMbi1R3IJNz7bvoXcsmKi3SSgKDENtaYa02/zoV5ymY
nLmN09uX/YqNVQNKjZ71eGEg3R3psLXmi3qnxKP0XmJQdL2Qefmd6sFAfZnCNcOVaq32tgcuR+ug
i1CXZaOMX9dixZ98CMrAZWnnB3fUs5HWxdszCkeJ+z5zZzHS3FEBRlX30G52ufLQGmHxcVsibFDt
gFUIwLqsSr84No6uPuQrMpswaYiOGOhEi46XrBmrWOmu19Z2SapHm4G1lcOSSfuavYsQpwh+obhc
CgI1Hv8u+kpv2sUazzJPaiA4BTtKhGZ69vjXubHJ+dIaTwPCkD9bfaRMw4FK7e4FAWrCSq0R1Qde
gip6CGa0YscsvaYZuSf+kHwR6XGZY5vpHzOoQP9HJpvqFN1vnO0argVpdBIcvoKiATJEJo4dbOhD
WFfGdn6xngylkbnRNpzSOtjY0j5DrkO+UBm/bWUlneRt0C68bgjjXnxdsNHZELVj6hvr6Zvv8vwf
lY8xnGDUXQY2FiRbvUrIhNh9YcfHKSNTlBpgmigMmHCEiZSPkHbONSeGUS0M50XYSQcYQnYQ8H0M
usDb9mECM9J2/2ouDNgh2RTXj/aZ6Pt4rMfIasPBI+fXhHbqOLbk0aKAdtrvUm+COiZxnHV4H3ht
oThanvFHWhj/HROSaxNeoQKPyCLrvCq5TrpV7zjbR8u7oxuBUKqOh152HtrRp+G0RXoduUnw5nlj
Idgaku41ls0+6jYBH418nlBWMS/ep5lWf3xAAN2QCuSBs5+QJ44ONWJpfv8uJlxjZQCROeNRYrJD
KSfYx9vNYvKaaIXO0TH1mDe1f7TLxryqVaoJBxKPYyu73utV0YiY35ZRz/B7xACX3p3R9wBoOlnw
1Fjea9qfoNKow5rRUiBA5L5hFM/0Q1YaSxZqnzwC8mcxZ/mlt7/60UlqzCoaU4ZsDdVg7PWzD1aA
vj5VKQj5Yh3XW8z95RiY/eYuKiQucJyDVXcABgbhPWa4cMf1HUW470OUz9edgPMYBKQ6vTnQ0gOZ
qBFGlcKVyz/M3DTpW+piRYCOm0P4WC1uf6EvyjXWdU1R/Hjb8St+n1l8XkldJdc92+trOkAJQ4CM
ed5dqRnB8hpwm1URID53wyqR7Ho/yK2wD2E3TPhpao0POQKXYFzoTZwBP+pS86HkWMzaAzyWlImF
9iqYaBwQSGUl+cs6xnV47MKzp9VujkxcaS0wOEcyRGRCwTeD9GXuYJkFv5IVVZ75eoAtbi4AoQCl
P/h1QPlDQjbmNGnxAQOshnyR07GhDt7ua+5IuT6Yo8hKHI8hky5tWVKniVTBYfR9/0IQ4a7pqq8l
ELd62r44VHh1w+J7ctlzL4yzI5MIsoSQ63OwdcGe8jZlJP2zYmvxtum8OxkAQs6K3hxGTc/2pC8i
y1cH84CnvKQGpZbEiHvOXiJ7dHlfv8SmMFutQApfPgRQd17bCS5NPZJqClk2NT4CPs6Fq60EwGG2
QnamRuQhCm7z9mKRiIeuD+niLhh9g7Vr+MPg5GBntpszVu4dG8M4QdzFyftk0xVFQMItP2GV1HN+
qBDbqrKja1QslYHE3BncIlY+Y7H80qXwYH+5tZPF5KLHs8BH1byffPZFaPM8GGhX7qVAHPpZYoxR
uGYVpkiXM6uNCWmK1jntJITLEhTsENXBFJlzmtEQ/gIHX2iABYIhPMFv1Ww2zgQq1iFoTbAfjFfc
g3ZTnWw4NiL0hF8xtsonb8TTlMPGx07wDvwancTK0cWxComNy2fwmextP4uK/c6BmUwjs039nev9
BdjZWkD6V1vgFVf8NGMTa89rAWqD4jZmFq8TdA1+sX8kmU2VzKbRV5nstThwIb1KjJzHqmDijKj/
o+qtV/3xLZrOZcOLzFhqh1P3rJFBp6CV28a6Hkfb3gQeTQlcWuKIGxnJD3ubN604h/5Bcp0EJRgn
jE73gHIKQ+70yJnUhe5Tu5Ljx0cGr7WaC+agJSeFf7TdZLM7s8jq+edBHKZZ+/cCejZxBXU86+15
bW2c59l6QsUb5av9yzz1SWmMoPynYiQwNgFHKgJBUkggKSBYZ5IcvKffVXyCE3Az3d00co8EckRG
r17yTZcd9LvYF4gilW0WQk/g/bSILcEPDdh2LDOAUZGwzmCwYts+OGA+rwuh3MIMTnMnTHP7ZzJP
AQ6rKaQt0Au2SeHrVIxKeHgoy5Rz8Gj3GKcOVj2MJBW6y3dgdEhi+hOhdTBS90kAOMEzOYP77udC
5VT+dyrpDd9XNNAYWwp2lzYf0d5C/X+9lfzIxNR+jVbEiszqoPITlGojVfcGuuOA4+yQ2l1N5I0a
NHgarRBtn2yIsE79yyam4C8BpbWbhQdaces1J6M3BPqi9T0nbFcTAclx5umkV9xh2zuXeDQzQ//K
AIgLy9g94iY5ljvmK3fF9BhhyIIU3dZx+ocN/IHBnsypgglPvmNUSLNs/LOQi08Ux5ayY8BeTVmb
SPUsBl9khUECs2HxBNXcbcboLeBydWgF816jFO6M57w8TVrYreda9E+EcafdzD7ZJ4TzWQExUunj
WRhhwbumLJI23WkLRuetGrXGdUgDmQh/wPmkjHb1cpRkzruUELrknysjCeNpr11KX0TBn2aUs1Cq
UiBU3OA1YFpvg0Pgr7LcOwy+OHZFrZeoS7MUzVvzAp3ZmImPYcHjTOEpFQ1ggGhbG2iXFLbk3263
lYPNejs/AMt6WGRZeFCVbtoyOTxO5p+28FZQw9dDblIFBZM2KzpAnqHGl+gZg7RY/h45NR2u+cFB
CHmJAVhM8FGoU6UkR38llgqrzwC3w0jMF7omZyq1zWl4OYwHayfr8PHG0jQql0LNbI4y3lIUG6nu
0Mp1/MG+4X1YT/iH+Kb4+cNq0UNLjB0ZDZqht9xE5QzrRgIMAaP8WwLIVCVExMN8JL1Po6nket/M
zZyHCwDM6eRS/4odIm9wNi+lZewWbtMHUJ7x0mXS8GNjD9ObAGTkC2GHeM7psIXmlHqnXir3pNyF
/LUB94TOZG3vs7PLBTKpqst5EFFz/Cy1KoBxd5sJvBQXGk99+cHyWuWFUSIs62q2WF1Zy8xqpt/5
Sh4J4vl1nMuqopegZLcbu8Ids7SLh5xOWw5rG5eyx01m1h3qTAVzhEf0bVPzJZQUVzdxMHrRfq/h
b52XyPRbj7D6YdEvxnsYFpBNRqYIvTYb6/T0H3toCA53kTIVRVrdUkOnln2LhPyDm5++ExPPZmLN
46kMB9DWAPooMcp3urzUqYPzZp/qPIFR/LRM754DGTjP4ytg6wguhJtgH3iGF97N2seMiCMGJ7Or
QOr68rRx4Y4jejiHFlcia4TOAijxRfcttqghFxd5U1nMrbhoGwpa9LQWw1b4s9FAD1yR0NbAcdVH
Txl+pgEs1lZdh06AHdjvYpMDHHAxfmyq5QyzVrqbITt8KAhXfQtJd4NXgkT4eiS5ZwKrfRTh53R3
aoT5Cfl20/x4UyM0FZguOmQNqInH+HfdbBwXVxx/mEPTNgPN519bzyuDy/HvQRPWNIIepIkpfRbC
Hek+D1cJrR3BTQIkJkbSwOaoK6c1+Jd/MY+4SAugmun3oW3Cvfo99w2UvvDSMxYkZB2WzPshBHNX
EcxN1u42mtePNEpcMromPEqIIocCj08Kj4qIiUtfDxAGrtfWBmjGgWBG74Bd3ClTSq1pxRxgVHC3
coxWraplWa9GlErsw+CMbOgaFnJYZ0H9myYa9fOZH6fxpnqmL/zf5U85inImfz5EAXKrWW7RozBR
JKXkkOieNbNioYj5xM2Nv2m4FTNHbRjCk9VRd9w54EDaBSbZgBioq9PxMtDvr0IbErYiHXIXEWoC
mHlBeu5/0BtClSnbrhC4Gmigk1LLZJ5khlOVJFxJub8RG8bAaGBH+58NgeI3/GYcRsWvEYFavI4F
IWEMPnE9dKBniLsfv2e/KktJqggn+dO0cTKBPDSXdE8FwkXvyUxGST6ZqStDPtvGgHejwhO/z63M
eqMhpD6Sbzwct7Df09Nyz7gj3vsoaWq5jO/ZU0VbM5iu9xg8yuJRt+Z8nGyhwdDRP4rhUNyHSclA
Qux/JosihQrbcLFB6imXxLQBuskwke2t1iRSx1+EITpU9+OjJkeC22wracqxqI/cuhYiuBrJ/WXB
0MYJzYvgHDxs0BOWHbSaXb5tFLiQotkYYVJj3IQPntCgcbE6AXEShmkYzA2DJhpVyHnyYCl0/BQJ
bk4LF73IMOskU1l3rEefpEn5oZAz4jHHhUcXAro478i863Qr8ZlRUUYoX4GL4gLf/uwaD1jape6z
0i6opJtbUAJ5kj8m10h6qQs0NjTii8+aO1e6+mxW4v+zXUzv5nEb2jvGBSqbPHaveZegD33bEzU3
GrRr6zebjW97KjDju3zZVfsTiGcA3XEnLqq9qYWYSzItAa39FvI2hpOloBKtJ6tZy0GnlyHJcYEP
oycRoytiXvFJA6HajsHfOPaAsqWtZIqa9+BI+FyiDvUX6s3dzwVQ2L+0svnlLSQN3k9fSW1Jd8DQ
XVQpun9//Kr/pUUMNm14BRUkMkzA0um+IRyaHJ/Sob7m5HDlrPmps5Z956lCZuqtsBVB+bOgJQd7
3+gfwU+sAEWiHoG0lrLQ2mp2KXYXW5T1TIhOAFJi5ccy/sFLbFqvd0m4ghR4FX497FyToa8rwyoP
i8XRj4nMckZQ/aLtY0CXKeZ3gQzGYjjrYUyM0k4PGqA0/dj1dw0TO4WMTkpi+RXSHpDz/agApH4I
h0qtINpxRbAzQJMbZKcW78ju/Em4YO3T0y/nGa7Xmu1iOQjDc6c/x9Jni6/B3AKKUTALLnA0rAvh
07DO2Bv1ysZLcabFf73Q3KqIeGMJVvWR1jJBQEn04S5l+XhIfTKgP5g6DZDfUhtjDNlxPkpRCF7S
b9o6dEdz2zTmsg4uphfn19PT/Ygs56mLD46I6v/ca1t9xTWYy+Z++cCY4B0jKnecgaDrgWG0jY7D
//WI/OTjOxckBF0pnCLq+mIxbpBngGOaOQKp5BQUtLsu9EG2dbjEtsaxBQkG74+Z4BTW5F+kHbdW
oHzbbaaxfl5dBLnFPvOuM0wlyqAg5M8N3szSH1HgrNDJTqKBXKjtR4ia2w5t/H6Yqka92G2TjKMu
p/IHjptaCSPRundJsf93vys6AqNDso4DsVUf4WNvI3CZx+w16NmmSomerTri1VXx3X9DYpL0QHsA
OiZFyy0fCBWSidAIsM4eTHvad0mKxHGlZguyswTTMwvO2UFraQEirudw5QvkuyKaAAdaRrzF/udt
umbvUVKQE8zEqhU9Oys9nLajhXljhuPmZ5xcriZQ+ZbZLIW8QY665SGVeX44ZEBJueLLryjCiOz6
z97qAT5h9rb8leCNKs3zKKXIfnsctUz1q904GCvXENxN8R1FJpyeCxF2RUaSqQ1fYrIfSLfRxMrm
SCj0E6fdv0icLMwMdkASZ7/1JOTocjQ9fSAm1qCCqQ7O/xNqGAXXUZB7+W7Yil/Kku/cD4YhXKMQ
S3u9Mi8wHKOko18hd/SxQUusKXNuwObWhzkx89aJqRFjChfORO96JhizCFlEjz5wb+/0BBIUtp/4
vNAb8v2oATDlc1n4gh0jVZ1qrKriMXVBeXlUy7J9razS4kEBM/EMqyJHRUrIqoj3Pxc0/IyuFmTi
ylxF6ZRx6nwnge1Ftx9dH+7Yl5ccdA/98QdrMuWwqyTL28OnD3KQ4hEUL86iMZllzq16CYHg2ih/
GuW+BChNR89za5Tt4X+S7Ygz+O9elbXUO546Zzyxryfu9AjAT/81/LzbyhgMJqRsj77gI3KcPI0I
Gn3MwGxMKfkUZaATM4S0m3SPoqur6YrFqSl35ZEbAR06BGT7fN9ZNya65fWcl+SjzLVsK7t+Bg43
55NIX5C9ASEf0nDxewCJGK2dPLM4Qwn2vIxHoPpkDV5d4AAG9w62tWbRCxlZyQq60HYsbRH5eQW1
3Gg/5HL5Kqg64yQd9edr4YGOow+TDD4GvEhcm41uq5h9hk2hj9q0WK5mVd35AO25vy25Qx+mVzVb
ild1KH4Q0mNOEzkqXOO9sQlxOKK0BPxSvSO+LvDARnFcMr8RTwcu3QYrJrZ9wkv8Y7GOwe8ERv9z
n7psOh0aLXkpnxEJPJg+LjX0L+iLYIAR9LMkYLNMjA6ZXPfq4UQyt1hpgUAWv5/tGqMfUrnOcA7W
Sx17f0lfRLCfcDPfkxfprwOOzkvd6JTGsS2wdoSa9qxGaT5LUObr3yf4PcU/o6MsSqiac52Bcl9z
S+BcTNWnpw/fiNq2BXztVacHXN2IEu3Lahh4kKCCCq64ZESU3GPSEXb1Y7gqUWbg475fpILbJPMw
j9DWWqY8bNVK2m34SQuZ9p6i4FJW0FVD9plLC6usWLw8EzFWacNuLJjVn03HM5TQRFOA3VymLnvK
dnoA3jAfqDJG487BD1VOgoTfE9PzNz/iZN2bi3g8KVKYgXlz0Xz7pqSzBw9hoFMEpQHbMu2jH48l
aRWcGF5hqQXUQwYxOLqOpNNsrifxoyhZ9Op/YkT02GQtZXQIRge52sDh+mIhrvM+KOr/kVTb/8mA
1k4OL+44VXrNo9PLqbHNpBejVkfusBeXAXtWLRVsAJQJloMmadCymNBzTyTuxpBrLDYYz2vh/le3
WCjVTvBLobv14ow72kjpj5jaj0HKc6pOSHZRkI8QYxtx8MJG09VhRISvFzimqNXTjA9VQHjyl2Xj
uBJ145SKJfZwIraEb4P8ymyNrN/+CPHGP2sdNEPfXBwi2zZWR0C3rUK2HHEtak89bUNkV5pJmhnu
UbIT7AmlmWRw6LtaqajosRHGppZQq4LQ24L9xV+rG9b0GowhO48QIL6SgmecgG1OvG17Ptve7DpG
o9grrFhxHGl2akyD7b+qc1IYkxNiMnT4ZX1XVToYIUz4qbvwHWUOs1djysDDTxTom68CJf+cXwwe
ktTzlIJyClvuTz9K0a+2EEqccZzoUi5Fjv0EeO0zB5vCb9sIU3HuPfOm7M6sDCxxDgxk6v6T8gS3
48nry/AvK/3w5fjYOp4ADVLl/1mgNLgSncotcBbYTsdgZ3gUph+8JtEPP2tIjtWyrztzDUdR7cON
Iv1tno5S3+gNv8BJKRMZnDth1T6LXcX1QhP6sjW7hkfU/ipRwcnEA+qD35Kw0CCHXet+4ouULELD
2O+P9ujotbutWkvvnki1N7RVUUgaC1GMiWlCYYvJKNkleAPtbej4zjxjk1PBNqbzbN5L2USVjowL
rQO2wowWD1o/Z2001wrYUyfT31/VesQXbePT9gokBHCTsMvdIWhWAD56rL6w7/1l+sy5TzPxN8eC
xZlbKboU2Ji3FOys5P2v1xF6+VFpEShSKoiM5T+O7KeNDnMr2sMh/6ZIVjVeeg0b0OYQ4hC00FEm
M3z6HmwF74xFHNtXFcBt5zVYTU/KnsBRcKcjTz/SHXmqssLNLRhaoKo7cvGNnrNWHClmlRAMZFhy
9dJtwzZwM5ROwZunZivyoz0tbR9vtfnsF6b0h4pg12XN4BxSbErpOnuJPVVMPPzR5MjU/Ta1HpTI
t5NrR+mzuHG447WDKDuCk4Sk0aT5YAAgEFFcsUq2PVQmnoVU+68MtgBnkVxlGd3b8EIzXEXcyFtE
sHovQo/hT7VGdjDa933Jtfu+Ny0BdPq0mRao+6vW/ImBghdnvPCd9p0vEtmrsu2iLWY5mtPd86k9
KZT2P/TqJA9Sbn/CxxF5YHMsFhBToOld7E0Q5BHtCtrE3EKKP8rSOpLJXGApkH0SpmuL+notZO+2
M1pa4e9LqPEqOo4sMTUifxeyiNo7lFZGYI/g/lrm2+RftBfsYpYMjuA1VY20CMNE+nl7WV68WoZN
8k7Iay9o6vcJujCRv4uFl1HKdxqN4spNosd855tmuDF8SPzoByV0hbVduKjaD2oimlneI7UK6Z6t
sTvQnJNLhya1PDzl2Nb4oCm87VnJ2DqM5ynLtsx/4FU4ZMKEjBIVbALLoxanQaF7kNG5zJVvA2ou
ZpWNJbQ9LnaMVTF09fLnvrr+Qgxtd6mfotBASFHuRdKr3iJ+ahPKGWAMa8IF8R0X7OAuz5queWlL
eYWjgNx/SIuLaohA4KGN7eVhcg970f2lLgL+jL4AjTa7vYl1PwpetJ2nNmLQlgvugKJwTUNTe4He
/0CaiRz7ugb3mRdHpeBisK3/cSwop38Gne7MPZTsnYKNIaRYOBxz+Em8Cw+h8JjXPq9ITLNuPVRp
NGHeURufAzjhVvpybbuxp+1lQPAL8WAvro50jwb/xewD1122iX/uFkg8CdVNKw2vbdXKrvweFnpy
jfnbu9EENOw0+/NP9fCTWwWvIafYaZo3n8aMq0xBfJJsYRYWq4SqsqR6L78CqWhXQSZGPSHN/JlQ
4EtQLRn+/t6S2QTdeRJ3gcMK4KLlhxhuZmJhQC6WuVmZ4ngrqZN77U2OQs75xu7N9xN5me7vHv0g
8tV2fZJcjMI/0oajPAm7zfoh1grfnoqQHHK9whZVCCFeqZsgl5tQHSgig7OnJ/RnEVIahfNb1uKs
cRnRadyHhJ1MaAGtUpt7P9Xd7kEdfKG1Ch71Pffyn7rkBJdf/VV/f7c+uFzXcMPbJ63gFmRurMYA
zUTPOeSFq79vm3ZEZ2/TdkikABRzgVcsA1lB+aq0UDaSlLy2r/rDjKixp2XA0CTg0LCINqv53JV7
+Dg4MB01ApgzFtmpm1+YiJCc9TfSmM1RTuWK79/drXz7v95BVANygAJ40Vj4g9rkqqRBhLwsVBDr
quKqsZKnrwDehzsQRIVnIuEvr4QiwqVec3QxALj8oltejVjSA0WSyXezYEKcBg5DRkJ8/jLp0KDA
IQUfAmpZZVLratvah1eqh/ltDvPN2GnRDxv2JZ0ZH8TtwBap3JXh3UW1Auyj80vVLMQTLtGjNLWj
ALJNlVR0cMTjm4LFkfxa2Eg1ZXpuelPcRN9xXebbo9yWxxDV9eeTWR+0aOYAFUolgAi6EhJWocQW
PevYEwg/voNdeSQisj2mWDG1zpA85N6qu9hAQPljYCQThzHduLFDaHeWyz9FRDVWwixp2kdYFcyh
HGrQf6rdoJpNLfQx0EqZM5DYRItXoz4tyhT5xyzKhwN8e1hBlL7CNwdIlUF0N4TQvGP6n9SfRqAk
qFM0cDu9Hwfst1sIDbg9d/CHuIBEzI5P1Sv8Dj4Fn36EF2pc1+X+nngoLUsCFi3CmSUnu7ulcKMy
t8l7Dx5LegaRu0HSWYYdDCmqdXFOvclNQN+ZP/27mJt2RBf95Nj+mDZEtktWmj5O6CZilOVufEAo
WyJSvbFWOChvV20fqPjI8cylhF6wTZcoH/magTURMQM59lZnlcSMIGP+SxbjXMKvouzN3VGw7aCH
uv876RvSCqaCJuWt8IyTTc4M2NJqwKzZttO8fxO2X76cYi/VaBrqgNuDTr/fsf5eoeFXtpxVDvD7
Nh24vENThdt3T7hk/3LXJwB56QL+azNFOm00ysgUxc+IV2iKdExPEWBue3QVlqNEmUZLv503eEgV
qel+pbCemQmdxi3NPX2soWYQMVGwPgVLPZW+VQQcBunQZ4MAZXfLgF2w5a5fiU+5h4mcQdWMNSoI
7RLbKWVaDqWwQHXmqHCs1gkHUj59fBQmnYpa2wlm90ND9XegmzM06JlM73kFLtw8dotXr8Xfz08N
DLBQN9zO7ugwOLWoE+elyZeIR/+3Zj+Jwv6PBNukoiRBotWDzegoA0nrzhQMVS9u1yIXouDm/72p
QQB+958ztRSsiiFJm6GqiRjcVMhXrZtdZwEiQwUk3Mhp5fGzjQ+bEeDVE9dz6B2+Bi7MDCgBnxO8
f0rcDpzql1pzJEmffqouGKFZqhKXdFy2GUH4RbOw4k2oPEGbLZUlDV99S5nN4ms4dSTB/22rMPkt
3g1nLIKubLTraiCoclzElApzbLFbVpNf8EUOASmQ5IF0wxBIoWOA/Yoqw0GykqOoQh+bLIk1qfnq
c/kOE1MxnCne3Udzf07zaJtG0iGES+j/RG432nU0eA1W/4pGk1hGAiEBV8XTO9WiWLzYOKtEl9OK
1R/MUYJYtWUFhZ2TWtyqOv9CMTf+666navKtQaqsg3LWgXv7+vAPKMIVHlycXCRhkRv084pEffzm
3pt5f7uMJ3ljbe0Xe7EieI5MBU2t5RF2kXqrjFl/kY/FMLuQDCHOktKzQduypDOFEjD2EVzyDysN
zGZlu3im5NGTIn4exsP9reMASP6wM74e16NEXBFJc1QhF4v0eAx9+d8zB7tp5H0LWYvoceplAZyb
RQ+o/jc5bt1atrMcKoNTVBeA10gzXRhQS7sP3aTgkqMr1L0wqbhNCMUUTNJkSiw5G/uSLP6nSzGr
Vwv18OZ9Pz/RY/jBm6eGFefuGdexB+Is8kOKVZNRcDWqxuG+0LZdo0ZiuwYAwLEcJk9et142qBij
zJfvq4dmUQ1DuLJudYVoR75Gfoz2pFZe62gvcivrPrr8ouQ3uz8lAAjl2IreOp2hjLQJOmrNFTUu
e7Sugc0NJR4gqrcjf80dD6yLD7a/icK2TEWY56+IJoOKioCDMEymB45+2x/Gj0a4vOrar3fCmOeO
UnDG8D3CmfcHJ3d61RRMQtOw4O0i0mbO8wwcPsZ9G5JAWxCN5eDquFMeXVpX8RhQj382du86DP/9
6nMUXjTuus1+vUAdr1DrcuigD8wcGLrKVUdMkY4pRTR15tXMffNF3tw2F2dO9VSJ6PolszhuAe8R
eNWjzRvwlau+HlDkSby1wdZ6t02/s1K/I2Dx4sgUTH7d5y/2RIxuCUpTwE/ZNrYbgHa+qKf0teba
OuudhJGCHd6kJ1neAymliyEJDpydiQp/PfsiEQaneoACqfZdROR1xQu9IVLBZ9KS5jV0xccR96Do
X1sVUqF/BYGsH17flZ2UalZ6/0aEB5+V+NxiQBz4MBV0ik4UaYxP9dvOK7PcKSg8JQpSwJ8LQQ4O
vxyXLbBScdrLINcD85d2QxTMi4jAVfvNyei6UyQOVWZrkSqna6klVUwRIaaBE82bRYdUhLhYeZD2
GjUl/hRDdS8y6xfYMzFuVMksq93UD6JxU2dD2nmYaR6iinFHXfPW4h6TLPcrYcwm7G/gmXiBhEsQ
Wgasu4SsB0b19/FfNfzNwUKDcuOM3Wt0wVCBcCcqOe2oV95dkWA4YrgZxwLH78Gul8uE4BvJUvm1
J3WmcNzXhGCt3EG1vlc6XEa41PynbjcoTXVwC39+42CANhEUHUtwZJiqi0uUDnYjHzm1YQT3V2OU
89Q7Byrd/5QtZN9rdAMuu0NEV1yxG5KghXf1Sb+FUaUGQsu4nzOjDZIiyBOySZn0sMX+dF6hx5ev
A0fXPdF+ZCBZbXcEZLxe3GL/i8gvyBlsO61Szus2J3hEia8JfYZuUdbPikk6V4mtFZ+eu7OFmUYQ
SG0Dv5/1x1mE4NeLCwlxdQRteIJi6pJaw3IanOltOk7I0adCUeASb+J99yvWOgQr6UuN//LphJ1/
hXwTunfilcy9wmvNqvot5yQV1hKBoRIOJacevM2wg+mOWn9H2pwr0FYZAHWomJrCXnXqquN5SSpX
CL9cBH2yDjrUyIPaOB4PGcJywgko+UGbJdsvPAN4AR9glsuDC/vXshTrNLJWIzCBd6NLHRbRGw21
QpaZ6kqxK3FA2B3JZFePBPrxfGBO/icn3FtleJ8yasfZ2pxjN9QZDAAaTKnoFz49fOXddY6AhBRB
edkFvhJKv6/OiWc1wxf9H51fAR3JZGF4cMJ5X2UIcRByPYzI8RpOteX9Im2G3Yx9WI5M1kxfC1P8
S4JE94Ec7VbgstnGJiQWUVAq2QzmU7D77Dg12AZ7AgX+xJHX4b8caVRP0c4AsPJj+AMFHHJ75GF7
fyrReMT8uN3ybgkC/Oi8KY3umc2xmmHY+WEPXQ9mkh5CKfxrZn9nMgLVOsUrNQHz7WrB1UH2OYjL
8au0Lc5XqKyHA5zw1+GW1K979Ne1T6Rv3RE2J8GKJvKlPnx9CV/+Oo4apaa5hJXOskNGcvh0gLtH
qGeklXaSQX5JoJooCnWPG0rYQHW5o4gopQtSXo8lhQofC4352/GcJcGx7aCroZfUF3wGTcF5c6Vm
6l6KJJq5joTeym3pvTjirRV5nt/s7o2KhBGuD7b19iYmTJJoqI5ZXXNMsGk2yfVZVPsyM+y7Kn2i
ePllwu9geRL6vLwGlX7GaG2hEIjI+dCwhefFy1roW8RuBDqrMHskoNCOBAakXpM5JcoKpPs6X2Lt
BDalPUyzVugLAGTCE44P2JN1TuuBkrGEnxeCcLwUyfQTNEXaH+SaVRHfqNlBPL43ydt50mw34TmO
sWioaPNitKvgffIgTacPTPKjvzAaI5HoQ6+kIGSvRVmftRkY91NA+LOw1whwxnzsfJ2sbRy+1Nuv
hj8YKwo279boRT6qI8MEUVx4MltQwIBxRTaJfErgQthdRbag3XX3ekjetipr5zn7XEKZOSftNtQb
X7pBwvca8makIwIBgVchi/JgzzmOeaEtegnbtmt2O35iJC2fd/z3m113v0PcQYtJYQloQ8j0Sb62
vDok6lsS5URl7jw62NxF13lfArsDR3Mkr0kBVUwMvEskJYxL6r5qoF+gOTRePvDt3prXat7iFqqv
Cc1eFbQZSfaBjvrQWZTgOLsorwz7X32l3iGzd9ZCzVNE1f8HaiV2yPpiE75lrHMh/pqmaDmGwej1
nLEJ+FUpMvY9hUDeIFdL4RcrvaXc3ffPzGDjSFuw0WSZRlSnHzv0LddEniwYNa1wcb7Ap3qVeSe/
4sFCG7eIu+su8SXIhFJQNPT/S72uuaD2ZTx5TssR0KRxoEzYwf5H2ngLuEpzoLuYGKUpzU9JSrmi
PeeUjZD3Okc3MkSrm3ic/pJQVjiCJr4h7xh9cXnizKKBG9iaSKc23fzXFanl6FF76sAC7/ZxYObv
3W5rm6BuBU8YyE+mvE3NFDbeZnbNzvuFKG4Ajfu1mTpqaM75cbg0jSqgsmsfjL3XAPO52HdF6jRm
IyBYao7WdalfVapkBkKlAShLfI4bxzmoTYa9x9NKODFyWvHyiu/JA5ZtzjOf/kL1GyBBpdUy5XPq
hhaBfLVh6QnW8ZuV5VKZ0NiIQwy0Q166EaSRsm5G7hLo7bV3xxJSKmlT+jLz7WDXp+b011spg4jB
Zu4QPkVW4MMADhJ1IRGpN3XnSIllF0xtzlksk0+gcBglmDcTog0K+YPXBnkvTux9coXIwx3jLnRi
vwEk+O15/SxvxeZf375CCQ7yKOYPFAw9h0uCvnFyO9FVufeskU0GozNJiBfjoPNxo88hMqTrP75p
kKUygOeLbnbNS4TFezZceP3eQtAx790hbgWMNj1HCCEe+6oS3ykojT66THxOLC4MV/G/Y1vsJh1b
iIlANYbi9Piulj/+F/4+5MEfTHJoccj1/L83q5RpHw8/Z/qz17pqOCek7WRzbPrmEmj10S/+Uqb+
ZmZMNhLryqiCYkNH5foxYrzgfyyqLNTQxwggwCAFZWqAOCbfUeYtO5Ilb0SswuJsYUA6pH/PgdOx
GBHEf4J+oYIAmVKF1aep/Ep36nEDvtSmaJShktN+/Vrq1M/A47RikhKe1YG+O97VxO4GTyAUuMat
TR2qDO4SbNZRhZZf96jwksvAjBVvEmfZlPEUx7Z3Goivr10kJiRh3G/bBwASLLa2Y3j8q+jVb2BE
s+wjlyT2G69SOOV8BUXRXXbXOtzoxYdP7STvbez24zgX77rLMHCcdRa8ANadbAWN6EaLIuuNN/XA
OKzq0wi+1YNAaOS1k3lOd8JIdmKixR1xBrbg92oS11vxLckQq2v8Lw9YEmRaM6vSYlNAgPSD50Wd
lSOzbDC/VQwzYTs5m4Kle28dizyOYQoIABzWsqBVV/XAsQ6A+8SEERZnK6qUzgdAXMGMyL4yTknb
+NfGY44IixmCHxs0bVt+oLeJgNi/4PagxIdtlz+9iOkycaV9cSEnxf/VFCMnkf+J8KaRYfTVY8iG
o45apP7ZNwSMtYC7k0rtGfIBFh9oVvCXZAlU21EYrW1yAB095DseyWg+EJwlD+1rQKtyuLMBPHUp
QzjdFTesRZ8Jz2xbbZ2qJu34M7f2Qx9fCGVNZuKDrCc/xBSCZ0bSFlOLVpm8M4xWLIKLLZd2a1hy
1DxztCZJGFpkkWpKrUdM1jp/onbGhMKSPD/0NbzjqCw2dt124eQpFYtawmC4wuEJ+zsfQRpEbimJ
iRgFvVmg0o5IaqX+kdRUJF22ame7OL7ksysxNid1YneGhPbsAfDOx9JXtWJJdPmL4hk5DDMQXhZ+
1mXgqejx6W00OMbM7EKYztGBf/1b0UNSBMDllsTMLVpmIfgQvKsS/jukP8quf3q7/1u1HdKAhwC/
jh2NolmlqB95iJ549VSgg7YeaQx1wOLTOewhtDXlCS8kukG6Xpo0Fyfr//zgBeOgZmofk5Ef7QQ8
db2EkXNGsgsEtRylcIAYiYOlvzl95Imh4hvAvgYVWv2CfMbHqpmdE6z/T3xVUcjwYRu7K3/sZCJG
Z8pyPKisi6g93bECG+FQGUiKMAahOtwRB0e4PncVdwcnz1tNuK9V/Svjdnfy2whaCjRVkYCCfcU4
FAq+wa/g7dW/7efvUtJo84aPXxEeRr8BtRkxiIbLbGtaBFr1s3fDRKDTrvVPO1tiXeUv/EN8j53J
5AdSq/YnMqpB3enJyksOqzj5+XmtVEM2Ru+xm2j/ugMAaWqRETTBoLuiQjI1jGKjbwdylZtuIIBY
clAFEVcGmFS2aK4zbrbirsGi9ncYgpqO+wcZdBxblLHM5cdry5G9gnvlfKninTfRPKFoSnu4/75D
Qp3CmeZFtUAGBhRcOy72YaQG7LZOVjIi8RXrVJpvYbQlLBoDI9P1Oh4Vd4cS7GerqUYoGVoK8KuM
WzlIZk7ccfBjP90x11Rys+kopwrG/gMySOz8ulvSRpDec3uFDDzMO3O6SzJPWGQbv60hatiisUAF
buS3qkPFEHc+nYgMwKfAvuHfW4HKekiSM1/PrAMpnGT9G2PaVEy7Y/ErdRNPi4CPuBbl0QqP++6D
Tj45kz4A0UrGhZv/97qTE53RVjvxbJLYzzzR7N+E1bIsntkEfaCCaAOG1QoEUPdqKtq4ShSWRoX3
JO4jTDxjWYD0Uk3TrQdTz3aZYDK/9ATV8RJG5m6rlqQws0QlpX/Dn69yZ1ae372deya+dD0UttrB
7G+cv7FPbQjQ0JLpBmyLUcQkl0lYVGkCv9neIbrHEdoitzgf1oaQKh9invtibh7zDCPL+6FJhy1B
VTsT3v+tfGAGAWIeyF9IIV78/i6IEykb21F2jV/scB7Fox8oC9cOvje5nVGceP2HnTBcZccWbmVU
usC/0EzEUmvyRHdE3xaDiy7HfEv5b9br8p6kFnRdL2NavJvhJV+S93JYLd5O7JXC5KZ1AaWYvwq6
meDu9aCIvSYgmoD+ZHtLM6KTSA12DrZ4SIJwo5gQN1HDvMlFfFD1MfyMOE3bTSEkDDwsM1Kn6+YE
h4yf4E1FBUDmNxzn0sK6O8X+MABmGrWu0KbQG+xO/4jrbSHTvz+G8FXxdbwCDI34XzRK/T1r7KAP
jj6cWt5IZ1BRp75zZWmkIU8LlhfNMKQ5zY+JG58oSILkpev/ChSt2FR8fQjpDNeIM5xeCPd+4ynG
ZbzmC6BTwnpdfb6gbswHzw+J+lnCUTO/eP7CeVgA5qmzbF3R5g26XJK2vV8WPy76exsxLqeGvcDa
J3xtwgLDMZes8reXG8smBh8CFUQjvMNwTZZaybGLWBr2sf+a/2XfPU1CJsRUxuM6TDUgIj/UVUM+
bv8gxv8M8jZLBeirU5Ou3xUMgckXdpqtunYhbSUI/NiN2LANPnejM5Lna80edVfdZrDaGD3z1+HB
4q974RfDxk+Xeh7MjwJ5shXW/rvt7RzjoKwoe3crf9vw//TL3DNJGF/FqwsHywtfzuezBWycj+bZ
UgQ9vmkfrepf9v+zCd3Y4mBk3F1Yni9LKagoFrOc5pZmmcUHU6sGUhNqDf1SSffMg6/ok2agFx5R
5i2gKFNhzAoB6IzeNFVJUm91kE1XeueZQs2T9SAt+XzNaGpxe2TAgojFMmJ7u5VUm8gN4QXy+ZfW
VuCiWsHZUedS2dkRjOs8L0eWKgAQsv9xaMN+rF5QW1F3Qln4tSwFuU7YAs5/8sPMsv0b+wyu9Tey
y9WPUGGMrtPXp3bYx7m0utf9z+9K2jwmS/ehaRiNjDV5k96oKC6X+IHt4v3BV2TJtW9gFQEDD1a1
yGSxdzL8KCqUtsNAkq/SYp6dsnI0qs68eWSKlBnUPse7x8b92lt6sSOtGI5VqHxLifoLcBmrDQyb
3YFctHusc1AfERCGWgRLtNr4QsLLOD9SMtJ72lYJPRURFdVIGZbg8hgEiMLc1mz4oJnQYHwxJOcW
PXGWGtCUAL/obcYBxBdlfRTjAKHnO+/5SjcbwkC8Dm2+CL7va0yIObsfYwD1rxctyWYZsNuAKbKI
LDAeopDFsT/mOoHureBEHrOIX9ufsc3Ql7Cart6YGHPKLlDWa9uzoEyB1kAkkdQNP5Y6FAi1bDDC
w14PdJgZYzAvuLh5g/GLc1jE3E8Iv1ROQsjDtmS29ck1UOmHmO011SDtMKkVy3YEdaJhZ38hjHte
GhDErebhUivh9F1ZkTU93Fk1Ph/iZh5Ogzk4qBXBI3PV0LWsgJW56gZMFYpMK6PMKsx5REKLfYZp
RJNhC6/sV23sa23GfTsk/qIvn11TKvL7rFiErhgSrG7hBp5Msbw8Y6CR1XQa0Gyb4bzdttTPnYRA
qXSx5jngf54Ym70g31FMnr0lTshkxY8UUYVlgG6lBfsXZ3VQyQLbniJNKjy1HVtD7xcTvSXRkEIx
0ztkhX+59E++/e9E1B6kjTJ2spMAjDYLqLp4DLMNpMTgQKdYwje+MbT8ysRhGxaMeaG3c8jX7qL0
22GdyRI1DdxTTDLSlJI0jq64ZsFE7Xp5fq+c44WpItrEJj0HwuvxyTwKz3gdb2RCtRgq7nNs5hLP
ArwLYWEc2pTFKSXRuhFKJMZteiYOtLqIp6iuo3JBAR7TaHL7WLsypb4q+Kfx98r53REnouosGL+q
59OcpMZa8+z462bKsrNumrH1dCOi9OBz+o7bpgrHE+hlkIx1dB4iyiAeMfu1BxKpZAfz4nXpvZmK
LTKoKhi78eBDOseJ+84jPAt8knKM1zovb9V4Z9Anx1Mqh2WpLf34zmZlz+tV1nzfDEZTJ+ZqEOqt
UDmVL/mONt4ZM3XU5YPEsQueFeRH5Z5zMmMj9k7AFVsSRtPpGR0Xd+/lb1ta0+ZANTNUcJWGPWAK
WNsyyL9svUMxDR1wtX7oGC3psgaRtPXyHnxcfgZVutuF575OS+fL7mmvyhi0vQ0OLWwwaVFUvFyl
NVTO8Arz4nUz1LExV8dIcDrlqbtQCHW6+MGwOWEkoaAe4fPQioMwA9EDGyjkZoKGeOkVm/xxXvqo
gw3+7V5kit25HUxdgGTL+zRNHXuudMYIzbUUTIT2UpW3K3E+C6kMzH9JoF2TBFrn0lwcpIwCS6TZ
7ZUF3kvk+GO4IxKGxga6fE1bQVue6B6bdoKpohNEsAM5nSngZZq3ZQQShyRxCNgLwBppADP2JNl1
KA3jUFN0mXBDMbp7E1lz6VZA1QOmYmqgNqCy2CkrpV/IQGgvsFwO8rpnEWyjBcp7A/w2K6ifNceU
dZSHIpDbARHwSlEr3tsaZxHdbP8lTNefZ/rUlG/lp9cchUQxxeGSZ3AsNlARUoCT6/VgEr+KhOYa
hfJUDgMY4KarPkK/8yB55TVRP8M6TJlHHmr2VFksx+k25lv3YAFpajt18FtjZNvqfp8XkjlVpABb
VQOtXp2kBn9veDakOJdqaowUx/9zNB1LQCgLqMLvXoHwlqli6BEC1TStClTvMcVxe2SUoPYcaFfn
2Rso4KjNZQm1aco7Z/kBdpkg1c3fKUpUc9v858RdJDIjwwWNXeO4FaPshiiSami1mGL9gYeR4KD9
Y0UR+L5OqQtfuMCYhzsyCy8b5/JWxwJNrLLudyPTPEyomoXPMjqsy1cvAEpEnD1EkukXkGFvxCSQ
JCl0Qk59y2JI1kitVB9XDdwY7vCwrq+FQJUxMwPitWPMJm31mO1dk8zUZUxzTHeiJRYjel35y5Sr
4P2eutnEUgh76s2cslro65k7VT5FRGDqCpVS4R8i6eh75ZEZfLOo/vez9mClRA0anJOVa1B2J1/i
SI5PZPl2O83NINy+SJqwBySRnbDGlgADny8u9eX6HfDkQ1QSrLNENIM6GSUDpjo88w6gNKAl0+tv
F4zVEZPk6N5If9vK7bODICBs9nrBnojn5YwU/GZs7BeqQzDJLCUb+109cSRnc6nVmN5yiqfQBBh4
B5pP6PaQlKnMsOg8oMxy8dSNYN7beXTSgP1cDU73SznCcoFhSWynAdCHQGvQDKRe3JJP8nWk7H19
ls23w8jTGLf/vcrzSZdb3jK3xuZ/v2S1HVzUynRhnUpnatQiAybpDcL2Lf8d6nDZImWallDnVSaR
PWNIIzV/mNsPBHHU3Yq85keuDoOUu+ckHoaOV4gIvFQqIUOIL+fN08YrZ4lUxXbRG3T2l1XFnkLt
AshajzOge3omgcl4LFTfjKljZlbD8b4AKr7Pyh+DMYz5+l/lZ3/Qhru5+FZEyXfPVzaxfb3oPm0W
sinINAZBCjnq3k/Ovvy7R1DDnS0sPgfxoY/98EEi9JDS/qP0smYzmpO0IHhdCxa4CSV5qikO2FAT
QHbk6wbIkRuk/S6mUnQE2T1e2aFa+uToLqsVYAEx9zQStEf0OwFvjlPsrA6LRcCqIbsi8D49kO60
GdOx0YzmFmFNUvaZ8PmCepEjT7JKjSJLR+G4dfkksBLivkeQKgyvUYkyixil+f9RPaaJQU5ztHQN
mwnXrclhCMLjqfFqsdf09GMMzDOBT6A2wSH4iQ0c21/Y0ex47zkc524iRqCyied2LWF15mEHqHGu
G8TZtl53L7kJeoMdC7n74uYcN30eCBIFXJUxeRxMXNmoK4QisQO84tK4zc9qiOd6Cu4FRpRtZnWK
JbV1wJpDIkTDTP3uOmvkhcDSYvZNY46ffJOpD/606IcY6Qypisiycp0UfVkME1syM42j8AdVuDqS
lMVH555hMP3fc8zEOecF/IXivpR59K9G/1Q+s+3sf1153JAyoXz+CtGqix94Ji+2mVrmiPbWvS9d
C/4QgQiVTgdDz9JZvh8eMf8EdLjcrL/Chh9uHEmpLQ53aRkW+HphG7Ew3ZOOhDR/qvYoLssSt9/o
DvHJ1Wu60eICSxNTfgeUGHWL8JTovAw2Vv7nlvRhFi10k9TRBRosx/nw+h2jg/xPSm4V+QqgkaE+
dfCETXpRZfK1Sx+4GCm8Xj0chcPpVUt9fUZG6zpSF8D5VlxFPJhRJrn3ED7rbETwKLKyJ0+OvdWZ
PIg+soh8udcRrdn8yW/rk3fBpeyikkYEU5uTaWu82xink0pvylSjMV0haETY8yi/P5uOoUAh7WNt
rI43/R7PDJdpveEqpgldCHbFqotgEExGZRr+tg3gdZh/doEY7Y2JwuIyUDZDZqxznVtZiUuJns9q
ZY9JYxwKFjqtnbrneIHfDW0BlmIVkYeBtFBonAPLGi15//VVDS+KdQ8rxRStvy99Tyli58iQqPwb
0RvGYd80QhvXOVeraRqHyQoi4KS86Nx+EErDuh8fCU77Mq5meIsUlx6Kmk7iffczGQKXZ44wEB0S
atx802JFrxOcebakrWivu+JYN/E7WFPu/cfE1cf+Wfy86HMVHWf7FglM58U+2M5GFJ8wMREhB9HC
kLcX1cbxKrVk4gBuJbyjlKjlgJYJb/POu4SrAg7AfqPZIRhJXcP9IFQ4hjI3w7Ni5sbBWjnA1ek9
2gdmAlpjhDW5NRKCg6LNlIs38P5EGYHCGpf9NUNNUMCnCgLrweHHP32erb+5k2h2MLLGP5YkLsU/
JfVzummwZddj/53SMHQhc8347XUZWHHZI5833eBuzuRcf8y2r3q8Q3ykDpUPaKtuajX7gDACMTc0
YB3L//hEoUyScx6QNLm7g4rZD+dL4rs1/yrXjzXxbRfll/gGU5N9CYPj07DXeWoLPmvXnoeXglE7
bXn40zdQZbbMEzkW1wcwQS+QYYrn0uFNrtSH7SEyIcTNOF7NxF8pZBvl+tHzQacQp8WmXwm6PVm/
9IC5pC84LChOQc5pWe0yP5Aduo2tL8q8YHhifEOhseqJVaSHIB4KdwDgtV6wvy5Bzo0iodLpAIhz
SUjWyK71n6GlRMA9FPk8Atw22xvxl7vB2BpTGx+a4/3xYP8BCRRm7gzPsfmwImawzUbteY+e0OES
gmK1xkdcviIc8BekhuyyGsp3hELlUWx2c6b3rf0Q/Ych656XZoh1Ql8yxrxQFf20PhvcEMJT9w9F
qLLwYAcX3r7I12a3iRLlJSyhTI/F7vcbmQ6c9fswZ7AoED0Pd6DaxBr/eqDIGgiUaTB7zCzUgaxt
hNoLT8o1spC4OrNgO3OWvaJ8mxRnyZNLB+6a4BsBomdYLdL5i3w0MvF5dqR++hYwCao9hVZ3WisD
w246IA93gZCj7k4RjZbvaKDPVqMkTmU9qh4iSp3sP4T5aInem89AN8Y/xujIuDuwWlLmYy1HiYh7
SXYol34y7Rau7MzJ6vLA4A65CaWr0Ok112zwtTFMTQoP1KOh9RaJCacf1Y3RNDg0i5eHWWHZK5D3
IOc1LTli5X6Z0XqM8mLN1e8UlH/yOof2gUeV3cdj4jkXGhV/GBdoMA+C2288A/NB8SI5RBnTc6nR
Wr1JJn67VPsCc1nZH+3PaPfrbkWmlyKwaE4aj9L4TAE9Dm1IDrBNtHQkQgVDTWjb6yrXmSKneXL7
E0rqdzbS6FLYImFJcqb0iX9KmM59I9tKuqSydWxuKBPMSeGYecqD/MsbW5722pIhlM5jaRdJExLE
NkXgaoW/nj/RB9kYbaWhJKJgqmuhR6+ENhW2sobZHC39quIudIH1b6Hx/c3N8EGYGx4iZcOzFh/+
vT2rfEmBvdJqc/XVW0qZcHWBi54qiin9OQqT+wPqljq0KyyfKX6Kw318o/fDHA4Df0844v+WBd6O
v11Z0cx70g2GDC6JXXhL1RyYj58+Y1kJu1/ewV+3SD52O9ML16WWQrviPFIyLovMG42trBDcqb5b
GkYX8e7gi05ujJLsfIEBlkkUikSEMOPeo6lovlKqbcSMr+anv6Z0khENhsPaOCIUv4NxRPqBQYDR
rKmxy/63PoYGbKY9BRJoRCYJheb1m23HotrPsQB7dkGwDOLyM4F7UtDKWW2UKlCRRnV4jo/V8q3q
ehIbwXFBKzrR5Alqyequ/mqey0vd2VtVoKOrcU2Q81uKj7m+M2OCaSeVmVBQDYHHMHVXUaaXMsNR
1LMMRD7mD0J2nL9dxODRts/aTCKDmp3Of3m/b3issRVVgGsZXvEKxnvUuBYxLVDWvwTUZbz00jep
7IcgSAOAjWziFZY9Pbi57mmiUKiiARlVteMp7DkC6VH48LDoPgKFdVzFBwCVpMSrZo2jOMtnj0+K
aX1rIT+VQySN2R1nJJm6RJ9ho0rIPAQ6EcOmz0W9noJg8I5q4af/T/n8JBmD8Fy5IXTFcncS4Ea2
jVzbey5IqRAlBzF+kns0Eh3G4su4xRyJyk3DzxaYJzws3OBw+uerDTvix9VGjM9Rimqhx7Xw19zS
ied7MeBfhBR5J+WivdLdznWpm7okVLMcsef0ZQjKaoEJ66hvMY7Jsy95gkT+FLquFqwpM6QQUrWo
Ng2MxjUdicWL0NtMwCNjQk0Cnxz3CGEYGXfHvHH4Udj5XoucsumaQJtqMG5Bsmapd9pzgh4CMEde
jYNquyEKv0/+v52Jzo5E+cSEHC3bxOAAANiP/c2tMjr1qCjAUf//FyyR6WwAnuYA4vlgzgaxwZam
rLSPHEFngHO3GDpUmw09sc0kSPFuKTuQH84FgkH5RwWCxsLChe6PEKASKl6sECYTl8r0bBxfOWMN
6rXiYuoOCLmAAb/kSmyhC1J66ZtR7GZCGMPEVstJX8LfjhZK1WwHoiBMB93KQ82hFqJUQgm9bW+i
jR/L8jsQ/eaozLGbo3ZLa9VOqY0ZDhvvED/0vwkyOsUw8oJY7t2rbYymBY7Oy5CIlRtSMPYxHE2y
/bGloSTUGSDd5ZqZvUGAH7+ZBrEFVvxLbF3eKgyciWiPXO010Qe/uYrhT641kqnnTldXsQBYXUpc
KhL7dvCKv8DLzoEJfOHXIrjvQhzkrByAzTCifVKo8lw6HAJUwFjEn/GI/SYjbfPAmo3Tl4ovtrB5
tsZimPzC7aGOGpLXjsWg1s6grSmg9UQVcxOcHl1Qa3lvcC79SDV9CXAlgNgM1ecAwCj8iCnDLyuQ
3G05i1Zag9qdhDtub73eoudKEul/NWra1bfjB6lk9RS5kTvRSZ4SG8pRbkx70CSOcnDwgz9zjuse
NpYGygxQ4sy2Eg62A8ic78j3+4e7Gu/54FUTxF5nO57MNSNERbbHqGynKeDQAhmnyz29nf0xhjtm
yzRMyuRRtpk9R6UK4koryeDJWVA1q8Ty3qgPXVpXlPcxSTgbMHAuGu3jPFPXwwSbToLtlUjQM2Dj
7pvHSn2PbL4hRf3tVCAFAenHCB6zSGQqMVoDmu7HGhU1GuxRALzAlI7iNBt3IL2sGa2uEwhcnc+c
YUChIHK70TbjGxEeYE4RD6ol9DmscGa2TbcguJNLiH823gY88YAs+B8CSToM9gmXFmbUzxVuZ8mf
Y1xIoEBgCTXvYAzTjkgUXwZjCB1L5aA3jHb5Bt/bFCoFq+8A+CzfRXuwMQUwz5BBgYuiEkCSORy7
gGveQ2UrSWRehcm5jXLawUjnPzsQcNhPaQigjM6Ch6TDaGZw0ekoNQBo1NJ7QwD2lKYudLFlLZDI
0fI11gAC32dOyD4Gs35JHXKJs8RtiTYpbiCHquMjhHx7EOw1ZxzwBu0kSKkIfcAGparBsSI5wWvm
kv+w0NnLtoctFbShqyzEsE7XcLEpp/jOdQe3W9BZWeBT8h19/tk4vUAKLaVAhuhnLq6DC7WDaz45
MW+PaCV0TeB5NYPonPXQ+jc+e/kGqM9yDdx6npfoHJhway+/wLBnK2UJuD/FRjJaGa6lWZimpsHW
halvn16AkioFnCllF5AVq4Y3diXmDJSBi/nRrip9YerSjZY4vlpZ3+ooGmTRondKqYK9zlWey1Vm
18SLK6sdNk4WhKlxmTQHAwg3mTVLnVeSCD/nZurdBqn5HaWK1zE7t9QmsEzsrFP7ZERaeVxtL49B
X9ZkUxkP67yKi6CCo+iOpGWafTy2GZPBs7WKPMnZaCX3kBL+jhtwE8ZWM5O3ltc9MlVsNJyWlpKN
0N39+Rr8SpOgH8FhORxpEZIJ+/Kj+ND4TiFfv1ynNBNaLthd1z7qXOzHiWC4cakgyTz9awFFF9LF
cJkYuqa+jIY6wPmNH2b79mPv84H45ZLCtrDfWkPoNyOKWHXkQHOVCGOT/QcKotHBvncNpZbFsH0e
LzRw5fwaDcDECzXRj0tvuPLCdoP56DQy9Q0LzaB1xLcWS7EW/w0bDY3Jpx1z0IdmLOB/BurWuv/h
T3xBli1zTtEOHkUx7qqQf4am1NzYHyFsVH5uu17/xFDWzjfNdM/MgAJwJ2Mmgqbw6Un2ImdXhOSi
ifaqMZsaaMn5ODArGb9s75DzpEvzZ7tFsRb+UqJZY2ZCR/a4tXeY6K8V5Nf4GR28Lv3t0bf/Lz+Q
xIcfDrKmrnvNlBxzoHzht+pW1MA8lqXWd9iuqQtIK2aqdrQtrYm66J5khW43tsIpKS5nJ0UKtJnX
xE5KgNSmlurePyX7wHeTdDXQhPgqNRdOJmKYLRMlJtYXBkrJuVm4iyq+ur+JREjelIyATXTvor5h
VmSiHAqY66EPCk0ATUGA60AnoFKYPCs+Av/Zo7iR/X94S5KlgPRha/hu0/CgXte9r5DG4jfW2QdB
VlFrQ/YnxVLycfQbUUPL33a6UiDjcnvDFPj8wYyokfxv/LlIzriA4KOOk5i/vROq5tPOxhNmXJbe
+VnQgTwVlcGCdqRwkg7M6Au37cSL+R4TM7L/6xwSEH3f4c8vITdaA/d10LRNp84NJRFcb8rjEhna
poqXfVCRcIcLC1rNQ09D6XE1KumRrlcYmM7F9CKBZHcaiYUe7rvLRxKmJpTi3/Fh6lvY7XCN4bbS
f2ZaWNT8Jmb2MDHVf7vE73EoliJWCpDYpSSwo9fyA7NiarGWkJKCYiwMBgGsPoBxIS9eGPMd9nDM
NKPCsmBO+TF47oExuUHNvCQJTnvis8OjhCRrlT8+RjFUZNcET6SjRyweUX7o93nTFbXEk457M31j
UtQPZpLKh62rJBQaHWf4xJqpvProsEudzDtoSiIvVv5UDSr1MxZU4j79Bkb1X1URSlfM8znCSdEu
rRa5cmh9kRmjCPeNBOxfC5bmc1Y+f0lihIIEdr15JVqAHUHWDnlUwVsPKuA6vHpw2Xb8O3q6Nb6x
5UATe7ref0HRABuUXTdt6AF3bc77zn1rFW9ADg3ZFUxO2V4NN5YcogGUYMY6/U7r2DLy1PzUPxAO
hc343gsksNTwmdRkEA74g4Q+jhoZh5B2tvLpAxHEa7fHNFjFhqzP6gk+tG2iLFqkDmz4HODd5oXJ
IS+Z5t2bzsJKlZyJ3Cb7N0DdDhUJNzUD2SUzd4zWBCBoBi20bVMF5mcVWORtHueYikAmzfEMP9TH
DOWMA9XaT3Gs5/OMo8LBYAMY9dx+jqe+3yLcQwzUMHEDlBdbfnxpe9F20q1tMslBS8Zg/YqTlXEZ
ho0qOR2FYPmS4W5l1oYwJIokJdPdaZePDde2DLhiSACMvPEZGMqtKwsNVFRgRh9XFsR7slFP4LQh
LvwR3Xi5SlOXwITQV9lPsiK3wqxngeaZU/SUpaatzam8p+ZLlON7DK2/oPszTf0d4uP4OAXy3FNk
hH7V6SKwyIBgSdw67BcG7exdKT7V/WdO2tETwmx/vbyWvY8w2LFwN0NXAyyTAyvUXw0hqfnWyiUj
tdnW+qJiJ+G3MiFJVCBDCCAvKxTv+Z871p6o+GgS0s6kXJoOiCCLbGW71d2x1ln50bXxCGSWscs+
m54IHPKJmy5EGwJ0k1SO29ExWfIMAAONbptgcEFLdS2dbpcrt60ZH00Oxdl9Kpj0uDbSdMG0r/RO
S7zP1PlllVQ8dwLp5ac7ufPD6t2f5eyixsFWy+Y8x3vqIyIHOkMglL8z4ty9/HXK/G1jj3zNFLsv
AG0uBWs567g4g4mT6aYvQ1e3QXS9N98aWCp9mWG39IFcbxGFBUKTEMPTyHOyPfFy2lenLA0nuYGS
LxwS4omx1kwSYYwdTjnnkpTFvUFOAKmb1QPuDtEnWWwSSZvKVfmp8oL7NyKoW4KcxwdaNIjJ/9rX
afRyK6sADdyXSeg699gj0b5Rc9axo/Xq8Uj5yNtZ7mb4CBIkyD/+nPFCoKJbiwF+kP+DJtdh5Ah1
zG9vP2MtFu1ZXKsbtV/CUVAPIibHB5tADieKVqUfyPD1DXuPZqrrWPNU6rcz5qbLS/9VyPljugMC
RPniqgcCLBym7mIz/nnsdJZdDxzy97uhM7NrCTDR/LZnEgbqQi+KC51M6XIttQV0q9dRnntu63d3
KUz1ScTRVmKCsgapLB1Tp+F8ofbFUYzsDOYmDJQMwRPfq+rXp9yI7aSJd1Fm7KJw/8cXIQ5gdSD6
SnyZSiSq451IsUtDVpvNjIxkHIyu4ndKeM3xdmu4uD8MJfe1NRP1pKZelU9R0q2qOxvyE8W7Zl8Q
NBbzQGTHEZDrfl/3zuCddLP7YY3KR65dKcaNZEukC6wK6rlGnQxwfcggqRgzzplbKOXIZin8uLhl
UI7Wez+Bffgldjt3ecUdBc5DNr5QEFRRWc4eLZqgIY9eWtmZ4WNIOf4fKp5d3MRRGKOUK3JZdGkM
kqmKApTaQd79Q5F5qYiecnOLKbcTeRPZ1BWW9GCMuzN6SsSsM18m1d7pphDaEW1rmRvANLRJ+LWL
lzQy2ef9TIWZLX4sEgRHnPBkniCF8oxQTMzjwkZ5F3SQ4q5g3XesHuSj/QDnbIMqG0Cx0XA54xAb
CZn35igfm8e04d07ajVNVEAgWlMc8T0IcfRN+8F1XLeMUOF7wCkfqagoERu5FSslWGsAQ3aCFKqI
OHipIz4AAXP9tHwaR9ko9RfoalLRVOs2mIrYEhnYNOcdpIfTmEDYObBFGA8ZFtjp/IoXCm/mqtra
hYNkhjoAb9hbGI9mFiTlSLJFhnSGbbe/7KaRjoyTPSck17R7qsJLUVEpx7GXo3/SGv/OQDp6vbWh
NiDkX6/KgC6cn/lE08GxJwayqHX4ykL39X9jU0S1eaG/t+s3hvHwrz/tiSN9r7B6mxd2EJeihcZH
L2u79fUumKN04P3NSXxZvd0X9MelDIXhHa/OWtYTat61YKvhbSB8Gvbw9BmB1hhSOeVsci2TEY87
JzHynEvLqWALmxyRS4Qi2b+t8oTfeqWGJnNQ9AItUVAEvwTl2Vznm0oLaF1r8gkVNQVRS/s+g4mD
WcPdFEpTrsjCgqNplZuHkyZke/6bywT+/mADyDUiQXNsjvzNWu1UQyA2nZqxSiWQkCHIUs9enPmn
3dd1hRh5LjL9R9ayxFhen40AesJkcEkEiq94hM43+q9BhJ0LHw83LTu6qa1/cUAysPN8Ftbxynyg
yD4Tu9jwy0SmW0qO0I7VhCjGcZlZLEmgMg/srEeJCk/OMyoAe/cgVGz0pYgr6/zTSC6q6FlXw+QM
xOwy/USI8gcn7Ni6lBvHqzrdgQ7IZVzyvjKTMPS9cW7c2tWXgFcp4vUyA5Og99dYeLLD07iG/jyX
UQSJRm+cPxqyWuz2b+gdfLVnVpqNs2U0GYwKXJ6lRZVAKWYkc4m/X6Gk0LYHe6eHyl2VPpJ4c7Uj
o2ecBVvontI3n61Fu4LNTGoISu3GPXmHD0b8HhHAycg720irlnZNnqDLRXXnB95iWdfa44WNnWKJ
r5hog2XEz/CXk7qQm3+/xlzf1WNe4uab4qPpM5Gr2psUYeySXSBULA+4AGpgeyebuttnmHmzyWoy
fx5fn3BXpKH496YKtZ+xqelvLUv2jyVBwnaoS7FU7i5zwbsKYik3lrfI7AjCeJ4ZH13utw3Ka4ub
QdReoIvHPy3QQoUDdCsppDEm9yX/y2lI1OfunbrA5hPOk61oVKK+qYwzonjzTdjtxMn2NrQfC5wo
vGgekfb9/+NyVLHOiDR0uzLTSn3Lq4fwDG/qrkG+tcrjAf+7OLtLlJr9P9KrattdUTVRMfW0La6c
1ABx0+SRplNr3mZh3tpLItdzds+Tm33yDAm8qqRwV9Vn6+93QlJSjvzVoV45TzyiWF4HpLnB+ke5
4Gc1I3ApgqB4mUI5LagJXtjtbVpuaHUtPZaoyxZqDSZgmFXfGz5e/qM5Es+WGx+i2sL5eilv2hcX
4zyk1/Bqo2Ju4nlM+gWctFhTOzbf1pe6Sd2b2dCJs5amew3dbDpN9AKLJh1y+dnVq4KUynrC60Sq
e5T85RaNGcHMlZzrcxGXZ4F0F0x0bLPBCBJD6M1glyQrT07X6CEqtM3IRHZG/DEtRIbF6NNdrALe
RS5FZYQk1ln+3G99S5LAgxFOEcjtEHzB1x+3ylupzYX1KJqg3a/FblkSf5hLLtlSDQR/bgYNyh8g
gAqTBT4A+bvh2Ln7N4VhQ0b1fVXY0nXis/eIg/TrzHiTf8cwTlt3Yxz8vLN+7wJmmiuhOWwx0gTW
LUYhUG5Su/T/uS0t0aJkttWwvx0bx8NK3HXMJLmyzTMGd58ksUuAOFEVdm7ZX0xOT3QZwZ1D9npi
qsa8BfUgkJgouY3umFXRt2JNRSMD7I8YWqYK4QckQ5jprGAUcAdZyNfWYt2qsepzObN3BMLPhxx5
WoWT2QH4PjSdEM4LShvQ0R07tzkrvCPDhyBazaC3/R4mxZJ2bEk6sArZ68OmxT0t7WpsWlS2ZZxj
Kp5SJqKGHWKoa0rYnIe17TywDREML+ZdFG0IuYT5mLz5T53p2C4LaBP9LqoV8lvaRNy2dZPM+1rZ
32ALGsbdHLu5y1Zb/6FF0xL/xqcG0DehQT9Lz77cACrPrcHPHIDclTfYAITZAKQCkn2ONoLTrlzd
WCBBsUHAhz8sLJiLKWl0OpNB6G0yT03Tsq1DjfrBSbuFTq86JNpZ2xDBbBOpEx0INpo+tWeKiiTv
KJ52/dplGuAO2QNQm2I0B9fBZISId3wzwBj6tmQWLCE5lyPqeAdLeuYCc3emsZCw/tZKOBpEELEY
h2NYpel4kzV6Dm8uTNd3n0hbEq3VVi6T6yvtH4b7TETq2Fucq/m2zEHREandvo1LHnPP4+QIvvUk
3SA+U2MgJHuuvzYNzl6qYP5Vslosj5NXpdeq3dudU0C9tr2ictlquwZHnk4IuXuEc2UIbT60xH7b
G3yHQbfRLGWn0X1y5bGR3dzrPSiHatB0GqEOyp+HD4+0SGef6JAnNZYzxOzYQmIozEPU5slaI1bG
FOWnQyskXq4ZugEJVll0mbexsJIxlQNG4OlQ4C0k7SLY/x0laILQ/9N5m4nk1elth5j89NnOt6a0
i4A20z3jhXdzCO48zaf6Le9k0GFL1N2IiHcc8t1DyMCZxg1Ramv7o5cet5DlbvuqZ9wEIy7I8XkI
5MdXTsLfiRxBv54bz9Twhz7KFLjjgyd+JovlxKyZ+HpiVPYToxDsjY/ZyrRa8s84lfERcXBi6u9B
GiewaLu8n4LvhsN/w8bWu0wUwolx6yNsEly1IzGtfrnU+F7tk/rVPwuTGH9B8CITv1+WCqDEPq/0
eZj6RxwC5KtlU6LoVKmeyYMp9zx4TIVNpaa2d3M8H5vd2wQxmNomykTVBriojbu1TGGfDdoe8YCK
4oRD9CQAhbWP4mpnCtK0gh667gzJ8I2eOEWfpeMZMQNX99bccJtwPWI2bStrAWBvW9SJ+ki2ffP1
lBRbIYNOo8uJK5wWZVz81pxcSrPL+i2Wi6FR7FViTZLx5jfhiY4iAaLCu88UtK2pVEpHaJnAWr5+
SaQScpGy0+KbULUjeB5K1o4zUiEZsUUbbA7iP3hSaUJQs2H9pWepEygnZJ+WodQ9GMHiJny5JcL4
T5eP+wEjJHGljC5zBLwFfs+2yU85CT1OyKqEYDjaf0rH1hip6yoIwCnmjtfqv1qZW6uB3eJLLTJs
ih2eTJVUvd9CyzTxyNx+fdzZnR0jAtu2RWb+lcZqFGI1tZjzss5k1JNLwKb/UJwf8hBDAk7TYbOP
YMqHOMp4TD2O6TUjmF62wTjY+vJ4lkr+/A/x73Ij/T7I8/Di4AjV9APxj0J4MP8UzPCOY45HYTaf
j0fOpwtbaPo2wivNzQFRuKrxm4z3UevyJqviKwMGPOoXqDpRLy5YcmZMILZFORS0yLZcOImGSb6G
uLM6QBRdNJMeW2pJaEPgr/Dpeh3RVWf10t7vsajxi/+3idShGQzURip42VxUz7AtMuXhKD+bbQv6
EzFL5ipRCIce6DkH+Xn4iJUqT5h74DQH1X780VfxSRGWSYUQmUWfNENLw6OcNzjG71ylCqhdOOvy
UL/yDnVUCkfGQc/gk/5X+oXXfivclveTfYfPztbSWEE8kRXrd5nzVNlSNeFqu0o5n+OtNnj4u2gn
GmGFsmbu+aCbZiWgEMVRgZxdVQ4oxb20QbdzKPVdrhYEO4MgHUgFeG9FKTzFM2FrGQV+29tQn9Er
sNgd7AhJNXZbXUlojOQkpSb3WgYwvJOLYyMtmrJX67KckT7WOVfb1duv+p6AUpYQHzEqxchNZp1z
u5BjfVHel3HLe1IU7yiOb2cahnT01vlnglX+8ECKIHgq5/pmMANDfYHC2C2M5n/CjKSYHVuazmVA
ProDPnGFJUzKaRY/Gf9APmQvLdP9+57lO4Dcibi7y5JVkkhvvMKPq6CsNW2HgPEL/R0XuPhRdili
rW40lVnzrygOKMSAhszu4XpU/xPfAXuIZS8mC6lXb0FPpqdaV4K5/uv6ajamDOUvzYvXINGC0eRW
baYeCkHgd0+OUa4DqvCPh8oVJ/iMKhjVv/+vEwNZAjt7uhTELR4Rv/uFmYtVOpM8VTml+3rFCOtC
KP+Jx69jsF/N+UOaCqweHkL5p+g1F4AS66YkOGMjsAGKmEAL8t8VbpiAlyEBcUeSDsjaggxXxL+B
zmEd1zBwGre8kPGJW6Uo3pUOiib4KDp5PJ1G1JuB7Xo3wznKqg7WddupD+42rT5KYR/uU0hg5i13
zHQVRB58osflzfFlgo27AAYEQ121E4yhUhLFPq8KhL4uGtTvmS4Ai735grxC5FmyGst5hHfnTu3+
bPnvPvzRY5D7mxjqwrrU36PSLThTju/mRtpJ29rRQk/TTL5hmN2M9ugqvEnHf1I1YPGpF5LCgWCp
yr812mZkCR0GYFib8vvVb7xKCqUyg0ypccvnH7xypufOX8wdIsd6Tr8qW0bgNFvwZWo6M8a5VhRh
G3Ce3kHL9ibZATnMwlJKtYdWlauRBrp75LECMTIYV6VPmgyt34TtgZZhb6hWtEQcKayD4i7jomHq
PkBlnRly7Pj0Hl99fnI9Bv7/ZRw1kOEKF/85dRIMPXkuDjiWpLb8gY9EahMy2Wm40wFn+2Vi1ZfL
4tYUaGmCWsk0EkYaHxtXY15N0PMScUKt9vPnrATo5UadzFo5u1UwiRiqMW47lVhqQ3buH0X91wJ3
4IqlBMhuLF1l3dM7VoUhR7S+N2SQ7EavFG+2WeSDn7gRxBC6JbFg46wcnNZesKtmN+fyMrTCLBpv
f3ki1nJR5kJiI/rwTMSAs8R4sKKFAdX2MztnHHu7fseymInz9HSEvt+l7+cN1pFy/FapgHbeIsVk
bEbfv6K3W5q0SNiMXANlWNyAb5PG/mScFgzXC+pKu1h/OFquWWHfFpSESDx0/pnUp5Z3KjNuHLDA
fbG7M4Qk6VMrLtuMtaSyDY9QvZdtQ/og0GU01IxOPx07itc2pXHIx13bdReO1Ui6akNzPjk+2Llk
QOT1cvO3FBgs109PtUPOp+kV8BJ5TQTAAGo4Uqbgz3DDR2sYNXPhhzcqGMyOL2nJ9Tf15E+YyxG9
cl9A90AUW17ZyG3GIfp2lqFwsXUpZY/v75itrZ5w0pivkA/YE1scMMM1TFheezgOBrGXmsVSnzxc
ZJ/Z/+OtUmLUfF5G/CIL0baj80zukmr++MKvumwJfgJGh9BT0etbgCqH5T14XxWr5jWdurZBpLCg
aKOEdCcoBuLio0fkyrnjDbprKuCaefbF7ZuB31tRqEuZa1Tz26/lsjWoEYnzS5LkICqloPB2sOMx
yHfBu8ee67xYWVhu9DAnjhhjeHaIPd7XaT+OTMMoWT5YXUhmZfEG1RnYuE4wy+3CE2eRxn00ECjC
LCXNqdotbKYhbLc/gQvetIJG30q1wgzSUNZQ9ozAuh0qLI0U0MadXJGoNwV5rDUIIqXNkw26QbdG
GwBCFhfP8ffuN5aY834pGiWuTYtLcY2QriiCrwwFO5eU1S24piSymOD5D6RLwWmx66LopKgaXHf3
IeCePgbGkGYTphMKwwmKAMD7RrLS3Q+8MGrzcG5QMklaobzr1vyDqcVvIkacvQvCzpENMX4Soo9+
1MsCn4BrYesVt7fw1+WmNayUyOE8UwvfogOb2+9EfkfLnPtr+E61lZIjA2qIGMQs5mhO0Sln+Q4M
+uJIQHPtSwS0ZbgntEiH4Ndt7hVjG8MF4pJnyAVucWCdO0Euq7mFbK4CHLRqUGMCzbzK0E+qN+0l
CMGTrqFY1FfKigWSi35sdGwRmchjiFMCdwBjRNNY+UzjMmXOFL0cTWBToQKimuYjNWSWZ+HjMDU6
7qagUsOq2yxTNeCuS4Pz0yJKSrYpkjXU52TzA3AE/bXkYLeY5uHw579ObhP/y6nMd3OTblni7y9v
YnT/OT3WUAglpeynXQI8pLr312V5eqaTKf+2HWlTxgkfuhECTZEKSIOMfnYpIFjjVx99uznmWAeg
TK2BMb5ZESC0WAF7pqD7DvzVJ0XdeRZl9/Bl8Ksi+yhowxxiBcNheEny0h2lnCcVkOYPGhuu5bc0
OVF48MHR0ZpJ2IM35XqDxIkWZTicQMbnRWiKbn5zTDGnIzl1EGi120kbnqA3O+dcQORhefDsGhvm
aZJap0Ev9mXuIN1kjZTIsBzJwMtP87pN1dpF5SKH5+6Zig9Ymr8wSjVK0nYirNkpJm9o4VrC0PhV
zONfP8mi4WvGIqR36zUqyOEVRD59nZhRSLUB+bHbf0qgfpEM9miynX3Wvt+Xst1PRMOV6Kv4TXNB
41kkEk+/6EV97MYNT24ieGanSUxiN9x83kTb3ID+0dW8ig2yPYmBqlkUmtoIvwAT3YakWdDQnw62
H84AddKSz3kztHtuyHLUR3eqqZ5x5kQYw8XODZhgRBU2x/Qt1lupycLsBx6mylmPqhV7rpgKlPdx
z9LUgIbMu/73cc91ON1JklJxPkSL4pl1R6KqhS11KaKlnXtjReQ2qAs7h68XDsUUJML1HyhP4DC4
hEBapoOGsI05c05f4X25N6jQvXlvt1TjvTp6To9nDzj6ko0Z5G9CkagFjnGFCtVWkUEZrKHkCbSN
7reLxQqqEQhnaYXjO5+QMZsGZumhYsSwVZQT3vGFjL2Ue1pQAgVLfUk3u8c9YiAM3g3Dmt7XodGp
pCluZY2SR1jAOaYISakp6OXOS6KIGhTeINpxAdirPQ9w1diWyi8uO1nDudag48NmLtFhIcWzCRZR
rwFTf2GXc+sktDC3qQtDptkVW7Jj+Ymuip8TX2cs4wCnsvxyN8/dWnb0Wc0Wzwx/ifyOxAMrYdbm
V2IE/5YzSDnvCPiifdmboeMOJsFzxpSzL39Iixjt76eU43lnggENB8gs6RJoxENe/xRjuCkUgmsW
jeTvKZo3dzV//aHH4v6H8Q17geF5gMynCeWmNPvsT+i9EI1+ADRXm77+7qojMnpTOOhSnacbR3tC
ut7cIAQnUITGEXZ+L6nXymeqnqce+gvTsbdnYrnOByx17de3MoUaxO0Y9toz3ghdnmFRcUG2z5MZ
/PuIX0oG1xLTLIu0XB/WvEZrrFEfeSM3BvvyM7yeIfwa+3kOQE+anWGxO/Cls/g1UfvHHlO7ucrX
5p6KWIEno71Z7JsLxBOAoynerzeM5ADSMemPk1fn/A3AUif5obBR/Ueh9F7ACUeHXGSDtujEyrzq
hg2ezY76AtcGVr6FHSaustRoxcHAGwBQVavz+BvekjgUKMBtk1nefGJCpg7pxBzxWGFPFYSsGnfn
HnmsamvfpMioxfFvcbRTmQaylJ0z6RInOnYYXJjpjXE5kwl/Ds5JaeCoRkN6FDTVapJX7sg+f186
MJawz1CyvVAOc4eMyYCmlhPO6gvh2aHk3A+TqTI7UXCnQrYi/Eh3QDfJTektbPlcd0+VLVg0iC/y
1DoPSGNclN/iVxATTidk3ovsdlu/FUn+rhLkN0HSEff8zZQFTgsqGagiS6l7L3BWbDM2L3dV3ms/
+0y+hI1dq7J5FDeqKymIELdsV7sSYGS20UhvIGForm0SNeG6JhUVA1l0Xk+nnJJpCXQpngbnOxRD
w3+/cT9/Pwk+5X0bWT+z7TnrsHuwxHw32gD7y56vCNvrZRI8+xfc/DchFtMDkK+nPxcWscRqUoPn
7nQm7Eyw3yvjf8T7qi71+eDZFXkFQ0WqYaduHXq3liiAYhslaFxw2a8ZW7oJNGIS9INv2meD4Ohn
cQLXhultcsgpEj65tjIrEHayLwxRXFjuRExFo0dIMfdx7fAY3i+XYNv9Lo6ruNFz29xoz5K4kGy4
5dy/d3YmfL4Pi/02h/JRd5z9MSww6l+ng0jjxazpfrw0to0TQTHI0ccS4Zpb0FA3G6hzi18Km9so
Wscl3+5A8xKhXxBgJbtSmJmHg3s581P2vX7gttYxM7d7LShbe9MigpYoWeSO4046WfA0cmjEJiRJ
oUPai98hgvXeL3+KaZprKLvfzxwDm2Y951xBse0Csp0EgyNs78DAAgME7emohqxWGzwYrlPPI2Xq
KL8OlWvqNEhLBv1KcNitf1m7FbdeMjfKKForlUuTz6iJV3jXqKiH9HV2rYdgdiuHoM6V/PgJjHcu
85hsk1s0kWLzAtoON8gDaHatWXglibR+8bmGlCcFdnmtCg9f0f9wfo/Jt/xU3ZpLbz/24Nt0CJvt
Vs/3B/0HouEAFxgp4pvYCbzfwHLyhokBAyYkTbIsX7hoDrhYR+NJB2lfFnQmn0K5IWhWjdoK8Ugz
QEqJq6MqJhe3PfvMopjIX8lxB0VF/AaHrQgg1eOc9qDZRYG2y2lfwsOO+jNgAcfICLBILavX/5j1
k5gFE9+2qgBtWQ4i8u1JkJB1QZY4J1WlxEeMTxr2lemiDuRtICLYgURmj/SPHflH59SoV7lz2U4S
6TSGAxkUL+5nbUB3GyiAxZGqxSkgbUTgQrZ7ANzQkEHJdS6cHdableT+33AfrlViXDkEjEJOLeka
+SKT1fyF7pILorZYP0dm0fO6EEi0P6PDmVFPDEZCUi/VsIUDohZEN0bFz8F5XYnjLEIYV/Ci0CjC
zuJJwsllL7CK60f9YyJQPknC6UCVpcG8gzsllwPQw4LH29VHpeFQUFjL3HTe95FUZxWLketIet+n
AFTAbXI6QVqEcZJLAOldfg4PnRVlOUJRhWRT+E5WTzBcT6s2r35jBuqwpnqXyU8dx4BuJ/FLgTaM
uR5huEpAu0+w8T+xo0pBKDwH98B+G200tOeGGmP8kz0yiJLwEM0Clu9hT34qGrStVRDCQyJDKXmk
bkcAOwfL2P9DiemgZSCGTTw1Iij45RwumgGa5/46TE3R+ZQNupz0BfBOZWzCjC4Y7Qt7LJP6s1+v
SJ2hb65w0aSzaH3oAPlx5no2IPOsuRGl6zkbz1Z312Ag5yaPBcb8KkaMbDZSHtUGFzRnBKpqiHwv
1BL32sL1Wusy+R7ogztwMMaPH1j+DNhmeY09uIV6CMwdwzH7M9k2GE4S3LEonX9CtrBaxqVh14QH
h7/bkKXjC+Vv4b3d4F72zvMBGpzL2//1BkYHtFjW8IPfnTkCzJOT2HuqDF/yjJNiL7VzRpdbmOAA
vvjzjhe7Y3ztBJZFnKddrsb3onPSodtCVJZjM9FvIizFAFXsijdccrC4eR0AGL2FyWvIphfr8aY2
aWZqL4cxEVFocV3AWuk8osMaWg318cZe5hejYj6wQfWrqwSjfvx8Ljo/+cVYIWD+rPMbLrgEuwSB
RHSkoPi3Pcflw0IkOrgdFQvR2LsXijassUOVU8/XVVvRofmiPPTV4eeYMZ1ld22s/SG5DGB0RLEL
DTyqlb77nMUhmKmoDkBbtDnMXXE4g/88yjAqA/rP5yH0NsBjER5yysCYLW68nzuzsibfNSK7120d
dQOWnKcakpoGvmmZwkD0k5Doqwni/dV5Lj6Kuf2GDaQXw36KniczKftAQLUew+UASb1o4yASBznx
Xvk8j1guBZwNtj4/m7gCdrqhoZlB8/Lf7r12uwsAPMsMq4S2VfD+Ha9mE4fiNQ69otWJjgpb3hnI
3hFBsX9c26tIfnEizahJVOuKlvKJNW8nXcOJNbGUx7R3oCPtnKPcEu8p46XggShzzjC2obFdQG1Q
/VGesMCv2WTVF/dquHPC1tDFUXPa/lcYvBWoMHsLrntEUArJQE51HcXFKNB6/ujeglYztuRlAVqC
Jzby/6gTdWZn/sh7Ifgks9ijDl/bq/hmrh1MwqCFEnwGxLlXnQOJMRnwty0T6syW6w+TS5vQaTpH
1ghKR/5rnAQ5pu/QeXibnA/nH2oJND0oXJ0JzZvzG2Hqo3iiEG5KUaU6TmPbUoxOH0FLoxR3LrAP
gSpa5TjX886L8dDBwpJofCwqMpwcOngubFXUhBLafk2RHhjnSZMXqA0LLHlkIoW/UrjIeCvOGFfX
NKI2Ax3dBJp4CdT4tNY9PZumCJEIHfiHj5fM8ImR8ZReJJKs4einXdeoarq7zTbaEJVluTVrqjPq
cXJ+Q+cTYl9P+Duq4c0pLvQY8osUK0KZvHmHoFmyguc1ArZ+4m4kcyyKUjyYPp81mHf8HbTkWzip
p4AzotlYkZM+HnIqskcOB9TT7ShuepN/jlcFBXJB5iKEfwi2OabqJdePH5EGITnE0+0JVawAodzW
KgBVNPR0p5/i3S8AYwNqnC587eZkUfNWR4iS/nGRyz+QGJ0VakTp43zAXrEESIMCy+rGqVJldwrB
ByUChvpSvwvURXM0+uCYsuCgrG+eD+/9la/KlS8U0Q05oWM5RzZu93iQt16eW+/I2+Tynq1Nr1uu
jU2A3u95nA7LAVPdALhCjJJL9IdpO/TfOgzfpRP9AvZPK9AyWWBSoc0UaCwoBJJDEoj7Jype1OkS
uHiWIZHJsHol9v/xUZTzWeWHqlxBNcaUwKCM9C0yCP8+fSri/UWnwi6Ji+Mg9V65JrbwhX/yT6EF
a4+FHL4rcVV4cKfTq2a2G51zHJnW4bu5kaO/gT6TNrJewyMoYidkOC1WIVjTId4uSrFC90pLbw67
uqejVGM4YDcMAW2yqcDIxpu25216RELn661PF2l2bQkNvXOjv+VHmjCp8fVUlwIa38v0KtxGYzyk
pQ/8jI9pAScf0gJwl3cEylBEp0nQRmXFTMkzHqwNtL/QMl11o+iJfIBYhMDZ04khJ9R0Dn1gRjjP
5Je4M0vVtYFdM2fFzX3T7mFXkM+K94wIxV/D8tvoFTWaGoUFA42x8gGkR76l2GUkvT3n8I5kYu18
zTNMpLw7LP8UYE+P4K9DVjiOCsRtl94vk1Xzkpag+MQTopJvAtns/H8OepMO4ULmsrr9M6PAECKf
bhjdA0FSgszOFHz4jCVGsvP+IfXLx7JVfoYBy3gEf7HDec1TcKB0bl2DnKod4AwbB0Xwbq2guiyz
nFbhFqC+WcFrMtSSU7jp/TDfugVyZTfcMp4FnVHEu7MNwz7KRoQXR6cAJ6iYgzgJRl4kWZBg9T0T
cxDtVoi4sT5dIzXw8zxPNNvpMr4uPLT1jfq2sJM8b9kF6YJYrbY0ZZzZo4dazhKDEOWjvQohzNNu
2ITBCt5SxETvnBn9/q7fiY1BE2Tsze1YkjFYUKHkTeKbli9zj7Htx/RFmxmcuaSv2thLtHUllfqK
R1YC2cVaIzImgLvxOtoP1Zb2of5DM73GlutglDmuDEBeBg5yI90qIfNzcDRv4lzzv2g27tqDNMWu
v6fxIH9hKFnSmZoGIOGfibX2473i7jGtNafuExWYKkWs1k6ui7qfnO0BW1Mk0Tb/nkshKeOhR5pR
UbZJ23hSKx00IHAtpnAiQEjm9sk/yjFWILsFKgYFGIO6Fw1EiPF/FrBGq383sjgmYgxuUILOfVJF
RKvEGxbgvawjYkgcO8Y9nZ8Gk0yk4c1xeUBsEQWZK6Z6YqK5RPef4yssWCakKWt61MoEO8Xj22jr
p2NFUNsQLOFnNF6IA4QmzOf0yYhqtXiqS/1ye/Oh2hj8jDAEJGbZqw9GAuKKrHkR142TKPFKjToA
SlweVGU0jdLeo4GR3C5W6HaGuGP0KzFQnvdxWebckg4yjFor36BVrPMb0VGe9Md7q15ACzjWnlX6
sK14UdoUabVQ0uU5klHYPzDUu8wAMLBVRJyI243oK0n0SphlTSOqTC4kaoftcbFYylVZHeLkC9Nh
JYOSdLJ7t4Fp74zpYnkApUTjXoMbEM6BFhe2vqEI7TL0DxWWyJAeZDy+GPz/A79F/4Kd6gaah9EB
gJVSzKbYhzU5soIin9fLSjfl00Mr0rr+gQ1ZTAxLltId7T9cu0iPsAc7dw+s7NTXpd59Z5pW1hhK
ddZJdp8SV40knom0fktCO+hjCsPNeBP3enyy8eVv1GDOWpEEmlqzW5ZrMCejuUbhWIxO7VStsS+A
jdNjJ1YjcXRr+iv8JTyce5HojtLY0v8eRR3M+xLwSNafnCd3AVCjipxw9Ogk/7WO3E+NoysvVy3l
p7cQ1M1Jr0WLdzYhRvfpHzY8bK8uqec4DZoPBf+5Gx4Nf2UzKYQNfgg3SK9Nw6ZgtJtpTSxCExjF
JremIZOrLTfGDZgQLs4cb1Zj4CwtLjDLXLehc7/Nb2Uqu5OHIRvCNHT3zMp7+BAgjgV2mVjxDfqU
PoRCTkdmlmhVEh/E2YLDoTRPsfoU0UUgkMtpm1ZfJNf1+WKVA8LP8SFMihDsrvOZ7Iv+1wdYMquG
c48BmNeHKhEcHNXHeKak7HHCEpJzvl/iaoJpTRi/g4hIzf14NJL7+ryw7NO0oIO8K4kom9cee9XR
DYjH+FdU2U09Bi9NKWnZsIK3KBLAkYXFkI0rRExzgnp1CPWzcrGAdgsqqcM3M9RzRoLtKFVXmBDP
ERlNPAyxukv3ru35xEPj9nwmYGyAll9L8yFy45JUxjq1T0BaDMew9cmMe4kxdH6EyhYo/qosNb3I
NlF478O04D6j3GgMHvsLnD3+gOEPMa+bcvi1MW3kA9x9TV4LWxhysn5hCl3jIfVfo15zt3szRxpU
EdM5e+m1zJbhpPmLRgTcJ2f+v2JAFCd1pWEzUzh9aNPnXCqYylmq2tBBdCJIz7DWcvGJChlf89KT
Q7kEx401oP2VgXA8iQmwsHDWePAK1TLozMLoQ2EL+O9zmyzCFujyaXrXbxs053EwSMVP9yZFyeou
s4egj1iwRRjeuBaN+Xa0M9yN9Ea6p1jIrcbjY8XLy7pCp2T25JBhPs56b0qcY0EnpqRzGQEuYsMC
GNsXwDI5MGbBNMGQflB0VMImx1zlcjHJR0wUabRoKLqsWtR7rhRuBvmEilCgusVdjiE1uaY9UtvV
zv29gy9nuUFkM/1c1TpSpiv3cAIOzhgwLHErC2KWutxsIRcWOXfzA6TASXIsV3Pm0GryLR2PARzX
z7RQQWCafsKDNVQOemnBHXloq/HLlKGyQjmrRNrS/04miqdHGORa5HjWbMyHpceov8PCii6vUJ0q
Jy9T+eGIufZrpyUxtRel3krbK1zrtZ+1vDly2QYgcirlmtVl9bns4QAj45/UdqfX0iUnd0wPJWTz
uEMtxhoXG7zM7vKf3l0+unfgEnjPGNl9KcldrYpdGQKKHQcYMQc0TuyHwfgWz9bHOvGlzcakxLzO
Y3e7DQauqxVDDSzJ3cA9+oEbYbs3viS3e3D+Qgj4whI4FbuK52JsrReGLbYj/cvaYwac+UeyIzDn
/IEn8cY2Pj8gIjKY6J7HfMQBvqZgkoBFUe+2Ifh4I5BM2kKdAHxaivDKAfBUbpDxhMmh5FiYfTwn
4k70eCAhAxDQ79xu4D/HMrTpa+YAx3qk9M2RdKMoJpwCUXLlyfCCcjXn0jn8556/oglf82qClwjb
9LDzXs8mN+2CYDqCTFYmEUMlQmRp/MQv/3H2lvPQ6E3fH8Pd0DmfPbVgdG7DyVXzSjHR3DiEj/Ga
kIK7ZFscH1fG21Q/8Ijwgv2yz0TRa74ist9+My1GjSW91M44GVbisQzLmsrLQAfFNLd8OMyGoPN2
Pbr55HsMPQix415gEgss2AT8WhkOjquaMEzr/47Dai0t4XJtX6iSEB9nMl6hvRBXl/UmJ8F42Ru6
uu9SqQsaU/zBOksEi0gh4swRFomXniwEkCux0MztvsIcoYKFsNbxCymSMNnrvwFN/DlaQMBES386
ff6Qr96Rh/XAukuVQsB/00Bgg5z+Z54AueJFaCkFb0gDSfQCvsO4nZpl0T7c0owZx9KBefUId1yF
bDksaj8gYbLgVL+mvKjsYNMkqTQXK7GLwVxZpZEuE8BZkhB5sRFc3JuSSe07sagXM8/zWMJwQ5Ud
Wf2f7QW14oX0CH2OmZrSVFi2/dHTz0thbsYjaNYka0WW+gFSN1Lgp16+GzoxIJNj59xL5Hixo9wn
Lg2cXqsq3dg37KKHHqbbvMEQKqHzyIh0E4RLt6RItrFVh8YvLnLhqILkurfJa1X+viMbOtVg9Dk3
0OW4gNgwfrEETy/HcfTF8rwO1HBtkxhX+Ti14trtwu+HNBjR+Scbe0J2VORA1bgPGeNpDFcIw3oK
eDxwsHu/dnFvMRWmmAWhwl5NE+0nE5FxlOdVgch4igf1jG/kvGk7UnVwI4hJ5rOEsTr5sfZqYMYr
NVSIlNz1QEYs1Oxqxc/zF0g04PKT0H7PN7k9AKueUVr0vLoeZoxmAjYbRDO0FIXKiawUrqn7OSBZ
d0aGldQffP5yWc6oRS2I/dtsbC+EjLL7TqIw9KCnpaRQJLhph8FKj7puBWakN7B+vCKfZryyjk3x
ZU4514V72WpqXuevruthDpS20WCO7fYKrz9BZ11b2nKvBodvsgOTcYrdecE0gMpVrst0N+oA4v8V
APjFQzR09S3yAjA8yf885X4x3n3ptNRIxwKAc0QVRlJe6Ow+0hNNOfX71EyeZidnd3l7KomqRcnO
e++bptOQjs4neI7aTrBHXbfSAFXPL/JtK5rOQZeZGyJeGTXGtpZz3bQRfMpvFfmLpvwToadlnXJl
TeehR+5YuD3A+j+qYfYtsPTa7IpnbtGAEvaMLo9ZVpkcQCVQsIXHqnhcrJV+OCaWf4PqTdrBO7TG
VLc5praie7koJl0h6FjmCJ62Iecq++tru7Hwc4dkiuEA66YTeumuVHPVvg2Z74oR0jegbgfkPrT/
+//ET7m7HGCMBIIRfPpBPRszfJT1cmfrzGzX7lu7BbIMDFyE+YKT3VRPNqDS5iUpsgH+icLjECrv
JO9dECeTr3h2ROla75UUn5P1hahlAkonu3Og8ICgAtPtSyqQOSYbZirKpxR8QZIOlHTfgXXd8RLt
oUnaanZM34ejLWt3iuM9bCNN3yrmQzw4iveSP2EyrcBXpOR0mHCJn6pT2+shTJW9mOD3s+4dNr6R
98kb7QREy+y2HH28jOI2LzWJJNvBhOSladT1VEtcpFIZYdtKji3THqSLkjpDfojjSwlhNR5FCM5L
C4etd0YLZIFGLKEDSgDaxt/yY94UdsvS5R4VdNaZp/FT5UPL4wx9OPiJ8YYoGhBn0uA1gz+IPg6F
N2TmEBKtVYR62hMPVDkRFj7YRS447amhEMPNkrgSDJyNyvBXwiMnnRH+JTR0sIuzNMe6Ph0sYqBv
FuP4E3uOBeUjWfaZ28OMnzebITkY0+GpEhO3NqSDWVVFxNogZ+D6hRA+tTkKCTpuqz/3js5pvJ+u
d3uduop7c71LIDEvC69h9k/t2iulfSXsh7CpsrNwfHxOFIB/phbMzUzX+S/yWqR6vCyNe8IB0CzJ
eMsmfbp8QRkrA4BA2+s7RdoSm/gfV0eTWbsW28ZF0aJTlDH6nbAfCYF5JFpsq4o/jU1+F5J+a9Z0
ge55RkFwN1E4mYVxW6yODq6fdNN688ulCcupEP+d4Q+GtVj09w12Wq9GWMbmYX8D6HAu762xpRd+
J0wHEUEwNU0g5wwVy44U/q8nG4SjjuxJcWIQwrVi3D6MMaT28tBPUYimsgD30U4R1soCorQ6uPLm
Zqgm0l3xO3aVWpqGo7m4lXKGAW3yWx3s/TA7LDfVZxN3R7+TkOcKBwc6ruNY4uhUpbBVeixyvPm4
SNK433cqrcOU2f5nNh9luaQs2ZEVz9/Z4LhW2U++pFjlLcc/2/0WZw+jMpf3BgU08mry+PnlsoT8
vIfAC0F5NPXU5oER/XIL0F2bb9R3wocqcjE+dYfsboLLBBZtkvGgbtmzdgU/+Q8Ti5cQFBT85L0e
Mgff1WnoS+UgezlL4JOjRhmO25HSssg5Ofhjnh5JvPDH62D0wHeA+Mz0+GCizy5u2SlBgYBsnaar
IGeZkMszQKN7inCqNELz+v+9FfLY+stOoaoFq9jFNVilyHaulTtJ9x22buB7RE3un18X3MXNAl/M
g3ME+KDQnYAAeVHouP4J8t2iMLOZ5JmHvi/9WbHPBZO98GEf0VpwrIGc6RQ262t00J15LMipzi+t
9Rh5hmat6xbcYr/Bu1Wqmy0++BisziZ4mlMaSMztK8NxHv1tqivP0p60xlYvjQsGdguFN/0lMILW
+FXksbu50inb4eQ7gsE2qrAPfN0A9YY+cTWyCnpD+RFI97lwGFS3gF4s2XlhByP3ldWGp8GcfBq+
/qtjBtMnl1vt7v7eud0OYE4BVLi9+fUZngiEkiXFmtUR1rtjb2/53K8/2UIynitGWfCu6Wqpvv7m
u0mBx8TmEeuq9mSc3/YS9AOKny8ZwBDINB0T2quyusgHCUs58Fb5vyKN+3srvVftVUVm501ZfDp4
ONsYI5ojUABSJ0PyY9S+ICt0otXYPhFR+UlXqcot5ssC9t8xQMcAzVot3akxR/YOdu+0+MHC/vRh
BfjmsVcF7I+3CRqpsP4L6JpItrFkmIkMPvZvbqBr4A0RYLgrdopt53nTlgUK6CoYa6aWlirz/hOC
3ruEHCAi8zaF9NkkAdPczNeGqfaKixQ8WoOPe6wZqsplRVG+PpCW8WHwFPCuRSyAY1AuG83paUtQ
tbMeFcf00vPXSpE/qDV1mnZgc2WvefCAEg2p1JQxkjwTMzuHMYFPcrWSgzYGGOwPZcUaDKAkkT+2
grsAd5L1q/rRGwBkOX9267/4ye3K/lHHLm6FeGp4nurxutoYzjD3sploiomrnYCxa1D5OhHCrtOy
TtPvNJNoyAQlv77t54gUobWanYGvTwFSNCXgtqNuWfIAiIzhs4NsJ+ryBHJFa8aC8crFu47O5Jjq
VnCkbIfO/TjQFQ71kq57K0wKlnKRndWGcGM8zW6oPSCHiJmH7S44pXVXA4jn/Ptqk9tZ3i55HZkD
u17Vxm/Ff5mWBOa5TG4ga33FDOUnkvfyoPEJfiU3PBAL+2jV5zUuwJTHUbsYGtN7Inu+Y+UDRkvs
SHYY/lErJg0HTCcVyn1eC223ELt1gfKrrbIF0t+Awt02RFS3n1DMO1vYdmWyjjyjq3jeq3hbTdvn
BkEa3iWFZ+Xbp2pxst++AdUhu54Jnyr8kP/Fwg/U2LedLo1oSGGC+xfqXPTX8QimrAh48cNMPPTz
I9ccNbZ75+07T8eAUuMy8SSA6N17NgIC/eJ7FC3KGpuISBZF2tm/jD8Sqja3RjlpZdlmH+ShndGC
i19rD1EtQ0t5vggxUczLV2EGCiQVg414kt0SjHVGNjh2bcxKSr+kpr2UO6lrM0MI3FS/5yNECy3r
pKSVacoProMzU1m0EqS6RONIAIVhGYoyGL0vGhIqLwzfFV8sNcbso4/dwBSUa5R6zbZkKwPHVjWp
jwqlB+uukxIkebTxil2izN9YSSe9B+/CNVVak0FepsFFssCMTUP5OeQpPZ9SSaEC11djbJvcleW2
WarXo5lB9sYbYtKx4inwaQsPKZVAIH/t/1C34Ws/jDIf8UKorqWe4dV9ocbFUhEOmZdrUlHL5tb+
QBt1NdwtMQ0K/kRBCaWzQ9sHdGJr81egdxg9rTDi3Ts40RtND31kLqW6wKosZwHXET4TRi4UzQi3
Tn1rqgyEPxIYjNA6NWRTMCNBViMxRHzCe5K+wB7+xkJeGB3FMGS5rxez8ZUuskfnig7CBRQ/WjYz
978TRDOmsHsmj+djqltQWfpVacAywvpsc8EwmsSA/ByiWQ4Q1Om53yO0rAPxoV0EZAXnmVnX5lT9
zPpbVDtMGSZJq1We0MYNtMliGIAoFjf76Rz7rutfQJGgC5UQn0X6ClPBBvhRO0HGk8/0Orj0YncG
ClKFdij1zvuiNP/PbpN2/+PxPb/1jETsxZnsjxwUQOV+LoJxw2lF7eFH8NS8x2/s099Q+4gYcVgX
Xm5gJJCkIOh7XXaS54iA4Pkx5f8aUuOsy6n61YC2mTBZbzI+uqoCKrpZHjSShowc4MHmgE+7XUXF
bLeIqkEOwc9A8kKHhZNQJmyKPK8lARKBKNghn1g97Zsdt5PpZDC1bC48VLdV/g2fPM+UAalw9KKI
x50ylenfaLpQFL7n2cBce0xabp3w3iyRiAWDEI6dRnAVCFQinb6xVFE1FTR9uBw8DCZTdg2agGN+
1J1cUH+We0/QAYeRFOc29hUswhM6RnrTKEpdht6nQYOgpUSRtFFpyLJx+K+sTXHHC1BhLBY7nWty
FQOsYqQU5O33MjAaqDQQ4kWAuw57XTxO7XGMUjMKK4sSz1tiLeqV1U1k55QnJHGEhvhTd7WYIsF9
ryrkFaVMoipu9F8uRxqlcbJ0WfAFx10IF4Nhbb8zAa/UjCLAesgRJBeH9jiAIuLbu7iZBCZCJLXP
6fCMEwYOSqWzErg9dpJcaUcKYdIuoY+9l7WWssMnV4+QDjBpJOgWZp4ObQg8mJWrx26UCz0hay3m
R1qSVEkDQ5DnAWwzEBA90JiwQ4UA6wsCLQzBLoPdEbwF3b4+a1lnHIcAbgtj4cd3X3D01k5THBeK
iMDC8c/1Mja2WimmN6LW0S+9rZSzaeaKTPijbQMPdbmQvPyNJRVkJ8cG+XtDRdku2r7RoIVbZG8Z
Ur72FTGGTTxJ30lo+ZgkpnKv9Gw23e30mGco5CLwL0/M0vdMKL6tPEV2CARhvseqLPwxGkR+HcMD
pCMEmSdR036pNGji3A/zkNw8BrH76AwdaBMXED3AeQWWkibjXkLxeoGrcAvZfVY2khNQv1ivfZg9
6VjnGSaeT1uCeelz6aowQyPCzp+tACVUObni/+gYZBw/UBS1jPZ8Ph6TU/faNHlx+erpq1wsa+Wh
CvumT3kwyQRYzqlNWg7s9E7c0mH31UFLeryOM6E/jxmOXwZzUGULhQXfzCuUUhvpeCOXY2okF0JV
anryThuVAZ0VIS/NdgNUiDUYDGProkUuRcb0KrW3lfGNbkXRdjYxGBntuxve4Wzvny2oEIzKFHxM
J6mvebW2zq3mZ9yEtcrnaAr2Re2oIgmIltStBpCEP07AztbKdf6My5iy999MifirChulMl94b+RC
IonIkGMfkhaL6/eqO6aTjp4CJjEjUclAvxtXzfQJtq3+oO8p8INuGsVw2+mo9Ugx4EWdPxU3TYHp
Vq4RrGFfN0nxHgGZK0VKMGGY4lrtgm7TCtBkC5pXWVnnKU5w7+5SVn/SQj59/LCSdpzCPvP1DNTv
ZUItDGxMZ/BhBgNmjw0WjMhML9rqZxO2SoakqCrxqNKCazpfvwaMBCNnCmuIF5OfrVt77PdTxH6H
CfUDnJNn7OfBqvNlt9GMyn4EHtLZP572zUHXXBYTNT9D1K8wXR1mbX1SmoB+so5YuTNtRaaCdrzC
JKB2HmJzaw/kfJcCmoZvE3UDHlIADVw9GspCbmYQjQPES6gF1J1tfMuhTelxBADZL6NA0vsMIBIQ
yUd5dmDm53mZ5qoKx5nZR24IgCwZHwQE7g4roy0f7k6aAqZusXo7OsE0FkcbkLwflav04odKP1B6
tF8xOr/MluhC2g0FW+nageEE7Y9qB13ZKjgzpCLk5d7h4uvmWWJJxCfZYQheseuVDKLU+HoHZ1CP
HwKzKt3h41Cy0CmAdxDedg7XJv4E8dcWCvBBqxWqe9fG0gueRDkWVRg37CWpPtEgFRJv+xYSFjlV
RHheQgAvppqGVIEWgwqAgOhQgCfYUw2uNPSnHMy+L93igyqLjH+Ry35oDleR5DHrQsNpO6RcDiGX
srzuF5eWpMqTuWduYOBZpjzh5FjTJ9FQvLnzAlxA9WPz6irNFvLkHlPBSDWxdnmH9VTauGHrwxM+
gT6zaM/ocYMEShlZ4X5KrAV01zC+h1XY+gFk4G6hpq8nXqlDFe9Kd8DOBxoluI0twHTKxqlwsko7
OBmXk3MiS1ugrEMqH03H44v2XgcXfzC6V8BFCMlhGgMXgKGB7QpdotqahnwHNa3AXG6A1JMncxfg
F8syZfIQOnv7I080nJk5pLAoS3jiyxD+G8iTWXPwZsZnN3blEPEemprsYHe4r45y8Dn8kLJKw+4A
BIw3WYQVY/kYX5gdtTuYf1+kQoXOtqojMMEMDxGwbjLDGEYhb4ZJAUX1v8NwcZz3HofO++oStMGN
qRsZowHpV1WgHenQOJwj2DvgOuxkaB5N6DpRqSAKC7JlamX3rh0dbioPS432FE9p/0K5Fo6JVCUd
oE3SSOsLxZ3e1sFxD+rcRibkCUz2fwls84OYF9GqWqtcJkXBfY645KKc06rOZqr1XeyLNUu59kq+
Gm5+dCSPCQSS/yqjfqqTkxjBwD/MZot/GuWjtf5fwarEqmBubvSUD1tyUhz/QvaosXAKFYlYwysw
jkfW52RTLxLv0tK6711IDOut9+xJE8prLD35bugvV9X2WR9NRQsjd+lC9YGG3hDC6qXeOhwmF8ZY
k/xVQDKXV3MgPLzDj6KyMWEyA2tBGErGezbUnYYoTqOkME29Xz+068zDQgeD3veg0/mGGysXeMd5
9TYMFnWTHPLlYaai+ePQJtlHUej/MTqoaLyM8w/7EcS+ytWlqsacTWm6DIGHGj3qSORxYhklVzrN
8CdimdSzZJktvPwBCnhI88Y22t+fmHWzcMfvI4xKrPTHsXO/ON0FNIRTdCJthsqxhE/0fnmxZ6Q3
RxZjwbWCmYFsG0jlow/7nDA4V9g1qaiGBOwhQN1JBUkWiKdjK4jzAV+CWaDUIxzQnTp+hn9kCXbf
xpH8Da6u8+Q2fo1cNH35aLurFJuczm1GPavtsHveFKJ1y1F6nRGbAmYaHVw5STehooIiZV05JwN8
VR2A0iLh2+45gs9Iw94lTZE2CnEJ5PEjIGyA9S4r0aIYeH+HxuoNesOy50BS4FvBP4wstyYi2rPW
VUvGHpeHfQXQHZpQE7ZuZp4usZp8+bXBqKCUl1psks997rNpf6rJOTu20v+RtSMrIYVLDQmYfxU8
317A6j2DAP4nEyxeZt140hnphaKTSibq0FTGZsrR2sGdrd9zilnwlXsA1BSAzkXRB7P9tz80G6uw
vVi3u6OL8cycOb8duEcZSwKH3za4mCD02SB8hNkXHcOsw8Z1CwHh2GMQL6yK2j7CHVdIV8WJ+MQA
bLCaMzaY2k2V52BcrxQqKEabuMDRg7RpD2dO+9y9WUOHxD5M+JRljzq0v+8JlBhlc5k+BrnsUulN
CdpVS3GNDaER8y1lmMffzZgXf97oyFwA6Wl0Pt8qR4Z46h08IvMhzVx4pvpSZ+/SRLHUHS0BEIpO
16V+IkGYlGGus7IiCMnLrxXAbgP2R6kJVMEhH7hfqWukpHumBz8K8CpcQbl+as5tUF9pSiqjtjJy
3HZsIKKQ7rN9tgXzbeYI+fNljXf2e+iwLRVzF5RyGCBDlvhcG0WvwKLkIu5lD/CAvdA2vlW4Gqgv
9lST83DgyYimEOkE6liT7S0Zsogg/lqay5nQi9mZczARn4jAMv07jIzyAwUtggv/1ONENppWWjeb
SjmDFs4EG0Afiw1V5yWd4PxcqNSKafFkV0b+OAfYvd+uuIiRcm2lCZaEkW7wfLz5w+R2l91UmkUK
Gl9NaUd1xwKNOZYgnLMis10V1gtSgxhbBrqMsXyXTbz5tM8XFYhklr30QVfug5w1JMTBWFJbNiV6
k1jbZvxoxktw+Ywq0Hhlu3nHNGpFGamNTA9EVkqYHYFLICVvFM+6VJ7N+fx117cZzpcmVPFyVdch
yNSdKenG+3gpL5pzgKyyVjVJ2yasC3fPHpRVJEoRA15C9mut7k2hTJAV1dH0Dsu9RFhXkFK6/Ln/
HFZ0o8zfT8VFnp0EdreFtI9CL7z4+c0OdstfOQc/UQuAYyXe/rgk7nKqbhsovwBBlFUHG3kMoo9B
w6HyT7UOpHuK2Vev4kA1eNWkMshxH7nAfF7otFllxuwQ8PNtrwsybgvV4oPK4s/cibwGsHZgrsfF
ZWorPfoDRiccYY7viE0QLc+PGqMFN5qqfbr50D7dX+fmN3lhY6wEb/zGxQbAV8RstR2keQhqmkLd
hGMZOEkMi1KXcYPH+DWoLbTwv3YY9kjq2W+mNvS7B0AfZa9A2dL3PH3eAe/TxOfS9xJK7Qjbld6y
45J9N43yhPxCvlIOAW553bTRv+B/LVaRZSfKn5jseGqlXWywzRwWklAzZ9k2tNbAO3t95ffwPSQb
Z5edQTjCYkpvQhHpK6Fx2oQX9GQcK2kcMELkW1AelKHpnyw+ixuTOQXKTLcmEdfcR+9YAjOp8hbU
dZ76CMzITOw6nmbwulZVsrBcfr+orn1UvJFKuFLBpZUyUuxcwLEBAAd0YsbGn4bxdj/9flKiI+2N
/TkoEVbdNZl/vwLLxosUf+4kABfbf64ylOmqdjemyaLHRnbC8pyy+gT0F7AO8prm/hHp3fkJjGnS
PBunvsI6jE/yZuDM+/CZhbg/TmHj3r22xy49H7mO62XlPckCtlTT9WDz3x6oUzAUawkRV2pRoBoK
lnudFLLPliiag1weyfz3OYAK9PKJ3BKdzsrSvYsrjglMz7dR6HPL3WX+enEPTYhwXLhQVbkChrZp
U/mRrVB5BY579mS8c0U8OGbWeIKKDxyGRoo2h3gUK+uhbQ3WgWMDLLsFE2mDq27i4sOEIkhnFC/m
MiSGXzU5/r4qCiVXSB35Eo3SBRK5O8ABnLjLorxl/syV5jWN721M77HhPFz8cDf4cywcT7dpkpya
NOh0uQMiA1aab0Z4k9Sc70oY0LE/DutzP6/Kzp/4w5gqMPGzKEcSUZWs+6UPH8Vfge353jDicjQ5
wUTInSlwMQKRAnKCiw/GlXcCayybG1KeHbOcM0Q+Yr2o5IKGK9mvZuaWlL/0BXK4YMpO22LtxSi3
K8dmMibOBnpuT0SzdiorwYtzwIR3NO6R3K+RXPvBG4otSLwM34Kq9DLi/Ojzmhnux5vpvNAnoQx4
cg9CLnRthTwGRaPCWvuGcgU4gGI7ja0x0XkOvbSXQ9DpMt0Y+RcjM8NKYeu+tfNODOvjel05hvu+
GQYr27OAOGz2gG9VW9EmrNys6kpHoRHIgEyZ6els6Ak1eL+1rb/9ePLwDkWEGQGvGPjNu8yFNOYv
k2scvDXa4uufgH3CsnyD5Eof4tSAC1yTZb7No2JnPgh5OSj9OSrhDPfzBWu2RMvTC/zQQnJjDKP+
i9vkisyWq8MEaxGWA7oThzLR+0t+j58tHfGKBbbXSRr5PtgEsjqjNnE/b43VDqzDgeEAexWbj/q3
X7O4+8nFTuvaQCgJKsYzycFU+UMUWKEhlMPWa3GcOcc4vPUquCu9tgMnmZn1JgdZil+i8bHZ0EfU
dY4fwDe7zQU9UhdGcGe8EEMwMUKycKLfBkwEqJzgGAVc3jOcSJyyCuujPMV1bQpqW73VAcvCbfbc
xF7VC/osj3lBGh0wVOKK94O5uTN0b3+fJNquDFl7Mv4n10nBIjnNJba6fETuTZlyJMVJyu6yWEUm
xlnICop89otqw0adF80Be0uVtonHoQApfV8Bk99mmUNdd81D2tjatlLFz8U5lQ3gO0Z+/RWF+hyp
AFMh4uthwLdibkIg+4J68wkfzdHml1OMpZSRG0AKCvt+QXzlk4OxeGemBV728eZb+y1fH3ukwzME
KpDRnif04ei3xkXaJFQyKjVU48atlF1UR0pYacCDzHRUQnpB7rJFhcdkvrYUwG162Ro/KEBQuFG9
ba4ALlqGatHwMGtlCqK2Z33Y6FNzvXw3fN1gZtcoYcz+tw9AqSdqzZTvRjqJkUt6TLtcFLywbA6G
B5xRWpiAEbB0HJyfDtlP4EtPIws36X18hLJlz9FcZiZZnbKByK2nkxO7bfZnMzEWfUqDTDF3e0d9
ZsyG0NlojN66ERwmDBLEIeWeKuK8RpsSBWMLn2dPyuXz2cihaB9vfhB/6/epqSEFu9qnZa2yUSyo
2eoIleKt4otMv+GNfHlVjy1v425UKUysscdT5ovxReiHYXAdMzbudcOxf5Uw4tLmPXm1B5CndpkN
TtcoM6ZQvOPf1q8/7ka+alJXptFqkQpI2ILKjcGDCfqcWy08NERh0pZR5s4UDHZ76gxwMCqa6r3c
ywkXteBxYIT5bkqcE+iLlaIBsGD8erBSHyXXWPWztazox6SXFR4aGfKPLi6RNpElnvKiPZau2kr0
8soLpuxuDA6Z8EWx8XyunY+Aphbl+cppTe/5Xju0vldJBlWPT0Ef6SK76A1uqVB1zUVZD/IFGKKT
cYePVmwbMTshLiw+f7KfhsaZNHmMqG9bY4ghUXcQI2btw6+kq7q6MwtD+yzYQbbKMPGcrvWpPdHW
EQQ3UrxMH/ilF8YZL/yWFJCo28LESSEcmInMLLl8+OWYq4BuZUMcNKCTok+2d1OJc97uKIy8O4bv
4rzbOlvwTqjMOO2H7E5DyYQaUyE435jON7t0VytHx+qA1Hu8gMSJr1fU67sqHMyVuGW4N2LoSSpH
pm3lQnIweyq+30OgjNorY7hWGIVsqvDw5CsCFz9yvmeHlcNnk+o6tdmzK9sL30vyIpEsJN0e+1Wy
nzqUx2qriN+9ZS9Letd9kERZ+0wFfCN16Boe1TEWGl5GCJLvcKYFvMhtoG/7CHDA0SyVP3iX59Tx
pjUlNC9pva/cvezIdT8Bo1cT7ZCS3v7EmKa7IZaK8idpCISXWvYyVMm4nbg9/wtLcd0mVP51pTpl
KZkXA32tkrHjGvWHEe3kVR1KI8eYoB9j8BYkDulP7G+3AYt6cSlzjSoSgHXh1s0HCT4ggO1zuXC7
2K7fDsVYhcy22pOF1McmrogEWDOWj4KAU8pPoSqwSAMZUTZaT/le8Zy0/CGGno9hNe++IEyT2vuJ
EttDRrExEsS9jcXuDXkKhYvNuuNnPhzfNOLxORluDAA41KmMCNd5W7VO40ZxFpHT4UJEeZzNq/Q4
VPRKyQucQ2Anupfm6M9SF9nP008AgJwD0QwS4xnwqrmIFw+/WM3Jot7ZUEo89eNFFHnAsUISSz9R
7s2PInAqaS39k9M0yl9eCmaleLvWFUStlRrSZMml2o4sGp4aM48Dh1xR1hrF5KuMErdA6G9Yw+4v
2/xqig6HbePyhtsSLqf/jg/dcbzUL6nMUTO/xiNQrlA+cdD0OpYP/bze6q2dpeDf3E8XJt2U0aX+
2OMXnrfZWAS4j5IGbWuFtYZ0rAGXtv4gjhBHfBec1q+3l7XxePfPU7g7HApnUd9L3rpm38D1Jq/i
KlaRLwvmeJfNa7v3O1yFNWHu/b4cig5LfhNjNB4YAgg2j5zXhJsAwwE/cUQZZpdWExOZwBYE6O+O
+SilucMUs7mRNX/wVWzJO9BSWx+fhr9E281ts1HMp2LXWfan3fpheFUGz7qFMLJAUmgrwmn0GRjW
fBFnNoXEySx6iR2DYQET+ov370iW94FmdxPDSCESGtXF052USG1NnuqcqT3yYkY83MSjw2r1cC3g
UqZ7b1kdMwmDtW9LAWF7kuK3Y7JJ8pPDQETbJKACPBTKQ5A0o76pLLhytYl4fFOJ300ip8PAIL9L
uDwCulw3NSjkRtfErwoc8Cd73gT1skcWe+3uRnsgScQjxpY6Hx0sWsY62bbM47yXKakeE8mlV3Ud
URTOCATjtXkOP5IGKF1luj6F+3ON0RyD14CtGbw/7S9ZJ3HryskB1j/9cNVWaRnroZ4u0Tk7q6xH
7e7wYa0aIyeayfqaJVeEIcy6Nkt10Enbmith1nr5/6DMwOPsoK5y1XIaDd51BQSh6Nw7oxs5AAM5
T0WJLnoOlT4vwhVC5HdjuFIMOAyQ1zq47qfgMLf/OD8sK+c8s31eEhZe5uWq/phmY4DJdsJMYdXO
3Xn6Og/T/+ztQV7NvvuGcQEwb/jA4Leaq0BCkjSpw2FeBSbfH4n7JyceBtgxOzkXsLDE4MUFZV9+
/XEpgNH5CIr+n89Fi6/FPfHWx4DbrH9+YPd8c9/XOQBYAiDVk2edJW1UE3XGscJuG57Xhj6/m9eg
uU+vWghLcqZkQPk1EvLS3MZ+Swnp6XymvCkKo9Bqfhsj8TRLaxzLL1LDt+KXwDvjKfT5TsbIkk+L
ufKTLQ6OWcI0uj7o2mMOuIvujBFNf8ZN6LpLYZIzCyPTy2GLRdQ1k3UEleyG7Jt4bVsssp9CXZ8k
ikMbKsB+CoUI/Ju3bN/zodbmEzbrL8a/qc8TaLfUDyDeyC3fqsHiAi62oTSexjCDjH5+JkENomjs
p3j57U3LWNkzKL+hK8kNOqqolWBw1wADMLsHhj+X0f4k3DDsF4ClmGRmeL48N3N6eXl5csTKo7sF
d8fpToJJmFVpfe/cj8q4kfzsELDgfb2G/jCjqn8u1q1j7mG9kZq0HrN5m3WajtItt55g9K1Lz7AM
++nxNr17m7a9I3D85RYXv6w+maNpfbg3Ul+ZYUnyILLVLVpdgyyx3SL3Nu77hGlRJiKFjdKUK4tc
2BsYgK7UJQ5yXJkCQOmO0nz2A0llo1Ain/0lpOY0GO2uRxeJkeLnzGasvRNZWvR5hkOQ4h9cwVJQ
Xmp2Rsrq/gt6drOfK7ddRzwUUC39X8xgNnK9X1ImHblNIeyd44WKt3XEX2dgY/fUunOMsxK6YHEi
jWcDRfqTzB5mOoBjwNxv7kU3B5s3mmpSTHmgKFHgfpMynLGXlsexoz2aeNWsvRlZgH1j5pQ0D2bV
FYs1o2yUe6Do28h/QwrNhCYGXYjMVrsAp2DOK3xiypBwXQ8Gp3EWnqujHkzMjbNfTT/cMhxNbDBf
7rOIudrVsuxi39DCwU3iwUpKA3qjjH3hhVBd85sEuZNuJjiVQG+bFLNq3t2tqMBN+SI7YPRW8AhV
A3lSxRJreXYpwYxl18DssTjgE4qFC+QScrsL3KBwABz1IMpHI4j7lgauZ/xcVofLHQSmCO5J8kPB
MTqecOxDJ2iTNenGOl3UZ09m7BoR8iPka2fLawfZvIFVVbnJc1FaGqjZB0dYhUEVATzYR2qGoyaq
+0WllLIjy8zLyP3MGB0AC5+bt+OI0q+delmnxSqmoibLpEeoDwPKUhejxOuSItgZ2iiFcyByhJCp
l8T2Rs556oibXyzIThz/auOfQfqPEzg3FsTb69g2z/MLXx4PzSxwyH9+1K2BMOSjPTluRezy/y1Y
DSR2O1H+y/MM/rpyDZBWC4soYv0U/RZ4AisgelBOgDw86id22my4DFNVXb/F7s/OLGN2WV5Z8M0r
MNIXWu5MTZhF7DYRoSPRAbrJLxA0bRP9XUEaFCxwLpL32F+jbvrCdwYFuTUckifsUiG1hiIbZP+h
ZqDZQezJ0LuFuU+r4L3moj1RXKCNP8XOrhn/V53a8H47nk4fz+nE9n/lGzfzlhLlPXxtB6gWSXq8
Ye8E7XPV5Xt9/JVwqhpHJLVUAPzv6yYmRhO84qGzuWX2922PJ7rfgGdpeBuh60Pv646YFrYhWHhE
gp3gCDFJTCqVTPyqFtE+1kG3tnT0rG+PM0kL+7wgfXGFT54gyBqqvZoKrRMIiSHPDhz4F7jTzmED
HM2PUvtbSmoGG+EVtArALNzgW6On7JGP2X28RE8IPQJlOdMmnHZvvGCY5GBfNggi0mZNYX067R58
IQJf4aIHCeavDQWAiI+6ysaXWDEaDWxoprXDSu+PJ6zddrpaOwXnxGfoKx1qW5BGB9ohkpFpXBeP
OBM5ZG3+6yD17rIZ4NeO0JXLrKcZ2W2+RcPO/cGy6tgYI0mH4R9q3hlKyIWIY7iJzUR4pZ3yC5u4
iC+6HhSAzWT4pFEmccYcBe5fcDp9kUQseUWRJtEuvQ4Wtp20QQQcVyZYuY9c8cBwlVBV+8/FqJo9
2407+EVNf5qGI0uUzTvN2lGsPW1hRD/voUN6k8kjhFfsYX4qXEwZN0KgOMpkfsd0I0Ptoh0ED0+W
vhhxdi5pEfTTFm3E1Ekom6r7AWTJztn/OIlxlsZ+ef6NLpJuI+IFcG6icNCNXrrwMFb1VApnRS2z
Ljyq/4q+DAgBzKg9o6ux8/ylUBOdwX7coeVcEIHsW8uHyQ2I8miBy4N3kAYM83D6PcqYDndcIl9o
5u/dQq5Ae3CRkZrLNtqi/3M+dV1u+f5yaGiwIdcHboUStMvd64xWX8bmJHyhDEuNfM/858uiHH9p
xbgZ27oTo38zKZM757JsiY0CzlfPvHxh8L3w9qnhvQpxdfYLIFqwOskitbnicAHPClDa+Qc7qpZf
dc2UBA6ZzY8W9AAOh978dFiIxLGRq4x1g9Ey2ntukMwz3Y1G3R/HZlUgQpZ5Nif6+ijWMDnobR2n
PVZoAW7/xXDpcrzKuBTYEVzq2zShWc0ItfAvu/Lk9fVG5AFp+xIBHeRKil893TYN9zWeSrOz7iVM
2JI4v0hiJaYAIc333nYMmbMAl8qfbikJCn/BqB5cEP8jTjH6PoARJfevBj/azDAlXlxv3kvTWsIF
UnDO0vSCudmJlvnQjZMUfiv5qXnWHnD5gKxg6f89qYBInLnwiKhwckoyX0TIA21VQPCONAtIAqtD
4mtW+bAyQYhdFSXat3oSQOl4HtqZ2iDoLVVkdYwQ500p0XeaLaoUwDYoBT12vWUjZ7aa8IvLwSXx
WvO7oZYWAUqpVhOc72AXSjj/TrRDk+M/+287HWlLfUVXdMZWQbF91JPqA0LR3UiArFc6EROVXwYq
F26jbU8UrfrvPEYwD1NKks9np6I2hINeG4yVjQCY4owYnpg+qrmgihRovWlW+kLydO6DRb82cdjo
a5TQUQcdAKMgtKmcybQYJvpX1WbSyvhTuFOxjHVgaD7wRsv+874Cb4HDKyEZhoFFc88cYZIvRh/v
aCH7f56DtoNOigAq9gBPEret52fOR9HaO3rHEFKSsgkdRGyOhUg4nO6vIptaSpXOURrSTN0AYwXP
TFSxRvLcwzvaTrPgJkP7BQGZA5RzxIfMqt2JwNynRr92aGFRzsW+/LHiz7J4V5NgUATvS/AACtW+
iwNmga5C670BJTZgizWqKs7wGMhmt03OwFJ0yrlXayBmzlz9Z0mKwo8nhyEXraIDqAgbWKz0JXbS
j4xLUL2uqaKDBVVk/OthAs+ATqwpL9hGi1mBzaOgxi1UcLFOLuwm8/COPx0KcAv5pGcDrdx7j+UX
ZfWoZBy7F5UygRliSzJjSu3kOUz1qhmYMWYgxY71OfgLDOATxlYlzZzfrYcXHAcptcEKiue6D5Pg
hbP1d7V94L3piTvp0AFgMdK2vZPq8PpZNWHkxMW/AKq6MEQj62Q6cILh7LYeMfNM+zqHU8UynTJW
KSYeisCMZMoZifw+cAit7y85xD9GITDd2pU4noE5lLk9iMqfwZBa7gSgxHySaBSaOnSAuUT9Krin
XhSUrf7ZRVw/MbEy5BeNrJsURhChbqlV7wthndn4ns1O2AX/AqvQpoxJxgX26B0OfQT8ZSNB6vEU
wQnIUv2w2E1s/VjeKK1oIE4Zp5d2czqKy2FDI88B8QAgt+G0SnfRks0K4Qs6OXNLlV1i8EUVZ3yf
5CYrbyNWNaWoycFn9yLTQ2R0y9EIBcRbZqyKCrM4V5ajRWHVCqBf62t+iljU4++sq8+aR6QpIAQh
xj4cvOq4eyA5O6q6rBdbaINr0B5NxrKYfStPh0CsAvun+FRUZZVep6OC7PuM1oKC7hpzTtGC6g3Q
CUxugLEsJah8CjM1ByUP1BTuqo6M7Hgo/QzttF8VjZVd9RCHxnniLJcju38mmm3BadB9uwHUp/uP
DoK3/ZAPSQpyKPi+5MrCxjPWYrCs06WwRjW95S3DsOleOO67S8+BT7Bs/zw1JkQ/MfBwFqZxV9Oz
n4dpLk8/yBLg11Z7XwBBwLc5z0ISMc68lCaSh7HnHVGL721YQAMMolZy+gMDIOa1/pZkkFN164Bx
zVCchIw29l34do+ZHnTbnuje0o3IGV7ru1H6M1+D+qAsobSylrjdOjwTHlnXvGzF1fn02aF+HUVL
f86v8KrMFcXUiOu4aI+wfPDPewydYDbwMy3hxFS852BVkf4lcZMoAefSyp8X5UW8vEgxAaAqgktc
PLgDv8n7qkJ6wcBY1s37mnRv6ncA+9QNsOlzWQDQ8jLf8hHJYM9UIT42sDn9c2yIVFu3TK2Lardv
QCvnFeIK8ADc3z9ClRjiJKpUnajhQmS+aianrIca0WS3U1OFAdxdICmqGsjQpMqCGhuBvr7FOWVI
Mcy4YWdO1Zwnr5/ba+RDkecY0/CnT9n7ACOziqEzPo1VVzOBufcxHKvFChFFjXPrD1V8UY4Tuixz
97wIwMpBjbBu/nYmLufRlkpxbmx97grQV76bYoIfcEajbSVdkJNYzlDN3fd6/K2NUUR3ytqNXOQT
kJOnMtpdIPncBJ4KkK/xiPvbOWacIxzSwUgOho+pelzLfH2bVcsuDS1QT65u6j0wNwAhsgCQAeO4
aRhGL2FGEbong3a+nrxgHcEOj7Rl9/iLHkS4dBugJLHmEIqG0jIMuiVAW6Icnumrre6Q+JmxeiWU
ZZW0ycxUe68lVLVuTG27OUq5BBBJE7WI0umfX7I9Vx3KeaTamWCPDoaFHe4HaQmrLoeu9ji9Mg9d
KhyMRci/98Bbxa6GyW7SCpSWZqUc1fYqkfFVDiTbroqi2cZ8uxaTHumKc4AatsTIDngbDNoWVMA9
sSybYMnXx4Sg/4kn/1vzCSiPML6ZVOo3vzpv7fGSRQ91hxZYLfviHqOi20sTumrFn2/3gbPmrGx9
uMx/erwqdSLPGRCZF74FOvzl9mSIXEoHabxUYck4alsyA8cQUUN/L2hLF9x5DMepp0SiiLABCIFq
BTmFNZr1pF6bIo+GBR7ellVO6War6uFpleIj1f305N0Yk2WdB6UVnIINl8RXeEl/IgrHJsfrswuv
Ho7TVArHjsBaRNHnTq3Qnba7jDaMwz4qmQldbzXXA3P/liFL1yNOCRSVTXCLz5VefbNISV6HRiF7
25UzWi6MsDnB0aRYpJYXvWZSuFTlZ0YioQa/9zqhcyD4OFJbC59TfxRdURZao10eS98KhXYkuvRi
/nempMUwSfSJ+//cavUxNGH8Znvq2A8M/fVawO3VB5O+cuoXXVESSmXpd4Jc2xfsHeoT8LjZC3Vi
WxHhIOOXmPT1mrUi0P9vXqNrJup1Vw67c2A3PlbcGefgf5xoh/2WHBbbkkDs3xKJxT2zIEtjn6Uf
xOk/GL6jtquTLiAsxaxBfzkPl/DJ10BVMEE2XVPY1xAD8aDt+R14y5dwIOdBj6NAJWvfFfHjPug9
XgzrhYgjC4lzZQl9mgEcgMy4rrER1Othfj/qZR1kxAsAbNtgc0271f4z/LkG67DIYOJ16MuMbogc
jso20Tfo/YY1Yk2fSWb3oK0B9HJAt0iMI6jH9eOLCqPiJHl7JmjqIs0z06v66ZL1cjvbEM31w/Tn
ivf9Jn34Ulyl4vpe6qZklKJNPv2apiQOiQEwhcSvZdaKU2MtTnykxTRZfMH+jsILgHh0hnXoL0uo
4AOdX3KLA2kx1ftzYZB02Q4WMx4EUHADtYezu9+VGPUmFE7Adw/xPkSuXSSQjsm1I9f4igYfJDef
JXcDFfB84CNFqyE0a4AEumKYBbGL5qOIV7914p8tHGt5Wlo3tViIblDxxmK5SNuZIBfZh+LE2Ab2
86x4DYvmdBrBBd3kAUUB9IVf/Efgf5qD4bXdJNOfckYxkUtPMnTGWWRh0u+FF2swo3eX7GSrMcYp
YUb+BdbJSqDVntw/UpX3eS5jCyC7gZ05mfFEOBGKSmJofSfM4atGE+rOpyQFRT3rklrYWo7YBnK5
2XvaOyCvJW9/ZaGqbPUSffdx0KuskVyCIOo43wx66k2uiYrVUdSye3/p0J1XCvo1E5sOrGc1s5bi
gbLtzL/Q7fWza+m3FI4QYLGcQYua0Hc7u3Ymt1UbLX8BU4v/u0T5QbdDr4gDe92Mf+WFjDza+5OG
nZD0Urcxxa/s40xbYFQMC/h2Uv9EaU9z5CFHO/wmCyhnCZm69dcEB09a5DgtABOlGhS/4W8e5kzD
NIlQeQYQys0OCokErdpZz0C0MeqmCBqBNpsTB1SfrrQBmyj+grRa1YScugjTizFPd+GuH6dUUejn
9mntA2gR2nTk7VFheEcsg1PTkfQhICWVAISLGRY8MCuUjc5tMvGI7K4nyLdgqnVVsPPoQ5nWDRPv
hUpisIT/b9QKHzEToXGskyoBvhMxhJvXfowtGPKK3MUfx+XPX3gtV86gRjGXwue1sXnP+7zR3Gil
LYJby5Wn9odeWWBDFyf21/YmHVDx9jca4e9e8tjIdi9xbKISrvwPHz8J1M3KsJrzAvorQWdoNWhF
e1hJtDwSpivnBSbclWUt85KyyxYiC/uAlbpiO5vJrFkhidlV6oHsEYAbyCcixLtyNlD/jroRWm70
+gNewwNQkkIrPX8Hb3uGQ5hN9dHg/chUa69vnju27dnFb+7ehXpg3D/5twc0L0EfuI4zFU+KWXMP
tUlGoyeYTRhtxGjuxJwej0OOoW1eHkQYRYpAggt38bbtMcQKmFfWvjq3NKmKyaV62Ijnc/kH8PqO
bBBA0bt8iZj7mh0UNpb6U4dxSGslhUxY8Wh1D605ZCH65R1pJMWhkRxSt4zH1OxnebBUfJHr/9I0
6F3gXEikmmJusL7o18/wNbB2B089/6p45a4z6PrrEHZxM6wXenVud+0zaOUOs4hH5X+cRMSp+BDw
WxGQIsnfHsEoqpRkkEc2K24iZWbJyewGjKeucWnSZc9DMlLpSBE740+g3t3sNH+u4B5uPMKzMmFQ
uH0ds7yy3aPZWvRLVOm3Pqr0fgwaJ8QsIK9nt6T/J2DZ4Ck3O3svjPF23SarOz9Uz98Y5bGEo4sB
SXlGBYc3MF4QYvNxhbl54QR/2M3RDKUWjcHY7nT1ocI1d4qb8YHOHN6DdJ/GkM0Hvhqpp0V64f0H
Ij/pn2eULQ/dTT48V9PSqqA9YET+N2dgER+EMYPPCUieTrQuO8jUqFj5UNDqVTtZSEtRFyLUOkuY
piw93iI8s4cbOhFsAhpOan5IldelaZ9/fBUpoyMwMgNTrWcSFsexyr11S9a3LDGtW5wX2cKzqjao
OhHw+ZMpk8ghUsL2cJWC6nZkfMAffDo4GCf7en7LIbhdM4nrRSs3mbuduFzoABu+4juDjqSxDw9s
j0pazS/HqtkIRrpyaSmwClszm4C339Ix2jrf5MT3RRnOgQhpmLA7CGjbZBUK2btRAnRODHCg5Xm2
ObEiqMS8J56y3bhAmHCY/Yy729dk4yT9wdaFdN9ye7MqvyDChzAaW+ziBhq0jYlJyEQhAM+erU4D
pFFdL/A7zQIFm8RWPqkEORZeEJ2aADkACibTcfJxEVDUwOdm7YRy1BdfJEO5lqSY/3xkNmhfUhdE
nvSMPo314GWUb0fjtuR+ngZjKtG7goPXefnG3Xj+Jgkb8vuzDCiBtuvuVnV5P3QedEHbY62CrhTW
y6vykH8gK+Yn7MGNbgNnt7iK07PY6O9sPGkDyoDxuYIOfQm9d3D0ZtCraifzEIPFtD6Sed87BQuM
FNU7KhlycQkqh3lx8mTtvO4Tj9WecH0NxlUp3b+5sVRwCCkikjS5sC/ECcSLshoSl2Pe0ls+6Xin
1Ke+ITMM1EhNC9JX6T1oIxRqUaEBTBRQirSk7Gfxd/AspFynd8y0QPh4IAIL4SVReQ8m2C6GYWLQ
2PMEIOE+/1rt+pa9A6fBJAjsuxyAGsHZfKsQyOAImernZ1Ixr+dZf7IDMe5++OfiqmmigA/cMQNt
ztKEjNYrCG48CcWsSCXCm/OeYrnYDzQ9/GYQciKop3dKTvAaxCCf9oyu099RNRX3VP59XuJ27rWG
CYUSB1U194twEmvJ7QKZT4r3r1iU11CZMNOiBufvx60Ia9u8CqcBAjmLRypkZS/SZ7JzbycItDYE
urjIZyc2AaHmMdGn0TmnGt0dbuCbduF7FG8kTY/ZLuV55gRzRQeo6zx4MI3CB8PULWcNjPBUWmIZ
j9ptw4xA+lv8StIMk3bTNzcD8Lc67+n/XxkpFCQMhcUmPxws6tSQqdX3Xt3Hk2TWze6lAqoSvPH+
JHbDohSH3vAIkLAwZBKHy3hqOPux+c167Vzjq1FUbinezTIsjRUK+IYjhlW6Eozt8YZ3zQx/fwUU
uD+6smW0CMDzkiwGk7oB1lKJ25AWlhZ2/HfoYW+8ZWBY/oSbYRK/yVZRA8bLg4katJ3Eirsbykuv
zzD7C2mjpkLWhjEyaSCThU4tFVPvjL9ENOgfg9uc7tAdTiAjSF+jCHiIsakadojhrNJT6AEzIMD/
ni6XCF9i7KXuh0Q8e4CN9pvncXzV+P9o9wCAdOD7USxI912qVJimL9bPdRp6VfFmB5cb/fIGyo5/
mbQTjDechEaEecRfILNrKFs8gLESh7Iyj80S6a2l1/Bjyr33eT6gTlr8ZhML7LALh0dcaoWTH8m6
vJboCjjzk34LS+0V4qmbVdvyY2PS3LXvx7/7aNUs9KVDTVpT4iC7/D7shm2FHI/sF4snjY8SL+Tp
xJ4UoXzXNxddi/97T+ShPbw+LYFz2viLktxUbiI8faPylYcKzN++ciphl62Zv84HT71ES2thonl7
tDfKVhFAYbwkGFs3t4r6ABYW41E+FZF6Jr3pXGyrjjtvkFGEZNWvfuex+YwRHn42hI0A3aATemyl
XtTI9nLzgHX+sAkGPWidytVNS37rAsDsbM3YyYJhTwJYKf96WL1+nRODpeftkR9ReYh6OAlE39hM
A7k7kBS3G3E7EaKklFT96GKYuHmmG7mEsL8NZ40S5gKdQJTKjG/qDPwoGwhoWgmP8Ed1NRqFrrUa
eYOR9s5dtPv4HYYYVUtXQPdB9LEQ66cGLKd0+N2u1mp5frnHlcZh89q4wNrfxNVyLGO2BEPlz6Qa
uLXEaiK/LK28QhLw2LE1Y6oJz74/K+dfWmXF1uJvo4C20FiQxPz1GWXZl1WnM0lZSaQe62m3gdaz
zK9s/MZNkQfuDy8h9Xv9sdgBSx1al07j2HpnU6B3fVOMbtOcioR1WYjGG8zEn7WYFfkOK5mg0Fmg
4M/PHdQx7vU2Lm+BjafianUa1mN6L5GRaWPlZ1lut0GoQL4WS5nXqquZDgBCvQ5rW1qbjpVjXQDU
/u6grgWl2//oS/qHHm1afXp+aolOEdVyTrxBEc2/eVv7zc3OToEUOdYehfcTDLhNB59eBNStd3Uh
bFNmParPqg62dh8pHMaxWAmnk9Cdb6wZ/PEHjjUfXjEVY3rLVRNHsa2G5h5Aa+Lv160GyIw0f9Am
4AwtMtOe2U/njKT9KHp+Y3y49Tg4a2IZqFO+41eD9Yf3phs+a7sf/WTrXIDBe0nw9hOQUwKceS0k
toy5j01g+gsmp7M/YImEooxhUC4kjcRc1qej2bBiOUbqapmDvdeBTh6YrXfDypem+LY8+oLz8Gje
b4ifNJPd8afrrg3SU4DjkUb9O4tog2Q1OTD0jLE+r7xvZfwBEj/Qe7+MbFFxXHxvy3S99oVldgEf
nYWkcvLH7hhxzZNw09qjKAPBam53WtGcN0UfwYKKkbQCjn5hRC/gmR4p92yNzKAt5746hVvIGzva
G/cGtrlV36pqZsUdwU44O/LGFhUoAkABN2rxHnx8cYxu2cNBZfuePg/mm8MEgiOSF2S8fRkaLC/l
AtfiaZqZpU+hScPuFbGJ6/7lQZ/zattg2ZTCxw4R54W/7FkDVoGaeY0mfbCmQ3PtAcu79aFC/iF/
27frobjjR/TxRDw2YYX7HzgCOLw1TXqNpp9rZY/UV5oAnec0cUNP6djIggp4+QZG7vLKX+RIGRcC
UGWU3kILAlnefxkvCGsK6n9HIgXgflkgbOaNi1Bu20xjCJO2Ngptn8p7kF/aimHzcmAX2cC+Wot2
Sup74kTGUaO/PD7RinKyre99FHyuf6ATU0UUCsadWY8XS+91ir0kNqEuMzC8p1Tr4NjiHmhdDbDI
aBTozMnNs60u+fxSDFZBoxhhchaJI66YKjLQ4leJmJZjDtm9ex0rd+nAHxhxSXmbse55mijMp4qF
Z/8EZ8Qon6fWcKj6wGWs/wQroReODlfDOazmqu696+8Qowo1xIUogJrY/SC5R6vmw3bhxTHYkUOB
8r8RHPvFe2FijkChM7C62ijdtgqoPFgbQro2sg6aY5tKUgUiC+MCTSPlK0bqrCo0F736SqOjzzsU
OcERo6Lo6R1VlNvR0rcLwyTdIK7AH+qo9ZK9l5h4dce/frwvrO/UrKeJoQbBbQdTRiquUrferrL5
QdYF3rJpnwtN1RCpd2JCiNddAVIme5QEY249tVaoBEZWIf7Es5R8uJ689YdHCZrJxNkvDAQxOv4U
bxiniJ8sN6VuowgYrZl/C3cU8vvHvKausOKR5DYHAd+i8HOHvl077/QvFkvwoUKvRfMO1YYd8Xjk
m6DRXE05poyEh+awFrPuOZ6SIT5VwG5SODIt6M3R0ZQRIyQECcH3UFiOPiT4IV4AUlF+CZ9WzYFm
lNP8+LUVUslM/NtG9uOlVLlxufuljqaqOjEjDA/HhSbSGrdb+Glh7ZKQo4tYXbq8+ld/Au1jRnWt
xFel7ABC/kGDBYXVairouHQwIKJ+RkxO4X6hM0q01q7EcYQFy1aq59wLr1uGz9EHoIp2j5Pf2G1h
FmAT4XWM8DwhmBnRAA1WnYFdb6t71F22qPjXHQsGRQ5Vki6UXsP4pXjf/Svf/LDdHZsx8hugqNgS
5IkzKSmRru1FkZWnGMnIMKqrDyo5D9CE+KuJy/LRtYhkjn9Uetl3mNKCNv2zMLRW2ZaMzVUxLlsq
V/lW8AT1unpY1O661vLLvZVwCvBhndBUV+NlZmKIL2VpMny7eg07+9mErFjV3sf/LZV5qgy+7NyV
badjF9vKfFjA7jO7fqoSQprhRQNw4Sq26h0/08iSPMNMvkqF3y0tysT5M2KrHJkxxw+2/ockIM1c
nDtHxJ9izVw32RMdUq8nz1wRVnGsDJMi9ibF/h+UHT789Z3NFRFHo89XQle5P9zG6f6mwc9sZZyL
58EyWso6W/DU+/HP/s24GLPUTTC6HEIsas8yM64TLANXC0EonQcIy2vYd89IHNmUsIoxIKaP5HzP
NejpTjMNLQnLfuw/R+sgP3epwQZXN0t8ZU6pfSt7NmyhystvlE+3NsKuHnQBejcFTJvw76fB70/s
qhVEbkm+QrTEg6Ed2CfHVTd8fvZ9e0V1uOoFUHpSUFhlk5MtSUqbdiqu6aae4OFHLqL76uWXSbBj
fzowdiOX74VRUMMgPKGkZciDS2JGOJKAvbr7FpeLrLo41WHW2HcqTlLIlNdSpGmPKndCwJ9shBng
bvdxr980jbqMxYlyOeMm+eVnhlKrdW/amIL3HY996O1BrgKhBUhe9Y8oswLdKMbKH4nVK2jH8PuL
yJrdwUlzDvjIJvKrP/drT7IB0Q5Ywi3F7Gd4lDqbSkql3SoVbzBxCDLVSD3cHJ2lmXz/vJpTO1mw
uhSD1gk9Hl/GI07Hb6fCNUqV8sYmSgfDBvNb+am0Y9MOQJM2Be+DeyPHzgoL8zonAXuWpEfyCC7a
psq7U2wa6lHy3kEC0we/0yc9eCtj5/G+eUrFF6ljKIImgKwKUcaxXh7tnzz66LfjYtj7w7o1a/Hn
vpMexIAWVZ384CkeGPA/VYgryhPkvno78iPXMWQ6OKmj4mE0vPMT9/Zfi/G9qwg9kZXDqEu6T8wE
nxw6u5xlOpXD+Akpb6KJSvC/u8kUY5oWImhsEwk6JAayD1vTmu8FKBiQDp069FrbGnVjT4sw4Xcm
Y2XjQDW9/0Cr6pmW5rrR87x6N64iXpVPzIRfpSfxwxTSdf5QvESZAS54x9Qghssx63uH4I5uAyte
tVTDdTyLbcRc6G3RcZ6BAdghtAE/sqogYyJf5fSudkbULLJzEcLMDyr8MUEc/eZZKv1PtmiOGbwM
Pa+IycTtGc7jzLz82rMWq2wSak1sVfNLGUi/arJXX1VLnYLxyvqq/d/1s2H3BIfctSPj/GUA22vC
UfMrzwm67/h4Z23wQGHoOqzi7d6Iy0N95V7dsa3gbBkJrXxGYGc+06nbMNiyasEWGV1UsSHw+d2y
jEZu8BKU6pAqpHuMHcxSk5cA5fhFG5mSHwicia84o007FX9XS+ivbu7UEs37ceNiVFWm623JEAn7
GUtx8xBRk8MxOFOaq0Em+CbBATnCzlH6fpxlPglvrM+xaNd5+zfJLFjrkYRqCH/n5kYBn4OdHm55
buGru2g7Mvdnp6yRaTeib9YgFDgygxCBF3esovGYXDoQKEd3M1pl2DRbxw4K4kxmVbFu14aqvv2I
3m65htD337vxr03ToyinOJ/7P4N+05KIcPGtwA/w4NL10mv+UK+DfEx8NH3oiv+Mfy37s2SMSmJa
vj8yBriCcJj5IeVPunc2LR9UTHoffQIoG0TE2WcL8PJ/feVW30DigLllM2Y5kQ1FqUZw4tyTfjab
5nE5qqPlgGtquA/0OduWVA3pEyH991IAxUCJ09uYBuZYlfMvxEJZlgXHgwX6ssOXhisvaNwA5Nwd
+VRIvrAIjgOIt1gow9e3CX8bh/Yg+HfrSAlCSXi1tbR4x+cDiagTqTaDmwu+hL/4QUA7FxdJ0RPF
kL/t5SjnnXF8tyD7Y5uVsg/hhnzPV7sCsXEn6IefG6TPlhz0ZF5NMU9OH1wepOqjloilORWccj18
zoZgHIhwlpqUIi3t3QJ3PfUUYed78LiEpBSRNPm/OaZauIS540a0hr7mRPAP06SP/XcSiamJ1cWh
xpOK8gEvxihwuhZtBQd/poeoNVRVMbwKzF5dlxVg5YZIXrXvH0B5hXcxNtBZ+j9e3RS3JZYK4bF3
6u4SmtbbMs5F9Xvbid2byCqj56j9AQGOBD8lKQzpvvQfJ9ULvloGGxKTgqFt+8qwy1uOjQVTuAuv
VVUlufIRCDnVmVJFTMQfDfIQIzZuOeEXD/F4iE+DcWWHc7YGq4gsmpbr4ems2CyD1XJ3Ek2U9q8E
UzisD89u6CiF65zSUaCHaHUARxH9ksJ8D/YBkyCqm08/9L4svoi/5qYtxxKLWE5lT/BaZxGSB99O
3sxmoauN5Ty00Bqt/Ad7kFR/tLkP8sfXQqdFFOFp89OojNzlBPHqzh1Mk81Ob71d5GlYmZ/oG8mL
yab51G+xqJq5ctRPQtjOOQte6tw7nlhQ96idREPkq49xvWmck39Z51xj9fLJnMjGY15d1dXAEWn6
x0A6YiccCrsGV9WmlMtLHuRTc0vv+ESzTEWb+NhmFY3GLwQhEkODF8r2O9JKDRP0y4FW0pPBAoe3
78gF1hAXEze7ilRZK4x9t5lFdbIygF506ArTyCSuNHNsVFmWnEDhmwmgCkvJmdPu/qOXZLlyZHEf
9UR+o2nQjumrC20RN1uhaVKsYkrwoE0wwU3h80MZfc/tjh8ZXk9fIeZf6fS2OxecUxWqllUMZ0L5
nsZ4Fo9txyMbXSFvHMbhW9HaT+/N9hapayhah2mjiCGT6/77owVPLKw1wyVqfaiwn/g+Nd13SNac
LJa1rHYDi68o7tpS1JAvMPKt0TiH61yIYZn1XyPww8N0jNes2CpsfAvT9/WxLHp7nW0ss8+oyI99
pzVqyGpVEuBW54D+S4Ykl3Gn3R2Gz44dF8W7CkcE8hmT1aykycqzYSMYJtX99VB4mHtOg+IBr80l
e+GZiEEdie2lLOwGdkzWJpgzX2h589mZoI5lvzsJBsM/4DvasThRg9lQzm+nJCmOUTyylniwfRF3
KRG4ikdm8WqJJiMOxkLR/rK2/ozwF5PmTSY4yW/I/ugh2W11JUh6dG7wNxkyQlT17VJf+Fkt/Jgi
50+PJlBHA5VRVJFzkxrPZbuwKhWl40Y04ihkx8sMWGBKlex/debZtlewftTloybqls4kBXEcQ1Se
dGVfrnGtg2K5kr9gQBeZLr4r0HUHXmaBPUvnjH0vwJ4/+A36UdoHTmpPX08269rSyOUUPB6kHffV
gMlfKfIrXtt5gXDpOb//ZBbx2wgnRx/AsSuuXMkbTuL9Ail/dDyumG58g/8aufI3/Z/+KAZG58m6
X95NjpHZR3Ca8WLu/rNfEjFKMl0NH1N0AyWRAZci0RXQn4c2pXZfeMfqFebyzZtkE3ulAVP5Vj4P
nUpMTlQ+D/8D24t9QqHW0+r9QYFPn9GHXoDcVQ5scaAOVfe8/is01Rnaw3pnU3Cp+DMl3pf9TNu6
cXIeAX6c75XdgeqkxDz7WlYrm7nWXb32cZgkyGX1ilhEril0avl9aicKW2/P+v7w4XKfj8zfMBnt
EtMf5/DhFtuSZ6PcDFKanQUS44AakIUkyoDZzKOhgG3f7p6SMyPko9QN7DdJl1x+Las8swKf0KKC
vZluzvmiy2Ha4/8ki4dszIXiHW1/7BgtFzX81RE3uGRD3PX5WtHSud/ZWr/mFSgrVxS1tB04QKt1
10Zi6zJfxsKX1Hi2daJOXgdFmh5s6D3X/3ENJ2n7+BehgMVtNLtkdIutgIGicwSd6MqM33H2jsKx
dla/ZbF2JAzQY9bu8J8MS8jQRXdagjn1LWfWkOV8ZVYXJZmsgdU0ShdeYKdjvj2W7UZS7Na2akxq
euwtWLegVrXnO5DTzTVj4Cq0Oz/aDlwdnTwk4FOWtRjR7WwLERY/ym2ro75O2aSZyW29LQ0Tpzrh
GKRIAHC0nYD5AiLcLeFn9MteKVhaPxYAqVRZaEwNZgzBospNBBexO6twwObNco+2n7aW+a83kThH
nBwEp2t2df+CjfkZHPqjpp9fEZ+51DUrEAaWWYRZ7ZaXStTsEv4bB8G1O3iwq02VmMs/lIdBXdiA
iUERe8TUYZbKbh+inWZlIIEC1q3/vdNHxigBPsqqnLOf+mclrp7kUdnT5KF2ocz6KRq82P1ecicD
gOW7wmkrCDPqJoY5eEl/BbKaAhuUhbB4o/C7tLqiKMtonsdYItIQMPLF82acIFHv9NglTAsIo2yo
IC52mGUScJXizxCVXR9f8+4RquaT+dJvjAqKOKaiLLGd6VosFfvFKw1OszXxn/WCD8TLhLI98C+D
he5pCTEhnBuc4Hl5Ml9asMKZ+ZyglP4ZKGRNTNQDeVbc1YxjCHxlgOByHXXwtIcDOIAYtjJC0uCZ
KYXutgRjhbT/fSLVBUIDpq0nelDmAja0BbPH+SSxbD0WOm+rvVhvhDHcLTZVF72Sd0BhwEXp+bN+
sd9SXMo6/j7vgh/xe63eF2iBSP79ZR+BeVTivzenwt35amwl9zErvXzHEwWLTBrciUNhM00ofI5H
ok6RnfA2PZ607cHyzNe8Y2fr/Y2DY3KUJj8reAUxYP6iWYl+7sMAJ3c5X6BBWVgXclpSn+V1y8wF
g6PiEYESkIUEK2daiBHQAaAG3VbDX09PIhV2FeMm8yj0uKZ9U88uZflWO+OgY9a2ps2tVZE3pQEm
mqDb8UrN7o4bdtTUAOBcTFtN5vSbHNs0J+2J0PsRGg4yvEl97RPV/NwkqAn3H4LkEEyvGc+oNKhN
5ihG+2nHhdV871ZSvWjBVXIu9+kZvvC+/GlPhkqS7Hu6xAe5J0hAPdqN2NOt98ZLAWZ9PnxeZc4+
kDu7aWyR+VFrbWQjIhOoD0r62fQKnaHejWHkQ93OfuWWUpq3t9/6MozoXYZG21Q7LWtszMwIiOOk
Jsyzmayj/ga+cShY1RRqxEBx5G1oWq8L2NzWUlprQHgkFNzakUsiCiL9fM8Htc6HPoXNFzUNgXrk
XNX7r9+yX6+fAyxS+crNAJzqCVbbxaG+cCvkY9XRaQIJI0E3P3KQ2273FtIeBDp0RMS1KOxFL7rS
K53h/0ussqnPGFxivKqukEuMl3B39ZgDGm0gJ68Fo8j3ylQ5NbLV57snxrmZuK+6PmdsGZj1bPLI
ks/w90BsVc4w6CqAzVLiP7b65PJU7WXJn962N/QGaQDyFgAsfQw3WmIZbhMfVO4N5+qi8mFTfE9r
6PLlr/Y1ViMqmDf5xViZlQh4WNOzrRP56h1V4fco76Fn4LdokyGoTWdcuCT9Ih6GadLMnFICRNT5
LXZLti9/Ut306QaqJzv/z5m0Fq+niapULQN00LCt6vDNQZEXhRLFzBvmiqvunB7jznsgfleS7hOG
u69HzpfnZzAcUoRYsZK92SSa4SkaetE8DCMk1yiFgSVELU6fCupGF7UiI5KVQnOGOQgOWgKJR+mM
1TrYTIOWSqzyOvczdrhoy+57TxoO8RFm+6+/GCENhw5HiNMFUKpF9h86kpu8Xbq6k9oGTQykVfx0
FxnelLQA4vR29L5+NfygLVQILGGyfalKgU5CpPzHvGvvxy2MTjrlzZ2uxvSv/5wOc1Yyfc0uXww9
tB1ogXkaVeZ0h+cPrCvqctoelnULpdtiiru9XB7hjRbCv1iPd88kBVgJAfJTSphmpitbmT9BmE4e
NbzvRt6A18glt3ZXF/1Wt7DxfZJtlGGRiKfPODfPK2xYVMF73ssqrX6Is0mOlgs8fxmEyfg+Q0M/
rmIMufUlCMPOfMkHN2Yb7Y+mvRzUlNLoIzUsO+Dl/k8MsAIalH497FnYIpyvlxVZaSyVH7yCuxyw
ViCPYt2273GhXsKxVRC9HHhSsy7YNVPvIcizH8rGV0de9nu0VyekrzNCp/nYYrB73dhVAxzu49kJ
AV7NGIWWZVzFvTbfzKBTk1MeBWl1u4JUG6AuC98qCBSMdUhwM01h7X75fUAV2h9h7iTtJs1bvfit
DFSI+8oe0BOt2zcKhPWrxeIAzTARXdbo7Oh/pMk2sCOuGYSlviZDOAb0F12gzJYjUTvUpekN3kfu
XyfCgrkQYYUrAI6H4xrS/mCO4EMokaSO2BRoeK3LblPPyeEYJqjz2CQ946CP9bLO0yggHNia1TJp
d/a2sY0PskVPWm4oKHvmhoE7HiiCXDpMzt9xXNo2gvydmfP/iKOJIyfpXSK5UZnEzVvc6e+hGuDr
gYEexTQf+gkoJcamLy3NSCSeJC7HPAXh5npLDj7FVpz2KiGGkwLTlaRz8tdayBYgEwXCEtq34uR+
3U8+vgGLpkMpqsjvpbbLuvmSAkL5dlz9vP5Sha26+YPglKLsGQRXTqrDC/R1dEeJX/dghdV8F0oH
huLHrmlA1WkhwCqLJ3ID3943n4zElCzKo1L7zZklLubjW1BAmm1XOlWxdzm+E6qKpBPHRfPvxoSq
1fy0cw0ux4Eg5PIFVYXGGtjv4XEm18lyzavlxT0ZkrSk/jx0dHk1NI95+3g44K4gJSlXIE0Lfvy/
AtEIuxL7ArkWglh/eXu6Gc5hHWjfQWrM2kalAz1QKllXHzC/lAE0rQz4UooCRSbOdJZ05PbX9EOs
Bxy/mjX3847+7Zf7nCFQIqKrczlsKa3OFyMiUdZmv9jcrx6/mzITVdZ4R8EKE83/8AUH2vjUaYcH
ktR/CdckD4y4Sz63uv+t4umvofEp40aPPdZ2nGHUjwBklWJQrkeK8mh4iH42sYa5Lg8nPhVfp21c
1TnLIYvvB6xdh/kRw+6tL6JezWvnX0tcHnBTa5fXOOICYNbVTJG36AP8PptHBMZbExbWfa0ndoYT
2JTLEtqSz3bEMpForpmGyJ+dMAcllYQZB1uBYqQozrfghPtATh2Pqm6jVpEmWSTcwjBFBjwHOTIN
wLFAZ8Vn11Lw00mdhQUWR2PCwYU54VEjU/UmIpdfxNa0017jcJa/gdc19R3LyOWFuIBtXgYKIs4C
6K71vhriHm3v4vC7/OFm+XI8wNP943YQaS2ozJmZbhUu+b0NGAfxbr76F/+vBTc6iUZkT8Hr8aK+
N/hyLA9prPDYMtWCOwyBdkQLz06tUo1AjpT/0rw98UmOjyha+JgwhkPVo3CklEHEEbevbWYhoF/L
LCI7sdt/XZsJj6lydYUSEdCySln+DexI1RwNSWA5MNmGpEXmJvDAA0m6QvzKTC2e2+XuM0izgSJO
czX4FEqg8xW4ic/vLoAtfkCjvRn+3rw/8QYcbA5+ii/KAO7NQvyWq8MimbwegKtxRScIaLmgXVcY
i+51dKYLpzToEtpAhMNHuhlQJ8fzN0WOscj0toS7RDFLQip0a3a+0sU6BR8WdnBi73dQVsUJklBP
Ivy70JNl853Ij+S68W8r0cf3wWoK5IomWFBHCTZD6ZL0bSzeRm6AzWu9OKh2rinDZBI6Kt0rcmIB
PIH57mV7EsjF83PbO5mOFfBs52Kg8lenVmzYwWsBluNtKveOxFg1NqWhn1ZULTcuSxqRh0UEuC5/
+Ht41l6n4+dLxR7pN5NpHeSaAkJTx/xrBvafRpLyjXW52VHq7CsHWr8d1i054hs8SNbmP/NCwgON
spBc45lgs+3RmRie3e3svWclH/BKhYCPFSQI+LPxnJRwQKuVCnzZcIjz9WbTJBit+rN//uhtF0tE
xhufjKpnTZn5/kTlWTnUyaE9PkMBHOcspicmPyP0N9TXcCj9rJM+yVbU5X8xulsWqRk/tgoZTvwR
OCCne2IIT1Tw/0n2+HCBnu1i3s57wxjt4JuTCr3iF31MB1IxndWSwTO7JwmF7Ru5Yhkd/m0u6Cmb
ggnJXfMF0gSKYaRNI/F8sCLcaPsfUr79wOub35WyjKdndEcI7u+TLpRjq2dZuq02RCyv79/zQuMu
C4fdtJUlVCKhoVYSGjbdtYW3ed8o8Z5nxwHI+Qf8dlCnmSv650KjZaLQ+NO3IozewcfGk5JYBvHt
OIlMKoe8EuS3YaQAR7X43Mz4dwGrcwzIf+D+XzH9/+eMCmmdwSpbvnv+0JQUaje6zoxUzEXGbVRE
m2GBFeB6uursDJ9DqlIiqV1WrGdmrkP7Xp+rAr5l9nDwAO+nqLl/eMaUZoeKfs/lLV//Muuyx+Bq
dmtljGf9ZZvw0X/z4IJClF+l4xplHAmoy3rwfrNAoAdmqW7KY8J/O0eEuabfxBDaWJjfXdxOiKNx
dgNJ1zfp9koNAZzlQ4pkVdVAHLVrG0yvXZFLfjN1lLemobE4vPhfVCDt0iL9Is7tCYJZteFQzbu3
H+R6ATPl68lXEU3jNkedLz+fLsv+zKcR7aJTzDKIOmZ+4uMusHAvLWYY8X9gIYVvgCUI9t8gV9JH
6r+Q0xuH4DsxJubQpe6/Y2HIza+gM/nPZqw1HN4bWeD5gh5CNiyYIbGR+rbFySDTuuQQhnTA6pGv
zNHkBPma0UBheeHnv/thxbI7KdgIaWWQCFpAyK6EW8Ecx3o1SZBXEpYUu4FI7RmryfxPVK4iD45K
eDsL4dmJjeTK7eicHoA3egI5GwgbmMbGeCkMEioXwK9XL6DujDmRssmjUAL+DqYBXyUc+siwCRvE
dsiICn1M/xFt2nLkkLHvpp+6TRn9NcuHF1/kw8HnClQaWBX+5XC/PIMG/Varz4QuoIMCSkakNZuZ
LyUXPKQguWecTttN4BZtf+yVdTg0+YR1CYFR/MG4TcFINGIFlgaser/VtWugZfoYxrKtOOhvMEXU
DFiLXg1qAnWpoEJ0Va+ISh5i+DD3OPsH2Wfg2FDEi3SE/oJ4a/NXMpr9CCMrjo2PFTmR8c5sPa4x
5wy8/lspbvgFujnCComI3osjJrBuEegfYvcoUv0ZQpZvRyQJPUkgWOvuhFWz7e/vbI1+k5pSs0R7
ejNAJLEyH8f4hy1Z+WTiWlmjb7xWBGs+LnSzXiZldtZkMT4GJHp6qQvWQ/9T68izEWnrljLKAniA
BWpVvV/lRgLo6a7mB+VRuO6ZTegz5YUv2QO8D8FXvfAgdpTgY1rFOep0PQ3KtqPjfyaADXDpLZrE
7iDLhr4V2juEO4NNIwDNGV6e7NWgUhRCusCw4AxfB5UHB4Rs8mFzaXeap+7vudOLPSP95zAISM4v
G38YfF5vzzYKO5/x6X6spwHzfLw+3hgGdwTd0PUWvxAuDZq/z516ej40IqhUJnrp2fYh5KraWzj/
ARYpC9qqNg8hhGe0qgjV5jZZU5Vx+mJxrzCaNRo5rjFyJcnmaqRh3EwbgPs/tkgYxRpAh2utRQq6
Y2u+kHSkgheXpUKZnia1g0coul9kgueb7F/acJ4nJvP14XJTaNE9lBKOH5Cn2+kXScPuzjhvaKB0
aq/UUG6BeChlZcp6gz0jQfmQGVuaol2E8YwDhgIM+UUWBOdilJZS8JXLP1KebHJ+g6phLiRdqMpH
nSIJYKyFvk5qyo7be2ia4T/x5B7mhGVZjc19Y0V7DHw6O8GRUIIouYS5MVxFnwczcr+6Ypi7I0OK
Y3tB6Z2wtELCWMNQ0UpEpRjDXXZR9+aBd6SAE9UScVefQTHdxcqtwlO3z5BO9IKvxdzGbe2nhQH7
O+EozwcP0RNrY1W22GrC0QOyTZLD3M2D1v76h6uArMqYY44n0AelOprnLss/3UqX0ILb9d6Wz5GG
IhqQBuGwaBO34iCbfKqm7DFGyKZBCjs8zthexYGQAGSyUb3igZXreW8reMjs5i/jUF8SQL8UAtZU
+HimIn25e4/spNK6fNfau0WGfiq6UoDMK01ZIO1I76TjvxvutU2YojujujSXgJisPvmsV4sJdyLX
3cxZIZEYXh0+iGiRsYqEmtdx+URKCdCPbbAiRm0bALItRPUM2RpUPFJJKOHkYSAriRTgLlmMoYVy
KobzD4zbOGkLPzA52RFhspYs0EktiaCy6HxaktpfXWmIvZJleKQbLmhUNcm1mw5xDa2CjzDMQEfy
/Iv4Wj/zOvGkb2X3Cok040l8TTCdqdBtAS2+vGSLq1JZAa0XzxZIRgQRNlnrfy9nDXmD5jeRvOlE
5MmkNzO+OWyNaYKz+66Apcpexkjm/pWWqwQyGIhlYgutXCZ4z8rO7AsO6fNonK9g3T+GxL7Ynt2k
MSBIsHVautiyO/v5IiXV1fj55YqUY5AvjGDT7Gdifn/A+hn72wTAFFaM73oFu/uuC/rXoE+CHSiv
SUNG2EJFfQe1+w25YTm5jLQjS+zq+99gTveC494ZM+egVQ2GFT1cbUDSlhi/p+6p9NLky3giAocG
MndHSePzoXvPi41l7lQU3D8PCEKQsspv1wcmZkfAz5w5BtNoZLpilUis717DmqZDZWOBMml88w1K
qauPfNRt08nPSGLNhQQiQjaTf8C2Ax/uX4MsXN3UPUAm0P+CD0bvTJ6yOWY/3jULAMxLUHAaeGif
/gkTReyK2a8c6jHBy5YbhG4iVfC7YaxFCdUOd9/tOTGc6SoT8x6t4sGFAFw1wVJ5DyTE6PZWMxU9
DEIkHfelqawHhNZEwoNSAFLY3aDWvXIKEVjTkZQJ5mvq/p5xogrbROX1A6QzU17ZXsYoJzq1mjOx
Uz7RlaEnprNpspq0Ni1lkTJIivz1b8DGSO2Suos0WbcdiupNwnc0+YCuzNBCzpx3+SJA4Zgp7luO
h++yTKAO7Z1GRQ6GPSJF0OYFXYh7X50eDhRS6uRQzsPip5hLGD+lPJB3NJoDvu7Yzuk0Z86rMYFg
wyNMyJouvRLgZHNwzl164kzqWTROv+WN2tMqtUvVWCqGIS10HKVJ48IautHrrm/6uQoyn2czU3KM
+zCt0wj6TCvz8NK+Ke9Z7lcNsxqp8IvejYjHYqVc8TuzNqFf5+hB/Q7JnnEktgTaVpUBv8dSqpMU
EGr4I+LsJ/ZGl4OJb+svMv6jvM55H8/CP+3doYBkTYqshbVYaidAoZbZCRgKhRZvqWL7D+XyddXY
JFUiEN37dZVGgEAXk/m4kTZqXmdPaIgaM9smIMaRFoK7JHgXvpuR9bEYcAAg+RgXONO2vnohxOqM
xIvjUTHU4/RqeggHQ+okAZEuDSpUSHGvWU5kXJvFDIl8qVO0JJq3mJJidVa75tyNmPseAD7rn3uU
MzspQ8zTvYY4yBO2uDF6UlPHyMiFYmQ16ygJLM/hNACnsMszeX2sFJ2j2gnMV04ALp5ApNVXm2k/
PYQ73pZc2RdSK8G6JlhigoHU3N3ciWMA2o7gEU0PdFf0BLSSzc5H9iY3Dg3Dn642Q675lAOaQDUu
hzhZRVptkVNX3v/OMeemlzXZb+JDHdMb8FQ9ZXlJCC3G+jQpqQvHJHFsuNybaiZeInsjAkKh3WJ/
VuBXeQLtCmJZt4RygmplVv0gVScnmDad1DiGBCWPB4V3Eu0jw+T7iJ/pGQfR3WrJkpyKoKjxu06u
EABhmnRxWgIESQjuoXHebsj6Pz5ARXHofr+dDqDGoB4Edx7habCbOrAFWpPls4NWKVQ/qmqwy4rF
9Ya6ET6J/DQTnE6IDzgtChzWWRNYqawDxLI61jrA0erNiy4ijB0opALwVRLaTBLRx0R1cd2/T5kw
i+6Hvf85t18WCcBP7XFEVzVAPvcnIh9GIsQuvp1VHs4KCbMt6kqA53DbsoV6GszrYWuTBAzse9Qb
+RYcazGH9nZwSsffJ/nK9J49NQ5b8O1+pYydhA+KuD7k88aXShQNYg/zOKndOhLCtkv/XfgFhNAI
UpM+24xWIpRiDNpXSk5zMlZ1Nk9F4WXHfVcs3W80wtJytHblfUM6qq6pJuZzOfp+u0j89ecgxVTy
n5g91tvFnuvR9oMZRRVF2gLr1xymj87WMkOoeibVYygrWKCVi1ULfvdl/Xjj2JAusy0gPvVCgCpt
PUm1w5dzfBaZd0Gp6WeSPN6qr4ON8cZmojslHYp5RMs/4KD3bRq5xQBwTn2Xbu5LOWUdh/jYytS8
KMi6eojxmxLI5iBTND7ESz1SeF/1ZMrX9hFo6zLPB4Qw8ex4b3LWrFHfxaOvQopobZRRd35eEZjf
VGSjmXmrc1n8GMS9ne9lR8Z9rDlPHJgyOT5mNfPuV7NFGwrIPALymm2zIQZwGiBgRD8IC5ls66wU
JOyzJym9zcaAl1tQQSXVcH2Z5n2MAcvTGr0IoGohtox9XswC4fX8w75c9HUEIBcaPhC8LMTl8gTY
qUM8gjDp+83QLXa/DILcqwoNBLlOaBWWFfEFANjCVBjhw4dsuciX38Kemin4Q+oodLNYEB78SfNE
TWqEv8GFkQfrDpsP/gT3ws4Ttwq8AyAbdfaxLZlhCUcmYgLl1JESvnCSuPTMrryZvMxUZrSPI+Tt
xiEgkwmp6WyZpzPx2RiNhsqma5JMLPL6p/lpTz/wyTTIZ0KGP2GiiofqW9PvfTA5BZcdiaDYiCDB
QeTUihAY5ps7JzRcBwOOkihKonlCaC/wVyslUkxVdWkXcXlbTZWPaM0MpL1pymbYCjcEYB32geeo
MmxgKqNIZv9lXP4joy7nM2DXTpcv0c0XsS99GCnGl13Dsl7xIaua2t6fiin9ilHTtHAxpmAz04sz
T7z36g1Aqk6wgFzerCwP2yKN81oXhHRT0N1Zq/IuX5GiOfJA0qzzg7kazZGC9kYEYFw9hLbnq+rW
7gClghxjp8esTyfIjxxg3CbgR0i+UyhmjOu6gddjytuz7T/m6kkkFOs8YvG7uy10TTienLsuos9u
GKAWdxDtjZQQRRrlmHBI/WCZVBadc+o3OrTBcYPRLwe00W8dUadYXjhpT7knTM3y7GCvlDTHCc+P
TH5/aKbQEbOyfbHlvCkXv9wa5i+9fkoPHp4ucjcS8Xp0emVrX1KgMfidjqkpD4DRoM+r0wedYpDJ
jHMrsmu49X+mKbdu7q/w1m8wNCJeqXqYqmQZi3Wkkgdp6W6Twy741thCKxDbX9jxelCpWWjkyVZs
oD7vaqR267xc0/7bNmByfXW6DxkjyrB/db+LqJuBeP6iezTnVnh0RoUSEOhgZvQxETw8meKJy/9a
o2yH4gWA/TEmzouecc0Z0VxZCq2iujwVpmbQGQk7ls9jEFanA5HYGOcoZYddMFSCr6tA/xeY/hR7
VbBvDdVAzOMRCMqhbYrBhSDQyJrnYP5ULHcXSFoZ10L0N0TrnYp3Jr6eFa9sN8EmCtfA31uCiDvV
zIsQZAnzwME2tXEtX2dSH2n+NFmTd69xRa1UY7U4UMjCezvvC0CInWOvkPZyoAeDvWa6ZU0phUd4
0h0oqyL/kQM6sxwVZ/jmy5MWBt7tmk8s5rxJdRI65FqihW5Hv4feMX47AynUpX59uMrlfNjnOusW
iI0LRMEmUqt1LlM0pJBxLVHc/W1CDWbEoyt6OJDCR68k/RVNleWz+NPmCHKLitJLe7NXoAbHrm5t
Y5t0fxN9wVCqOM/AoxgEIRODYETLmaWtpUAXLkRxH+VhKFOu9HUOUApQsUHKY/t2JZ2IkXKurXD/
WtVt/tIrCSZVJ1QcWfaDc6C3xLpyOZF3V7jqA8085QG/S4ldDLVTB2NAas2rJICzrXhJzzKghj62
QFvAAAv2r8pht4DJF0b3LsIBsKxTMaWXJTd9VgQ/s8KuOpNsWeuEVCBVQqb0y/q4+sMgE8qJdDqa
UwIMGlmsnfRvdbQ++pVV8nucBTw+0lkBCYDcizcOUmjsvMGdV9tvZ8t2XO1qdsRWR8BulFUW+U/j
aLv3LLYDHhwfhqkKmo+Jnoy3VSIVaDJeGWzUXkQCTDd1rW+6dHi1LkH+jopU/6vMiV4+68hu7KvS
uc+WWcBwakx6o481I/FvuAIc3+ksgbHOKPUsvPbE2y7fYG/w6IYU+DuHpiFq26G7kLVUlWuKq0Fg
B8py7hYneqnsQN5aGNL+ZLdMaOPqgDHwhIKxNf0O0z7yy1D6E2BIYQ87vj7w6T2E/8epbUAE6imZ
SgXuZJkMPTPExvVOGWVmvJ++TjnuReUcXCddsiRAuZ/JF9oSrN8d+tCKYaTn9dCVFr58wM+bH2U5
dFaOxd9a4UKF7V8jyDKNQ4IYEBikV8b3NAkV6aYoMBrocsBnKoqD0HSvxthDwSpAgQXdeYGNNitR
vs46F00P/3Y5vUgNGokh10ddYuuPI+gdMeT1J82YNT0vGZcgjFPA4RMi2NDfceiL+miM1XKHk1Va
Uano2Odc0qsQdlDd9z8nWfKw8nVrGYnADu3zuC00pce1dnJec25amhnizc4KwWxfa5U+PekxjBQR
c1rGA9pIcUZkjBHqDkxAMsX9s2WgiQYrTJbR+VlAUSrGGDtsGJHZSvr5D8CjCEHlMMKF7U6u2t8w
fl/hwsMpECny9JDRnPb8+UyTfznfKp1PmqRO91dVsrJDON005wWaPJZeeP9gJwJY0muhwruYRnxO
nuCBoRZXaCdjChClQbDX9BbvVm49/0eeEWA4I6zqoAvIXbzT5zyrPM7mYI+n7J/lgbkeEcps9ZaZ
x5ayCvAbB9tsuWs8D+5wQBC5eIj3WRGedKihzaecuIEH5Y0JBHcYcqOQQ8ydxFDHUiSl5jIaNSmj
EZbWb8lF8W7o/IJAsP9VU2lDIVKnMLzCeOJ5/eQh/58AUsdSrEsl1xmTDUtyWUzTKEY4EAJt2gGO
9PBbvF6crBSEgkMQyLgGTAh7FPIJ5rMJ3oHHEAwwWX4xncdmD6sV7jP1yVatj4yhZz59SgjL8ZP7
O9qRTRHhq+MG81NWwmrXY0qiE/5Xi0hki5h8DZvLbX74ZbY1BAJAkI9/bVOQxZ+vHqR48UHztJOY
rBMjlGZiiS+YqModX2mabIrrK6TDUrCSnd/Cjegu5iavVaLPgLsuK8fS8ZNRVWPOGfXdnC7b9N9M
tMX2Jo4nixdNtN2DE7PrXEYbY+R+nLqTYn6SEpCC4nrTp13ZJEVEmzzq34U3MQWCvtJH2Yn0gsMf
g0Od8wtUJUcIY4UrOR+ut7n+pOtAZdVRAv1qfEMHCJ5EQFYvE9vSdiaMSZyeQWgasCxrvNcCidmx
KS/Co8sejM3uNt6gZPk0C7TNbAinOSa5lwuoaVV2+ZSUPaKTKy+h9/dL+rDiBLnot+VYLQ0I/xxS
Q4hjGIJzTMK+BDZE6rKiUqUxYscFmrpFeWGrEsSVQkOdJk6PEdVk4AgxD8HDFtFCtqnRz40GvR+p
dpMyQsFzwGGCdnd5sXxfbZh0uv5y2QH2/5A333diahQ+F7tn7K2v0ZHmNKecCQu1QfamH6r9qOin
Igrpczt3iQQd1EI76yteCjs5Kok4bkG4kJ8uiz83HcUDrnbClU+SX16C42zNiET8RcLX1HoqxY9/
ixK1UGCEg6EDJw8KQdvf8HWGvR9dEFT2M5APgQUJkZeqGbSuhPLp36s1guEzX59/ovJH/WUbqMLJ
YS9EjFNGlGKojkCWv41NUmIwtd0ZjHN6C+G+xXD8ZPvORXTduiFHiMGYMHr8cxfKqbFcAiimNNE4
O2GI0KmuKVknf0w0GdqYZTqGE+ZhDJfX0n9vJX+VIF526KvibGxpQo96rsVkYRUNEvAfG2prnOun
Ubg+9126nzHaFuglB4OhAbmg61JB0YjEJbs1XeJu6Q/H8ZiAtpSj9AQTkIB+r3yi/5JeCb+TTi4U
2m6Qxd1DIyd1QsYmYzprA2UWjrF6Qb0wO1WeKUb992ZVSSUCKDYUnMtx3Dq2cp5rGH0nkYd4Wb5j
MVy7a2aGViJbxjYNCuY6GoEFNV7hGw4w3mHxk9m8d79RPiOArptOJ1vw8PWXr+XO51DsZ9uRf5di
KUvs6fytht8GkZBufOwdknewcsUm4bFT2QvskGoGN5iWxWXlv5mXU+R8SX2rkRqtCdAoqg4dl1D1
UNR1JCmw8Ej2+rYLkLZu6L/+Ran0OMuuhTeie+kdkFzlVHfaM7Ety1QWWJ8i3wcBqK7YfLARwZIc
crc9rWrGPWtdGSCRiop4AfqKg9ENntgx2A6aFcCojVMABU6zxh+PRVzkUe1cPbDPY53cpDP9U11v
l//wgiDaG47AJTbP7vbw9EE0RvZZMrok2rSwfb5h4XimRA9/r856gQkAr85OEBOsiq9B/FVQBQrf
1hoKvgnCyaxsRrBI/lCE+h1n2ygp7HEq3zdd7QU+Uy+uftunUsirkb8T4O3E0RV93fJmzP+jblwZ
lv0PaRtRz8nE4wSKWyHahO4DcNQdUfcUnCVp0rbvrtdz2vX9XysS3QSjutoK1bcFu9+AkIWzw1lp
TJhhDsZlODE5QP7RzCRslxn2MoY0qWLEq5iOKQ6P/FCVI+L23eXFjrTVvSz3zIEuNOI11+Xm4dKh
UpIo2/vjVOdolj59rrO1+EX3rYeocQZ50aqdFEUrK7WPsJ2z4KZdzmV6klqDFY1lruhONeuR9AY7
Npc0spIDkdL2bodboNxjMEqs6s75qJFjxnOtrsk95eKxBuoXs0XVIA/qvXieO9b8lYWAQT2LhtXg
qUtrpH3yHQ+KExHsxGSMWhzA0ic3D/JWPzgo2qGVjdbx2vWqeXGQbfLpSLQBRkNkQUeVeRN9KZkE
lHYBeKY9ZsvCofRZ2N9DAjFs0LSTVLEQIvt5opGHkrcH8Cbm+36onRpKjjDDx8pOU1K9VrzxSxvJ
WenVrADGM/CqlqxM7jNOxJiMYe/aB4FsjnM9Zood142Zeb23zfvCW1EudTFLOqFIPdDkm0WyLj+U
HZzb92kn5gi+E/gHvGaBxgue90aGc+xJWhq3XXb4GlewU0Mo03TEXVS3h68tXAk/ujz4vx58Z09x
RIno+Y6n+sCKR8hVmO8ldwr9HgGt7gA5kU61ihJmvMqO9GwZ4fUlb3ZKpLe2ahKicvho12kSmzi2
wl7NADlDVzgE4RWcb21ni2gtX5LUcXeyyNUcwErKiR69F3SVSd5RX+AiZ3TO2xhtDAD0Ofcj+3sc
Gq2OxIZTjftipRVc7lZGz9oR19J76qA0fUrASrcwiFIRU7NvGqbKIhBCsCYG3TP/hx04NYXU1DRH
mbjRGIcmb184HKqZ3rW55jPzGddl5hnrJhxC8aqKtiCaK6a9873LmgHXFNHb/K2Ot7H33pO+eEoi
JGL6HxjS6jqyTNfLwVNRzjH8+Bjo+2+rEM/rmtAh8cWHmM/NNi6S6+tIXM6UVX1JzAOtyASx9sfi
c+j3R7BOUdgkRG+YszR4Qz583bxL8WkuVX2JI7O0CD8nsdGousnb/TOul7drOOwMeVWdiq9Zj+F4
oe9+d/jP/ipuqwzew2YpUCY16/idOaDmzv3LgwIAmpzknb7dj/Yr3otg6/buDyiWEl7x0/Ff15Ed
9S+hY828oMrABiN/fiRLoDJI3FkPnaZFgkC+cZ4oisEL5zq4s+OWLzM2+sqoh/S0RLhrtrs6Chs9
OGAnvfdWDWKT7j64V3l/dBNIzqZSmU/vGDs0vffIWRhQtij9ni8DbPn/mI+G9T2P067YrZJxJPiD
asMoyM7W8ElYVPww/PwMSVoGPPLA5ULslTHPa1G8DnJZaKKTejGVCKUwYjwOnoh8nv9brqI/UgNH
Jw7e+Ysus5l3y6XOMwc9nb2+5bdVRUu+tyQ/hTZbxLfh4Z0sUlbR5mO5I/b4yjsGCwxMrjg2/Nef
MxJuQq2nxAgEzayT9GBUAVcga1uUcPKRZfZ73ZYHfvutalpPsFSlnoWl+xGp9tyFqWKBdoVlTBgN
VeYDsz0qYubLJnBQ5W6ShEXCKGGRRjvKz5n34I5so7p3/eKOcQ2eqXPGyhSM3xr56DlPdNb2S2Lk
fC4+VIfa5vj3jYOOLfraiOQyXvwsxM6EduR8VesklhIUnm3YZMnFcHFeOm/jIQPfYAanRt0CHHj6
idRQeen816aKYtEfmcFmzBF2V8a45R1yvCd3b9O13mvolTMPFwfmNECd3xJcj2wcFH9sltBOrfxb
9tu9kaGtuek16KdRZaYW3BIC26Sebt7MJOl6erx6kWU3BTExyAywtrgKdq0v8aajUw5Cqi4+hVpk
iJVmNPE4rNJosKdr/B1RYpRgR9mvVHg43VBSJeeaj3Mc3/RUXGUKi+Us2seP6L+RvImEMaDdqn8u
/+ps1q4nY20tPfKs41l+bBBTcCGRjxg+rAX3MzMj7WxiCJXOJBmGAiDJbYzTnxHMG2puhmfuafGl
ItB2g5gUDladxaT9BNRE8yNDEUphwfna09QobzcLF2sLgeCJIRWz0U76vclUgcyNxanW0XZ9uEEq
QUdFgwSRKl+8IFBCzNSjxA7xRfIzq94X5HFdWWP8cmZy8LUusfsEJgR4yzfv5okyWNbmg4VNpWrY
vM08ksNRg09hzuMVhTKcQOGQ/fG3LHE/2gMFzxqdKb1yfA/alFgnWYhkWiyVTeHv1eKEmlFHjM2j
OIUtg2dBytZ4gJ/FQeFqQ8Jw+LkeRT0qsPmLMHRNTd4Mj+8kGtQo8FJ1GoSRTQPNBqw28pCC0hqP
Ew2CJ1HVggkiwA1Fl4nUy0F39dFB4N3VTEOib7zZ7C78XNHgki6xjcqtFUX1m2iHjNAQbyX2B1DT
XZ7m+Vv5bASh4SKsPR/qaI8L5o2WaNb5WC6gTE4U5rs1RzVW06GYkYQ7fvTZHL6+yMFlU6BrRziI
gOMBlmDDGja+oQLb+BavelEvQA2a+V/gySz2oeccv5Yat62kj0IJlQimcHhv+aGx1gojIY9U/A8X
rBSpnOOLWD79qDlwLOD831UwyQH/JmpHMS531YV3gEa0lK+bZqqBUK1sUL+/O2ihVyx3erm0ki/1
YCMQMOXsgd0w6C270LaQ9DIq5JKqn+KmhqYCdp8UUyw5+usHKce7idzk79fllbh4lbyEcHSKMWI7
i7jdF0HvTDpMa7uCvIvIye5e/mEa5A4em7Si8P3fw1swqEqaC6Ci3pmXOu3Y21XkqqTEI5poQ597
WTaZVDvNuP+dKkW1xf9+7l0p7nsOpcf2YduxTS4I+41QUuTFpcYStiA/q8HRXKXS95bMX6g1kNTi
pKczskU8o6F6uhjpT+j4RUIjfLjU4WzSC+xF0PGoHfXnT3I/w7mnf5De0lxrOJzLtDXBQEchc7GX
oUxnv73BQZrmS+d6b+CctN/goPLKIqz7ExhsXKNNerR3NXKGxRmvMsoX7Apf06n42Rh74kWChOqW
ALWoCNpQVNb0Be3BgmoLWGm634MhBnpz4Lci7stIC5vjnOSurzaJLG4WBUZSz8JSAkUPQfCSJ7D6
2lzeQ3EN9u1PhcwneZaWy/D2xVACtrNE9osf5kuOymOGt8bFyXvb8WayC3rsTXi0gxG/JqiiIXfy
0e5onYkN9yzWPhvLQ6uF0AJCUn9r0j6pem/SfWuoVWj6dAdm83vp9aK8/Z/dj2oX54QBZRqNdFxZ
zR2VxQmupvLPeo25wqhWU2TmUAbDRivHNyOVItrwvX8Lfd+D4QxjQZ1FlHU5OM07ycIJP686S4Qo
6glgD5dY29CPy7y+7MT1a36ADfgjCiBk5d+BFwbPYNhWDW9GQmyHbvmyKvJINlRjcKYKrc2OcZxa
tE6sxrXO7oHWOW33DTFw8Wl/f5+abqYsPNssgHclmDp5TQLkMFg6B/PocFLMlkf+RBVdEuKwf9FO
0MqWNBC91Ox21NEMgTebZWeu+RIObIstF5iQH6QOxetjq1/kuYFQ42BLL3wUJGyrQXbtIRLCuzzq
sluwk3xC07pLeP0LVUjeNe64Fx/A8GWXU/8gLlt7Zz034iRM8qB84MdDP0DJ7d2M30yomK6vAj8N
ac++nMRiLVXejX57r69p+yTs7OtfKJYVbdn/KuxO15JsCiIct1iJuxBdzyoK+5sBbc1KTAbOtSm/
U6PrvGqj6tb/+KgnpHaQOV4/urBachr9vJbsS/BM/fiqRVBCQ/2OtdPjnjqueSGqGdvBdduP18CU
cn/DC61oo3YGctWth4212m9YGXW3UYSZj5mv7jsOJPFdsbvs2z95+Odv4u6bvB4TDZwUuZOKD9Rr
TEZJbFVUar8AHkpp73WXdOeOPVa2vEt0HhQ+igwRcwl6U64qeyvj4S13GbZ39p3yzfagsBNOpsjV
xSkTYHy8Kk+WNbEOdNyCA95v5xZuBPn4BwBmxxOBVWXwUI2M8Tsj77gTar1d8grVy8zNO72BB8/m
uSHxyXDy7mPO5mCoEa35o3hHaTsWgWImLKenhQqJVv1ypXUXigU036Rk9LouTAuHgJwmSCJBYf0O
k+CBC125WBZfsP/lMYKW033zrfK3PifHZwdqELHsoYa8++I05dO+OusLsnHFfKRIVXye+CoRdE/2
bQqHYXsKp9xUQjmzEV2wnF3phHhXhPXdAycAGaRb3ZzEil2iA2KGy8Njm9Dl1sEEPkRcZVoSpiBF
7WHGVtQq7UzUTgYQFB3oXMWGt8X9k3NveZ2oEzIACAZTPWUWG2mSRSPBTqT8wll+O6KbgZ6PiHuY
dWht/owlUFoHiM5lT6UPfgz9ks1sdeMGBWyPP13vdzkiNumRabrvhVucN73jSFQ0uoz/GgwpPIQ3
6RYTU7VgvwFmq3Bddefg5PUfFbBkMgv7wAN9/vbKHkR29R2pjz4q9qXjf17j463ragL+b06gPMbv
N27BArue7ta7wN70kOcKdQF9e83o7Zv+bV/IhZgzH3VZtYOVjrstW+X3NzyDMV1Z9fN92Vznt7nR
YI2lKcDYOpO+P6e73f/OgIQOLa2GfQK7VlMFqqbJb3iNetmPTx3ZYUqhpGec42VzHfLsuepz7R5I
5u6DILSdrTK/jFceN8Rj2azLp6WCC8fpVdnC7YW6kqIQNzvoUUO+Qm9f60aqr9RqLwAraot/h+v2
hsZVxlTScd7MhZyysrZTntMITtqB2IP1HSOxfXUD1CUmKJFDpEaxFOJkHdCK9QOX4mmm/mKBQevG
bDbwVaFW5EnRNdUuXeIxgP/Y6Rt9cDehB2e0JGnNIy4iZZ4wzgeOHnT+rLg515v/1sG/ZoU6uwqJ
wQ7+Ei725Roda8WnH31KUjKoks85tmGan8mWyEb9uhNQMpbTC0CGWeurFhmmQpjorpQ+q8DWubfP
gpkL2Q0uM3K1MkVUiPNIl5qABlrgjXq6m6yiAXvHp1+Da8n9ZokP9VvQ81gpBn1Dv/oBPkBdX4+2
MrK/e4OLER8/dbCEglfTbX1vsaMeuhfZjDgi7teC43H6XWzmkLdGvN3mr7Dpi3PfBpqlFSrPCzD2
yuUng1I7ULZjuA/TzabPt/TSnEjL7cV+jV9zfHAPoj6W+JVps3otj0i0zbKNfNBQq+tJQRqKZf/w
IZ4uNlkceKbhdhA7KimCy5mFlonfzhwGjlgepuMq63Wq7PfxLqlGoA5UYrXE98jFcSZmlP5ylMVs
MFAH2jr8QLIEzl0GLgtQffOpBjy6J+VLbvYuUX4lbpHmSeaG1KOjmbQWa962pAnFrYoFd+8HG+DR
XTDtmWM04SwQZoU6nIQ5Bgu+6a888sMtZV7XRChU9z5mfU5eRPoQCNe7n1CGqDurY0qmRK1k4Gt+
MOsqExlCM9NymY8wvw7E2TS7sIQUUw3c41ZBP2KuY4Resfugl3BMpu5dlXQioh+U9G+2BwloK/EV
Pf0YM51wvYD7OJDSffkF6k15J/+D4Y3E2BYkVfKAkmHYs47BSNbk2jQG+khnVAcYvMgKpjkBtarb
2x1SkeAeqb4FyHew1xrE62WqQ2jf0WU58ee/gsJt0StKOm+umYkDH7S7HYgGagPR9nXZhnFVg1/0
zZrDFMRJA9SVzTe4Ep2EaxnQDcfKRQk7151iIy16RuKaQCg5Zl5tZGqxu3IzLPJGeEFb6OgLiM4S
gC4W0JtxNKees1PhbLOuKG5DJfqR6p40ofsHbobU7l0dgxxN/IO+kAkOQJPkcU24l69JPeWApFxR
4CD5omyL2O8UToIfYzP7n9B32nnJEcEzgxLPsybphtM3ceu1bN6pDbsBia4ljtgFJTeRHoV1R/pp
c0A2luvCYzR+NWLf+MwMzXXutS9dAqjuAcNsnqbHR21l79xWx4M+1VhdvpIphA0pmaeH23Z4UonO
Xzt9u/NVnC/Ban6u3J8Z+C2MdSH6hxndy3VDmoIYG5G5YP9f6ri6URIVK9WApcL4evzcICvNwhP7
/CZDlAhdxG7msSBkIlWgEf37NtQFFiAkb7m6NECLa8BY73zW5ssX6JbiNjXpFxpm+IWRWlRCmyEU
SrLelX7ovoQPvLEWU4CUoB9pjVvWmIWyrxeDCHCD0O+MiXhbaIIkSaDlMRG656YdzIQDW9GbXyTl
Cvr5jPowC3DAyBB8qdnNcBCYZUu5Y4pm6tZ9ZqVaOwXSwFNoYNL3o6VW3neK0wmxDov67KERnMQF
kv6DO2T39CoFsz3Ryqc4PpY3eWQ2lsQD4U2HOgBamkxcs0QjQmSbADHARwpedW1MfB4AvNTHAh1v
JbMf2NRMXHOenVc9YnL1en0jmwzjCkBjdCDkm97hi5c/bvLmk+izlEl3xTWC8OqDOo2t9eKMrSU2
kRw9NxnpI6WuuK2pmHpd69Gzn+RmfXLpC64pQYi8y5X7bqbm09cjCoJt7jHFkfxk55ATki1foRd5
fmZmyWvbsnZ8SGVtSZBfifSMeQjUZD+qy6RdoUyexBDIFFOv6GiyS9qHRmC6vB+F/sQL0A+dqpEU
8TRVKecmUbdcLBZ2IWi+Dirphi/CEUjF5MPwUELr5MzJOsnvTdMKNtuXQzPJZdOnLippha1sgWmQ
LjDoZyk1eF812E9UwmfUkygVyJNydj12M2IDtYZ98RQn/9KAZdnB/CLs7mWZpHKxzN50Je/G4l+i
RAvUgASvLV1/+iMr+Vj80sxfqjzSVTPNeE0KV9vfW0dvMygUWXcSBBLrJdgUIHXUun5RZSRC4Ow/
o83Fk4g39T+xhvxtB0ZkvP4NoMm8RCgUdhLnNw+csHMyQV/+9+ftFZqT81lePQCqnbXOMIkN+1ZY
KS8nxM/XiwVxuE1mOT/PuxqyjxZFQ4B2gZngukBMLNw+TJZhPTfX/jSYT9wKIaO0plbzL0wOM6p0
aKaYt1CWSjAgbARyZ9OQLhTzghuh+FAyzYvszh5CjPC76wWmwvTXgzDOWplbmClxq6SIg/57LJAM
hkQXJRNfQTbHxjQm74+sLmo6h27bhaLh7KLG+3LD1DrmkQF97504vgmPC0rBpYGpfw/yFoWwu3Mb
Y6ql+8VC5hApiTAz3C8tCgvoL2dwzRyaJKlR5oadxemFUi3AaqiriPubWysDBbdOWrWwohPfpB2A
j2WDAzRMZU/xNqKdJRtmPut2g4hQJcFtxvICF7SVV9N5q9GVkr1tzzydV9inR4R/7YxhGCsF6XRw
4Ruls2LNi39V1najglmTfdSLfBwj1aEtW2kVwYhb8UYROz7R5dHkJdZMwmoM7jO0pEBcMLZ4SYID
l8uZbA7wA/FIkZ8Lrf5uZQCmDOy4ByyzD0ivOHeeJkcYHG+RR2Z4HT8ASp0GyzNwzkf/T9ccyaEO
nP4raSEsSNBtXTBnTrdcvjGBXkjmpph3M7/ULejt15yQn2g5v2ffWrVEx/G/bRa0YEmCt0UU8MlV
ebC4JZRNQmNXnHTqdihsTPsW6IBTFe04ZUsho3o4SMr3uKu1O3jg84nK2tqG6LspuZrej45HetaO
b3RlugNuGRU9AU9wum/1mE1IYNstmIVtigShKbPrq1YE+HgKheqc6OAeDlwdVvPzXb8CjoudzdKZ
mrCK9ZxKIZ4P/Gz1d5E5zWcVJpYYhdawwTkELzm4P53yANzCbfMKXr8TwDeWcx2lTIrx9Ku/nqpQ
/InhMEPhuy9wYBKtfY5V49DeniYQSYxjppHhiVKQD3Z9CKyNkeZJ+P9OrvQHmruXFzCeXFetMSe9
uUI8h/QYMJD8aKlzUmc6L3nG5nIiNGNpcvEqqE4CzAIXhO/UUT7qusTgh279KFxZU9al5gJdzSMq
kf3NVhQ7v2Z2fHcrBtHsi87ATdQ6qLwnHwCCN6YrLYvWPNKOTxnmgl4FblFbll3PHAMpReEw1VVe
BQ1yt90ze1bK8HnHEAY5CY/GLdMK+DVmTb9mbGsxdRWMCrjrivz+jBH7gSfcbSKgzorpM59luAyo
aqVwD209+vCQSpX15XnuUBVgDuFwQjuHL+jiOZcvnUaIfxdHerS7/y1ncN2jpA/Nm4AYoWQPLcDc
Svnw+qBKMBpEj6Tk3v338S7alOEytJmBIkpjUpJRLQTOnIkqwa1VudK+xv3qtNet41oYX7lHNMXC
6F/6LhPJnm2p+L6qNP6R9/134jNIUYqnxkzvwHJ4HVB6g6B8jkbaIGHSR6J+xzjsK0yacw8SVVk3
BmluHPCyDdpTtaj6OHZ/qPJpnWi1LyiMYDZJB8u85rOq2Ea95/e0G0qAYe2wU5KUHE0IOAGyJPCS
Y/JrDulc590Rnr034jAGDgA29tEvQSFClM0q3qpVCYheSavF/2Q7uHtZjDQ4paFFXNfB3dvqfjsz
PWdfKwQFrTPe6m392MlCHFYshrZ0LSBKwCB0E7gGEKzvM9ayDRfKWDwpmi8N0PkkceSR6KG7Uc5C
FVxfTI3OYG1lyFB5s181Y/SfVP2peD9cilv49lWo9nHqQ5klihu9I4MPIQlrh7ExohquJTG49mN1
GTUkjlCigJ7I27EYAUYOFnyueWfjb/5iMlQuaUAd3f97TSpnhL6nYjrTjTwskLF3sqoECchT9zQy
mMGVO/6cw6SKsbLM0oi9bqmrOytpXl84BXpaKxj8XOTf/0oZcuvsvY3o2Hzs4Cf1IXiox+lLKbxe
vYHJrAX6XmBYmiraxR2vQkgNFl5sJtNFoRJM1GB0E7O/yBD/vmQdBDhcuXHLSwM6pgnHbq3sP3SI
U6VFcMSmTi9k3Mgf6lzY5SOo+MU5Qm9Q3PTErybWBfF3g41LsOgkAH3nnzRL/QIb/LAC9OqqygBX
9+MTlbUlPFewRt6jNIEIq2Y3gSSvhqzdNtUIaoejlc4HhQQfnIBcEdD1yNCMm4BPcNVJ4IJOFQFP
bfF/sqiDQXUYyuKk67YQj8m5+dwqk48LYleZ6PGcvuwEQc57yZWL14ewmGVQExxSluyVACSBZmwA
IxqETpc54nvGQNdT3gxxPUO8FEKeDZypG1xhBpxer77yVKWCmAhrRZdjhc6epXf69pFB1W8rW0gx
hUHlGdbGS9NHMqqn3jmFRGzr51KuyYK8yPeEkeOspvOGV+XEq98i6TA9RQjyDu8LgdvGpe9w/eCF
qS1NAwIsW+E2giTukBKfnUhAb3vQG34LMK3q5nszISsgfhqxhnAXcQYv0h90OVqTmQKP52s4ZqCv
iAuWmg0lk5AHF3UoJEDkZ2lx93DOICanQS7GsdMY3n8R0e5TuVuQ1cdYyI6Eb5V5La7WF0yeUKCv
8BsjNJfzNOz6jzsg14VRNWasFKFJTHhk2Qr2SLXYXXugaN/9hbdaju/RL7Si7eG6xBSWO2PNwR9+
mvfNixpvL6OHYnM4LS1Xc+kOQkQsqBROF/fWbJye/A2UnIKfS5oBJJfML8yw+F0YGOuzV9MU0KnY
/CVn3cKRNDEa1eoMNNbIgT96jo47yLa2luedDernwFSV+o5Izn3N52aKOB87A+/dqNc4bEZyyYQ/
fjdNz7tGPro9SWJw9kBWzGQcnv7aKB3BbF3OOcVbUSuJ7ivuZz1dUqFjEuLTQgTvGxW0PCFJ9Uu5
N21exF2YbZ59rEh4r13Uq2ve2ugIAJ67RkRF9eLfoyo3QNY6PfZtTuE3GvMQpG6nfapR3Wvia8j4
Nz0yzLQh5ljK22MQtR2cK+DVrLgW8AE8F0ZEcwZGkVk4tr3CQS8SnS17kSdJGwcPwwc3rOI5o5mA
3LC4ZdfedJ7hjfJS4nKg/AMuAYUz7HRWrkpBy15XaXjvoeMRRWwcQ09psF/fEFuwnqT5K4JGgt+f
6nxoaJ1RSIuLlqv+98hrwXcHU1OezWRT0XhEogJvycirMgtczdESZxln2NCSzg27hulVJoli6YyB
ZsbW+fYvaL+ouqkprITTwIQN5UmkjyOAG8FyDy5TvqJw3WctqBRblbHdq+lScfpJXwmUzqUau7/q
C5QL+z6xWSWrIz/DTFpdGqibMKBYLq7XPL6eRvtIPcS4Cw9OtkVq+jTHKB+iP8BnGqRuJrR38cQk
yO4mzXH7fFC6Ns4wjhVBoLIoO3B3DB7M3ETDo0YV3g9fZXEwjnhlGxwiDyS/iMRa58z/ijk/IRCB
In/riq5cbWPi6zlD8ijIgkiDZn0pqzia0zdHz0rLWoW/PeYspKiby00tXeXb7ufSKgSrkREqd8uw
+3ssZuQ6YVghIKstXQMB4MgTtIKVlmKNbPf5IjQFbnnlCxZoE6eAdLgti6rDNcDBtU7HRe8S3hQ/
YlRjFzz14yzUBNhVQeUkzEU/0Ddko96FoRwSwkRpSlL3E/2N1oc3aPzZb9ARKWryGwanXCxCq2VJ
LAq32Cqb/seWU2cPDFOlhG4E6VV0IMht0DK5TLXVUWpOMuvj8eZ3pV6bi4r7/PpCK0EFGrD3xJC/
MFr95r2z4e4zaSAILkKY+aSKj9Gg1IDF8pGZ484RFPJFe813dBSD+NyqSdy2y9IaAeF8Dyu1mp7r
oVlGMYG6T/O7jEvach1yRBY/vhxBuhmIrjMrJ5wl4CkRcPGuj/XoC7SIvcWQ0D53Jj05pJHwuilD
TggfuSjvZepDsWdCWfLCWpB6cXhbm7+Y84yZg3wVQBKNsYs4Cm8aOFe0oU6DzKYWerYFsPwnkK8H
w+EpEFzvFLvknVrIhjBUuDt28oY1M5Ne8cD3BJRjA1hHOf1IiRGEB3ovbilqRWc3Thl54HAAfW4z
/A/Ly88eoHGodBhXB959TeBw7qhcE6gisLZoMvH4GChGa5PvAkvijDoozvS1ivL8K8v0KerhphaF
8qyIl74SvAf9rzCMPiw0nSkZvZp5i+iMokMVkgEVOada3znv0pO7kLr962lDmFa+G9ctykbYwAEb
/OdjBdabMdFuogb89PUilG/dM4eR+m4MxSkLv1lvBq04ynrvSbeCWDDsDOoD/oLFk02RHFjGkQsX
+u0bgmsLCAbDHMwcVaTJyayjoGf47qT+KGlEh/zTVcXMFimAbUs/+ANCNedSLgYlQTVqRJlUuroF
77SLBaCm68ZcYb/mpoBztrSdA/ZCfNxa/f6R/wVQKM4nXqTZbqgif2PLs1FlNMYoK3nZYZIpJlvy
OVJHHvxF9GqBC/FFCo8zqZEzrt3fFX085Ab9xoFcH1leXzfybEy/u/JY1mJYRsYHeNp2C071kfL+
ManIkQOvsQF+HdQENuPrE4o85oRb3FjdlbQHuBIDLWJ0KMJ+5tk2kfpNGRI6HIS9ZW6aD6tqDtUR
aW+fFZI1Aa0PEetG7gS3Xwqq72j1gQKxjzDNzsJ7BwpV+9M+os9JVXcYqizJ3mrJ9WU4i4l8cYIc
UlrYwJ8gIzUrgqPNVTTfn7fh7KeQaV3UFU6VP0nLD6PoPPiUAETqqTioAFtmRO+zabQt3SQeY0b+
W7SHw2aixd9q4GH9QfN8/+usLyEtawfRJwJVc/VSQp4pWglAXL4ao3V0WLhvlbGqq80ziK+2OQ28
zV3MXMpdoeOWEZUeB9lb8D0+6/Ki/1Mgl8YADHNHR5LYNjGYAMPyHxsDqkiOiKdbqrDHxGuDcGkH
7XEaAGJ0l5kdsEySm7IdN54L91eQs7in4LulmmelHMLoVeie6auDOMa81flmX7sTH6dspzeD0gsk
1FtTZXoaYBP+dCsvcdbiNsflA0gtVCCntNpT8Nq3LgS+wsG6h8eU1a9XzwNX3gK6TuPBKHtsHiG9
RZINsxS2vMiVBDeXTGNs475cFKJ2M2N3PYHHc6O2cwc2CB2oIWBFJPDtgfmkrzgGAvGE4GT4W3Rh
BDEt0Da5vnZrIg7SZPBa3p84cvLsl+DhQ1/De8hyvYoMiiHoIAA5GlyZ53H2fg/ekNpi7nIkpi5B
gAf0cV3sScIRY57nkzYXmdCH8Y78TEdTHJq2doD3xk4TBba8KUgoyyj6POtFJUBd4kq9R/CK9cuH
t6ZSjU/WZk+PSmDJO9YRYYjE5DRpyIW7fRUwKf1ud+LMgBdsfYL1UPHAY0jxQF4KGqmjKSFJLrbg
cVH+vthrXScPPqUzIyzz2oXPsLodJqzUrQ+OvXrCs8Ph/m86t2idP6Bhpzrz1aU360CavLxJdswu
OkBE2UkQjFZUo3CVBl8OODiKzZNbePMV4ejRXpK9V1RhwkZ0GQ6bq8SEWAj+lqZlol9Rv1KeIhDL
8tKWrYQXmW0s42Z6SzVnz64nFA1AFdjLNIQGbCyGr6T5hw2N0hG3YJ0mr+snAjuKYqvMj4yE03L8
BqeM93IKdJEc6whF5yAUmu44H5nSWJbWe7hoj5C9hr4NNYNZ6kDfolbxICYyFqhNJrDWqOvl0c7r
YsL52B80TbK0p3l03I/BNScNgLN1QppCubOLO+15KCp1G01ja0uxBnF7CMPmPmDTB54wjF4XKtB7
ro2S17o7Y3aYn9ot2ypexCBZ9m3PuTyu3VyCnq76wZiInU+RVFb3X8awv7Tzc28g18Z4ZD7Nc0wn
Y9NmEP2JfTVILyuonDijJhZicvo5w+wgaou4IpMJwYL5Q5zojkx22nP6zEGeSx7DLiCsAQ5J5tIv
lF50Mwor4TjOtwLIDKL29H8Cc2lLaSND7eAuxuCcUTHDtaI3tUGzc+FPoadL9b0DSwPV6xIuwzai
GvQR3JoJkCh1zeyEM78+Gq1dob839QqvGDFwdaihJN2NVOvv0rZmsL2Oy91VP4n8bgRrzf19KPzs
oninob7OTTT5BMS9q1bMecJnJuDIoycH7xUUbg4Jo4sjv4gRrsW3SRN44Lj7XH1fibPmB9YYIEmT
GoCArXTn0g8B3HwK1nSiEMSUxy7EvFxdqDT/64jSBkaa6o7OxqYUPa3LbIrQWkQN+Gcfed/RQ5NQ
VpX0LNN2JJVQzPtfE/6sSfyLKrR1hka2VRdJb7hp2rp3v724LF9rCCHKRLIdXkhXbsaLuabnOAJ4
nhSwGmxAKy1zKLmoZzAhPHS+3HYqjt7BYkidQ84XqMbBCgrremeZgc4dI1Zcr+W3IKUASXKYf1Ts
NkG4kmCJhslowJvFPeEUZG31nkcDBfg9yX6hbNrPG6x4COTbjS72dPA3UH1wDr5db8HF1D3VdZWl
bEZwPS5GC9bRg4ZJA/XrJCP9Jphbl/ieZyMKZ8+b0/4zoeN0NOt9KjLaamD4ThdukgepoLFrQiNL
b/gGb/7PYag0vvTc54zIXUVGmdrqA10RXVPcgXllvHosyrZRhTjMSNyBuWqg3xlda0SYPoven5zF
mwAG4159A4gTFNs8BAjYEe5+pKLsN9KuVRucPzIXk+6SY6pMjUCIJ2QBNzffteZjS/T7t/NlqRhb
VwBpSVdbu8bO/ScIYMtiQRvQ9MfSID9Up0uy8CTlGZ95JFEP7wWvc+N+j9Ds/7Vc3WHj+emdPImO
j2Jiq3dv84kbQ6LFk5cr5qUebY3/g4vM06K/bZvLkEZJEZV3QbSXQAmOOGDop7zqibaP3G8vASet
WyC3CG+FMDGHaP25PkM5ILq6T90RMdEgfFhrHXhI4GxRn83LjtyZU6eRDnvE0PPiKUYXAZiwwfpg
vZ+D3yWNubArOASc+7LgqFjYvUy3K6M6m9m81jG6nXaQcLGOA8y8HbqXyREJ+3ukk4mEvVeAKp69
owcc5PvnIBXjnYUcHjSFaGwcoxyaDD5asITqIasCS2zyBbllkLnQLpINf6qT4LLn+xhGbBkmhb+z
zbkZfVvsMZb2/+U5fFxc+4V1Bw5lK1U6aKw+SKpOZ3LiT3doir0YSvjYwUaSeAXMY9iLuK+AMAAx
pH2S43BJRMXdxOXc2R7aiVEPrGFJPrEbNOyvlBR4ndUtnXdz+tVO7gq3NmqSUaekcBwx2iY9dyNo
rV4uXGL49Cxx8rdAeFpHWzTf4wY4O+925ydhYJaajlojjcs7kSzoFXp13f2aPz35A5eN98Be6gWD
FOBCmzy2t///anMOLaajbt/EkK78wNnhc+gbR5Mels+c17DQElyoGfQTrY47x1Pe+kLv1zHeu93l
QaGksKZgBx3FjOmkBwWQamrBxuadbwUIRwC/8WMTtj6EjNWg3NJ3ETseQRt5RXIbi858ix+CgWbZ
o9HMw7+Qxl6rxZAhzRLq+ah1Xwve7dkQG2opH++Xh1rxPRznJBhoqr49MxcEGTvwJnYab89iDk7O
+TlSGfbkw9UeZk0IJUUQtqd+5E06+la7ka6X+pktMbjt2g2sQhJ9TMk49Rp5TewVCF6Zqhqmm6Lc
WP6HFGwdpPei/1uwYLTeeibYbHaijmXZY8Y8pVs8xHCqXnU1ZsYBpYDBfn0eV9O0KWaaTFKVPRMp
Z0MgvaOdeYiGVpeFr+0qCJ5aZiUUxaWPkaqm/g3w5/qxR9/KFjkh4nmCtWRr7f1WBMMac3qnjFpV
yZpwUvbxmMrL9A4z1yA2stIT7Kw1tMRo2Lo9dhrx3EyydDsIGv7Qh35y5lSrIltphVWxU9+hvPbc
uQ7ZMav9OmftqxjO7Ddp0ngRR2Nqlp7VRl9ogszym7vouymqlHHc4Do+2WiJA2o4+pq43RqtRK7+
Q4NPeU7ajoaTCLGdk435i99B5wCWrTiJM3QWDhRLHzf3jhEwb7amc+JDPos9EFOG+HfrXfXJHORq
9Gr0qUWUqzCro1Wy9L3pugMLFnOn+yYgjdL0kJ2eszn5kWPpwk0BjXgQzd9sCtufMkrL5cpUWye0
pFlzZ8bdZM51/xpF6DMOACj0Q5fnNmqAP/ZIaTJTHeJzpdU/Fx6IKrFWVxiqFl4ArhcVMeZEyOO+
SpSmAC5BCx6/lmp38u8riQCG3zgsd4pNJq6sYVyAZw6A3AjCT79zsHW084MA7Z83ML0y82PpR5Py
Kt9LcY+XbHMRFD31/GIRgcwUSxhNI6JZfWt5wCHwhPYxsK+Hb8KgiYSIerdj/7+a0Zo/qNT2FYOB
VCDNhxFRSpcSmROhSszYDuA0GLu85lkLj62iOXOheJg0upRQ0O3K6WeYRipo2cpY7Qm+aG0m2CDH
/k52nBDSV75bISEwsdFK/P+LfrYSXgVeyjrqT/zlt7ceUS9+Cm8k87ZGdx1DoE4tRTG7OyuUQTzm
kxhdbv35Kuvr4eezIavrUNZoH3ELWNSwrWYxbX8EBH2ou40ppIjGSEs6BHJP4IlFCVQbQyAMo2nn
kWKkRdLfC6lkBLvEqFNOGDsMV/uLNBFABrBDcz12G6UDkCGZ0Ew5kXFkPRbqRG4h9+uRQSz5tW7e
NKElOGwLsxoxI+G7obgUgx7STAhHdhUwZgV07n/XyIhTuCn2QDiuCORf3Cdcr/KyKLtAFtVJhtn6
zI7IWVhWMqBDEcKJNULIf9BWMA/O6xiy8fg4JRzSxKNtt9s0wyn9anvuqxyofcVWKqwUsu8wr+8Y
Gac7wapytihzhDZ7Ug5kkOdCxaYSMrlKS02XIMieDMqjJEjTrLbqElItJgjBS9uafzHRG7YvWXdS
nG0zgHUds+9l06RH5yIrvrz4VIFovh7S74Zm8wydZUYRYiihIlCMR2yXE/C2tXBDGx/i1Y6/eY1z
81V0PZOd0WCt652g0I8QktC0c9DxBuzgH6YnQbHwzpgDo3btYtaBopw2sZln6icNojjY6lcfkmBB
uF8xS7bxriBHGYQpnqmkOAit6nzWFX4oIvKUYVBgyXJSMLrP2E/Mm9VA2Vg+pTgDrUV7qp/PgVOF
KX8pUaclvJBpdOcAEGnQEBFAsjaD1kYBTHdQvXBYbPXOw8O0AoqElxxNr0lNNdvb5iYHCW9V41Kf
sQrIGmb3/T0l26CmaeciS2qHvvBz0nK8qzmHzqiI5nhPwxa8zM7vMvgSqZ68yIJH23LF5Kc2Pp5s
aGUCm+LC4w/fW3098yi9HPCsN22GhX33hBeTJ8EXKmiALbLRTdvMTEDMsE1z/Y5i9bzs3xp6cbm5
Q8j/ORwoUqJaOu4tBOa/+2kp3FH7Jp3Ho4HTzqqveKAm+jCje0q+b1h6L4SYyj3teIk7mumMuwNr
7FI7WveGY6UdcNmKdxDsZHtXYQ03sChdD283rVrBCLkjlSwqfJpDC0I/Tj+TQgFAYq6cAW8zCeOt
e9sa+bn9+YSa4INYhKAI785hFkyQcRy6L+3hBr26P24aT7iZCkDYMG5XSKep8zlXPTUshSSL77OU
bIzHOou8hsHoAtY7oUFebNoog8gY6oL99IoGeabFO4rKjcQ/kvpkmf3BZW8WhvsFiolDHLDAkeha
WlPXSaJXCLAp28Ed5T3KRnXlgeGKGlwbxWx1hKzPrUlmRwxham2/geOCgrosWWX+boNTNB3JRGmx
Yhzzty6qoJEuiF7mh/sNDgGsKkfbcIQFpJ1NbFjc7SBvE106IQA+ZQhQ/Xbh8zf4VR8KeQXR5vvc
T4IUn5VBQB9IZ8/5nLQMe9fWVKypRKCr3HM3AWEgRx67RGJeyUkBBl3k7vN1t0+CYv23j46cz4Dz
oaM/zMfsRNTNc7fQfQeRpCmu/+u/yMRhsOveIJpXDQkWcm/0LvVpkCz/pLNfVMSmQXxepGTqDA/O
e4DYJ5q4EBe6Om/aq3jHWoUVyQr1oG6/EsnvBDF0PKKbGaTpBLP9FifdhQw2OnhMJDFqgBIdAXQJ
6Z78WAjCqLhws4x+qR11gPmFRdKqZ5FhlZnZwMnxwEgDfMKGFH4MgP+YioulMGJM2DNpkjDcRKWV
hssu1jYkiDqAMtI8+pPDEnXubwpw/xq1xLdDO9kNEr4Qc3IAp1R2ZZTFiTstgDaTj6+eu8UTRgfs
CCRZ5XhlSWn+9vygXGE1RCHsmzUUnHP033auiq8WhMr10NFJZAENYnyiplGmG3bJ2GSc9V2Ehrs0
hvw7HaSa9kj2hziFBzvU9XfvwksJM4TsWy6DrcLTwzxB4i0HPwhztJcGdJbkY2DZjYZf41FPrASA
DSXsFzSDO6hDqUx29TRx3LHRf22iaiG1EVJbxGMoVKhlC6O2xiMZBjp9OddHedo4pBAi2+4HcJf3
OyjYbwnL/7V1jEWMxNsoTf0gCluBcc+GARsi1f2x0AYNwlQKFyHClxzK4pqD4LzFQAXuEgyKuda5
/2jfgcvQ1C9algNRwz/a05EJNmWoiP6/FKmuxKOmM6WxArmWSH+9PIks0aerXf09ysdxe/K7soDH
gQ1y15ddpIYpHTlEjc39gSxFp+zeSdUxnKO0qxnriNsf/fwwcXiEXnjIH9R/OU2FxGqZBe1zWAnA
XrudMKsneb/huDh9QK/0YqApBns5KxPTvA/chutOsMZZm8cbJAJdMqvAO0vuZ703J6n6UgGcdGNE
b53N8ySoN3WPAVpZZsD1haSLoNf+2WlOlvIecwbKtxWucpVZjv42jAcDviKbr0hpoE8WK2B7mmNg
vitfpaAGB/vQYlVkQinVm82UbtpR8LUMEk5dF63bpmCyD2Hm2+9RTPINcLYbN+gQH0WYtogEEa33
lRf2J1ZxRv7pYq4+wyLapV7nV4doaMHHw2BjakhkQGTvrg5rFKQ+atWP9ntIr0rV8TK35ScTuDFl
JCCKf+ky8pyr/d48hDELQPvhnRekjykd1BEmpGNu85m0skXSXmjHsQnlivmhqf/VuDilE4DcZDzx
P82sRruph0BCYsIBydRpURgCILs2xb54h3ojkB7PMgdkaob00C6d2LsY/SmsXlGmWOh5EWepFPds
JkZq4ka/VA1vCPKVyI4uBMGDhsSSd9wEsAyTxdWIftSRLn10ME1xPkyQi/UH3ZVDhK1VdiSDPRhs
2I9X1MX0IxrYCyqE4Lyzme5dRgpUH1AnMZuRLveI2Ex9RtUcILpYDbY/O7mqOTlsYtCZBE/HSsL5
1SJnSIrb7wn3pB3ioegBOeVr2zxCW2ENLiotLPzzovQ/l9SR6wbQrHSkSUh2NaKM7iRrTAbysTCm
hIfsPFl92x3r0bIzxhcKzsCE/wCuEaXAYKMbavnVF9sXugu2nFAwi4/7nRwtApsJS61dlBsRilYK
WM6YaaH7GJtLP0M149r3+AhhW9TOlzsLnz0b8ljwBJr9ZIU6/xwajJsvjAy5wydXVrfeI5PfEsY2
Lg/Z1/1qrGXM8eMLGwi1IclfP075JTpEPInRfHL/veACN2UEQMpYNjpiTNC+iLMM4bx62hh9pzSL
gFYmDbeGwZZoxR9rRZSgFHGTOcNTbsT/+tSRZ//LnObyR9TjLoV2N5e7H4GdeN/p106CbtsqFb5b
pA5JGZpAWtHrRsQVAIFrwxRfEeom22HPkDORuIIJs/T9ynfZLAqdQdqJSpg51hooam6VFI3aYMHM
34hqwaOd94Qa3vVcxYZGIcKvoLL9RUkcfxIgrRNNtkuCGXIhHXa7mHazP7SIqXM7jBgKHmaexStN
oMS+OMfn0aLgCpiPDAWWD+yXfqEMJKsQj7Vz472pGwPV47qbk1aeIEo4j9PX2q4WE6bbvvPYUEJI
r1jwvB2ZhFWWVN+HhtsyhGvuPO6mOyyGAkcp2fYVKM683Gng+CNTaxByrrW7bgEelZ8KfOlQY75U
+yJnRTQCKfqloDo0mOKsjM0p51N71RpQpOQmWfgWu8QLCle2WrCjOr9lBo1oz0t1YOK1YN88XzKY
IpZhn/RnYOXVT9qoe97HK6Z2JVeg2G4W8lefCawzO2w6ZTzue6YsjnPxByqIRiyfA/87bbYN/saA
3jpXkMiSMIh1Stavxcfpf0SM7qh8Kdme94+ChqMtk7PtKur2FIIHynfTZTWZt3u7p4iX8lOk9BDw
ol1qcW2OP6hgulKOo/nrivx+dW3r9WWpaMgcJft/J56PvJhunTWtHv2Kg0QtmvJ9UJ3xtSG6e4v+
oPwQ5iaCqSVlD+IZffNjNuVMkKF0ayHr8cv1uFrMN8NKuQB6mGxd7QqulRc6S0dYLZqLHtfFqMmH
Blkgaes+mC22m0J9KIlqE2Q7kW9KpwE81ncuyrpP2Z8yk/cMI5EiLZ+FuyLcKc/4qJew7HYbycDx
t5vDgKu1CbJtp3QR6upzUe3yi4PqevHhCHN+OgKhBkmQnamYH3vb6+XBhYYtNzLWilhEGmUoxFBS
ltNZ6/CBKsm0jEK5mhwqoUBrRglsUayx38tJD6/X29egB+gz2BSBe8vuv7NDhgxA4mD2wTRrpkuL
GA4tFN3t5jaWB5B/Tq+kYVzpSjZIYb0J7q5zZlr06Rrv6qdnKG5tZ9SwFqrQGYNHf2kh2dkBd/7F
P/P+P+at1WJo5B1c0G2yO8rsUoamoWjbF49OG+Lku+He5BqUsia7khN3H9SPxeRad/uB3a6Ysc7N
pq/QCKsVTjBBLpcSTXzyosg609si0ZrtFrcRgU+dXuUdzj7Pc+CWWbItt81ghgnxT4xmlCtBbzSL
xbaJslwuVDtj8u6iS7QTt9EGtJUhN4qch3gXeYW/6AWGqea5kALzBPobIcvUVdYVMHeJ7yc+xhha
jnTkiv/Uv6FR1IY5T2lXNm3L+n6iqHGYGvaW6KH8VVL/2fIkI9Ot5y7EGY6BTdt6wDGQa/46seTp
MMQE/Fs8Dw9pVnB7mfak1dY1ZHqdN0XXonpt95txUTwuP9HY3/vnBHewZPckoc67kCfWndEmol5m
7y4xVtW1Kdx5tVnzzl6OuQrb+oBEkTYMyKHwAotw0Vt/gWVITQzSlsNbSWTcpGzRxmhdguqWeHWh
+4LKYEwZvrq3JcCnj0uXNd7huLak0poiYrpnXGW31l3djm3juSLPe8t0bya9MgHoFPHDLaiDyzEi
Ewy1KQsizOdVkB2uHh7fr5r0qLysaiPucezDK6P7dNT0QdDA/WD8TchpwtL6VnL/7OAvZXBoIFRL
Ma0+0/k3mj3/x/3Kg4nyvQjw9XCiYI+LHEl+dyXliJj/xx2XS5Gxpen7MihmArMeF2KI8stKWRHA
gPTGLaWVZzGXV94pY+habAL/7VOu20Wv/mGv+YHUtpmKnpgilCWEFcQBtk4JSA845rpq+M0CQW/J
3XLrlCGRqyw/rUESJAIkOaO/245bnN8qs8hTn13pZDXadBxrUYyX3zhRGinScsgbUmqz+e9ClvUd
x0oHZ+WInusoLwN678Brjc11dEIXo2CSy6tGmQp2h0P61VfB5qlz1s3eRjb/qbIJCoPZKVbF8jrp
QP279R232iEGQ1E6FMYW595yKdsOKADTdywa3u2wQ6eZ+EGnBF6lC98U+fny00bWnLPYMMA1OQpd
s8xUuV3OduaYaLZYsFckqCar0X6j1CDousgEL3nqWYbx1PsFe8CesTckX/+6BfyxY2KGoyhO/chi
D4bq7KPOGCsu5Ds/+fan2FaU3Ivrq4W/TYSHHRmMAtCnrBLX2K5NHqd3eAlyLpUbeTwrWNsLGmG7
czKtztmT1Qc1cMJrflUgsFJfnGuUPmvCqJonnnJr6yx/Eg3anaFrytkvAVOEEIXkjFftj+ZaXMpx
KsGiVBea61w325+p6EpYf/69GJy6BpZboAr64lHpgG5A141GrJVlTd3Dx7F9of8XXvkEJ68mOah1
hhD4wuQRnOBAoJG8vvEAJUJNV5IkXHHNg5BiwEMsvRPeY/P1WPDc+7pJxgRsICr7ucBMYu7JfnEF
Td8eIIDWI6ng6H/OjQJTo/RNIrQcVHn2XLbHsq0aU6eUiYwT4sw4fL15LTsTo+VJmJ3C8/CH4S6s
p973Ykuhe8KqaKBkWhtXMdhPxTS0o7llDYjNt626xy4LfjixU2fJGD5YazsO7IRiNWRKGnzDM/HR
o5OyirO0UxT/njHLkBqASRUfPjmZ8wY8MeNGbrObA27QcFAmYpsQcZjF2HXWnmCmStXlrLG3yIKi
ctvXjP2WJlo/jjwjnsiHEHXJuBfUUZyeJRt4hNEP4xNBPZPviP0UmCQwdxjSF2pd+GVSUYpXhWOB
S9kGj+j87c8Vshx0I/7p6NEE5MEWgKBJOa/fH6bzPn2rOFf+Sw32UC078xuczuP2xfF9BhAqTQl7
ERK1Q8Eslox4EqMknCRkE+xvIctWDMY7O/rR+3eyLW0yB6nMpY12//hYdkfUKgdg4ngLFxMBJ7ix
3yRcEoykAot2s9UHipTITpN4kG18EKMGiJoMnSsQr6mKx+qAsLqtfOsh+G8ggCnX1bOCZo4Vsxn5
F0+XgQoR+iAG4O5vQrPJ6TZJ14vQOKty2ehWwXLfLTrs+Da2vwx2bKp0CtVJ/rvIBNUTPU1imeNa
LnJH00tjijxOAShNPBDGD1fv/9p5jpjHU+lf2ZLkMQxHtekRCj7KNWHnHRW6PMc/zUvVg44Biuaj
cAbmuo1ETe9EfuoaJFzc7m7khzLgDeZE/0B19006+lr3+8h9/gc3abfTshaUAos3+40gUR4EGiNc
csb8ZOPo0fmZdz53mbwQ6fnhNuim+KQ+YWR22sGkvuQr6aeZubL8FlpOMYlANIz191HOtNhoNERz
YDWTVuYPvGGCBrLnkWbN+zvOtxuiKxAtsO0S/Xv3utJ3ZHEOw74KP9MsqggBAjP9HGhcBbFUY+fj
22CsFS2xP1ftzSad6rAr0OL1wCi73JLKgmi5S77FPVuSx9Ti4E3gCdbLCye/xCXCKPK6LExIopI0
fweDOSZJp0GXla0e2YcDZaVj2donGErc8DkxR4nstWkJggEiF1/bKuRIy9scF/Sv3kLDVw8G2R7j
UVc4O3zKYIBsWtLxzDWuKo94gqa6XJNYiLhNQYJCG+8CttF86rZ+YFvd1j1+kxnlKKdn6B9UxtSs
YTwDT0Aea1/CHCdolQ6nogYFV38Vs5Zwmt8xI5DGI9yoclyt7lypY/JSSaFhmQxNPZcZzKKMbyXI
oS9awogvnq6gkxGlSjdYmbvm+E3ssEk2WkBDEpC80ErDGOjWeeuvSkplruVUXPBqLUOrOzmHlEJX
b1j1PWBLcsLtLe1yco28SrwgShLx0DkI53lwWskF93vyrPPj2TedZEo9uFKH7BaORkjZnFR/fwJL
5uH+SW3nGT7TaCNvF/PT+cCUEc22X4UZcSpFgVY6JFPpl/agTAjvWFFVGU37uLQG1wIpYy0e6wko
ti9ptfy3kilzQSGsHA7L7bCrw5LNUZrqnKPn9AQSmu/i3n32UHWKW5R8PAStvA5tYoL0g/wO80K8
68yVePJf85kANVDELZx7SPAtpwCRixhBLsg0m9ei+YTHrNBi+VywKRdd0UC3dmdqEC94eNDygUU/
/an9ToVlIK6OjaYij9DrY6LNQJ0xWQ3A7llnwaf/bsgJGElZ9h8NUqlI8OZzwm2/D58njS6XA6+b
HA0wU4PX8asiQUizd3eGFv8ZcOzomlG8CHmczZvy/Mvep/9eFjOaXNnsbXx1YeZ+lpQxcnAjjqJ6
1OJ5CKrnZ6437toNAQs94tO1DdBqHHSL2gV5H32fJT4s88/F7CzU35ZM+I7JPbjvEho89otCq7hc
PRc38k2fWuUFW+aa38JQeK02hnjv2BYNfPkYFKctiPp/BBWdAH2p54wjsBnZ/YUUNdV+1i5iw1vn
uqvtG64olQ69nAUCDjKRLH2CMKReWteNVKSCdOTBqd9suSypeGb28DBz1DBKB9wy/SXE/SPCSoca
D6w+MB7Sa8lrJzLmRdxqvnnyTwzlD0gxqLM2PtNbyFwELeXq0v1HBz0jYp9VpHsx3+kT/yE+VzWR
VnRCc6F/cHq7ZunX9S/unbT36q1PTik1w1rjNN6ifP4x0P3CgE4t/aPYzyyWmnzJlnXutkTaaLRW
hYKE3XLFASZ1oedbzSirE2+wmd6WM6WMtiDBkaBXZd8kvXhnTdm4nQulpT9HZBy+X90NmfbAIkDo
CzJN0KsTqGB6RRAomcnPwyIxv8/SJPUYHszo/BKMe0G7WsPSj2bfO+qeroFmQgTqIMUEZQO5jZYu
/REEqkh8IVLDvQ4BLBYiIGZEOoSnAel6KWAAlEqvZkJo0jIR2PfMUz1O2/NeG3L4yjs0BBcWvSDq
AHJQoC1xNyFQ4qYkSCL2E9f6Xa5QxVDZ4Bc7PnN5d1zb1LAszLh1XtyqLu72ZDvOHFSrJgaPGb8n
P6tVidcaumalqJvg3UiZ0O1tqDIFE1IvgDfe8nHv1NAnou8ONzuBBEBWwp8iyJh8RHlytQiU0gfg
oPKg0bULXrjFCih9UTLyyDtk2UhGzNbdhUzp2KaYNYa0hFdgdeBfrRsRX/ZsabkBW+h9WNN2n+D0
otgAWgmOMjrZaYtK1mUroDS57z/+IIFR6m2gududfH2lc6YM307Boq16SBneS9xckyTNNdjntevl
UB9iu5mEVrtRHsb7ZSJa7vbK+n/99MkodeLYIwd78nbe1d1Btk5ppx/e2cA583deT7E+rBbS+P8M
sFqIZ6hiqC19RpFIpsl/Kv0sqn6aODg3F0UKuukBJEGIql6AsY4U/Q/IzS3iGQDJjDBIlWFQQsPH
qm1uGEUKR3UssUvuMq1GXj2c5StaBwlK7Hflk0dTZIEshXoEY4lqYNPHEQXj/bX6sNjHwrB8n26c
ErubF4AeMpfTha1VYGrQmlvom4/6Jna4iqupLgOOMMHGq/Qv6GxrZ7QU+QDsk5sPVB3OO/G7l0kJ
/MNhYletnlJAIh2vRUcOyCeFpa+DaCHY79chY7YVGQmyv1nTFXoem8lFe8Rk3fn4yHfdPrHWIgAi
l8CoN3BrJ2OaLi9nfC8WTw/fmnqVmPnLgV1cFiKFxwR4ZarjDEOqPyF5h9jzEzB0eK+wJf5ADgqz
stkdxK7jgwalUPuv+XHHxzR2/Em5Ih4nyN65T1fy2fPYe6XYBW4s9G+VJ4CHx+2gcdzzDu6eF+f0
VvP4dw+f1+M9Vbz7TFRFSyp0fnlSXBn7vPIhogvmHGwqaTN5nm4s8BkWO+y4PDZDEHQwuH+/wwv5
w4WPQGFfp7rU/JI1cvULOODRP0JxKoG2NLjGlMF7DfNKZenYzsN1M96PyQ4zSOgk6usUBC9fqmzV
/bCTTQ4BqGP01yLJi9e3BK6PSfwQN3joHngXgOgfTKjebAyOyDBUmiWawH0bFSV183v1MeVYEVdz
7linBbzZq1QiWgUSU8dYYVMOsPTtDfsgxSFFh+eBW3JPDAbjr1VAuxkqS6bNM0TNhxNDPA3E3IMR
OfVxlZBO/BLaE2xECwLWh/HWZGzUo0Xczx19OsAdsA8IKyiqTjt5ekLru+UQOdlkK3RhknQCdt/c
wddlHyv0WhMdNMgWiKZBumFAn5VZNVKPmzf6bU/2OSZITZdYFZi8IrJ3R8EC49mX46RkE6A1Cf0x
5aQ3qNH3freVyGNslcdI5Pp7o8CdP+tSLpflH9o8pA4iOtO6ZFc7/OtNLSwLQ7AHfDzc+QQBdaEL
36P4bnrbPWEZmFmU1jBOBs8fIlt0tehzdCMDNnKiKKz7vTh/U2vU97Ym4bWEpNL+RxTn11MUS9U6
R0TOFhT8HuAp2ZlF831Vv4c8mvMfltYmIoFV9mCN94LQY9h3iwMroJHhB8eB0AITno3i7Phk1NQu
sJFb0Q5grAa+rc/bXNd4DhGb1VTvSGpA3OLx6gBnGegP5AL9XvGup6XGrgbyvfQ+LNqpkryOzmNw
83uvasAoeHIDoKv7mad3Zco9k0SxgxGqj7Gn/HKwyufNb7UaPq7KVmU+853GRWM9/qOE9J4/EMkh
hDzODrYjvLspJJMamUCwJvQ1+9NUG6eNCysHsyzLtH+vYhNQg+AtvdD+dDLNnjJxTdUeebPLYlII
nYkyFmcbqOUZMBDM7oAEGk4yfEeplYfuwPvzfxCO+soMib85lqFB3kGyUj4VC7awKvFo+2UyJP42
rB9c3EH1+6ueP9RgcMq0kZHHy+zQMxxZfwGvvmBwSoQtoJnfPI3Wtr2DN6EG+/XEUzp0T434FgAM
ZvP9BinioGmZCGoSaJ+ZGoxsI93+UCyaxPW9AoOOHKKJ+LO/9LzRW2U9ddQLvoto/9JCreUgGbGD
/9Dxk37ecblEg/DEFdns02YnuH3kzVAnN+KDCxVz2tg92nZNP4YrsECjpOC9ckoh9lqQQcWZpUbr
Dt+z3KbFNEXeoBB5kZxcFbb1i7PGL0Zo+oiYKarwzzcggUvZM8zZUWCtDXBx94yQbTQVnXSV9iY/
JSXobH4zOlSPu5RtOHIWutEnaVD0fObGlPLaXGS+GSAfPv2xnBmx0Jq0rin9QHiiy25M6XVd34sG
m4WdgRhS679kEOGy7noKBNDLge81TJsK5k3f89BMuvfpkvPEvCEVtgf8GcZU0p0QSrx6qnF9S5j4
K64tkgd8ICax9Cun5jy3fzbv2T1XXpeu7T3ZPW9d+fbwmsL281vbPpSYJauiTpnJqKwBdvLIzUmD
n90ILmart+/FSEoEbzsDX0mkQQc6CwlRNgST0+90hZPUWfAeyRpDbHB1C2PETwzeolHb+5oBlo6o
s4+pisbxdZdVXpktA0+fc1dA5pZBmv+x4ja25iqxDchb/hMunIc0VbzfhgAhb7eISIiPcIRB61EJ
NkXQZ1lN7NyhRrca7BXWAA6KZRAfpqIodEqIkVZEM+DGyX9eqNOYCGwFvYd/EYSpJ63J/MQ7HOUw
1DCqXDCtKRxuBYOIoNxU6SgT8SUslF4DZKTYFovtbn+QgjwRc+vHE5IAjUu1JMct5dOHYlgTfZzk
Z+UNvS61NV5TxIPYptdaABt5M+teP+INvu/OmMDweo0r3Na8ZZw6iRj0Yfv5L93nHVuNIZ9uBJkH
EqK230UBhpjTC/c/uL8+/KmQPOdJqEcgW1K/UIsB/eCbzp8Msw8c8qaGJhzfnkaCZapNuss/IkBa
zc7cSnJPW7a+zapGuvRXCTPI59OPmprYRA1H1NZsKi0kRb5sdwwhZuqBQX31N/CrGWxg42OAeKOM
EpFjVMwlZjw/7QN44caWgOefmJjmY8zotYUFI/p/sGqa7QZLVA54BaTfZjaP1SRSQ+pF1UJNqxkY
IbHgEQrUwN5lLKNjEziD283R4nV44EDux530F0eyjp9LBksTCmSmDpaY3S69kagNtaAhFV1fl9+P
V2kPq3AqOCZSy3fM9rJSer8gDZg7so4PfJGckus/vJ00skO+/WxJ73MRSrBSRWBUslhPZvR3VL5M
SI7YRyDMWkde2oNx0c2STAjWTsYamx5BkgNroHpvModga3JFrkCKC708A403zdCn5tTUXnbzOGvV
Jruf2NZW0+6YfPpAlLoXIwFjPryXuP0w+cC4QN2Tt39AV1GYOSMuamv6/xVf375LR12VmJ8W/o3J
EYPBvI6ortUJ+4vjffrMFqNsVo54nDl4nVTFAuKwtJ9dFTnGZ7ErN4KVSdoufhBWZKr827lf9qxr
m8Q21U5sKbdcKHumGrBU8Xr3CjGSW6Y+PehA77LYKbj9Sll7gzQOJe86FcIU3TXmuix1l2v1Zhib
t/+XjYHIEMif6E0kGRkd0jf+ks7eTIBvmYSpmFrPUH+gaOwqviagfOxMdPQJ+vv4FHh/Osls2JFu
p/zad/AXnqh9DUJEL0mat6btIXD5VkvbVq3tmj9lLtu8CI9ZnFsbuUjPnU+93azY4CstmsF1jRtC
qZ4600773YGEliqL+S+mGYiq6pm4dr/IHBMcn7MPiRqNDk2GM6Sk79nZXOQnFY2G6FlSliBbxqQf
S3/Q1B3Ih/RPQZckAYG6lRZHaFXTTaRpegWGUl671ovSii58AkvrgogNtkWZLKVg3/4ndO6xx+ZN
SS+9mVbN6ta1TGDJnhYd9nsz/v0XaxGkfUkYRKiwIUzXaaKAw5QPz9IBCfVMsZ3sEVWDj/NDcE7v
aDZbSEg8SHYkE4ntb5C4tMEtaD0Au7nsDtOm/Jo1Gjac6ntVgj8xS7Izb9Hgu4a+NbWRZnJxklVK
d2Mf1Hpm5mlIBVzV+LaP9HNkMACXhUllaBRbqk1tlP7p54eGO35vE+Qt4KWpLU56o4LPECgsNgId
/7SgVNpl265v1DURl3CDrxzb/nDQj2QbUQ57uUOZXABnMUShNdf5PjgWuT11mzxRiTxGRmfUN4IX
BTelsaHedsKEoTh8GQOOe+aTUyhIRJ3JSUW3HHMvIyCeppIVZSXEXxhrso+EzsRSXMTj5XdMqrhH
M4+UA2Zhn+mAYt6WYB6HGfo3SrDHm2L3K3RHJboeotfGu16mTmF+Eb3DOuKhzxDFSlk5Zpnsy0S0
iCzlZEBTAyXYE/pOa+OlagFmoWDAODISMvoaZEy7IyYq/wqX1nSUH0GWDwRHqP7CxN2MPgBOtO/B
gnZrN/bVm3cgd5vUCemrV12Lg3e3mQcGX8sZCiw0dsfZrRSPu+y0wAp37NjcLaM7QBq/MRCrhT4T
Hy8h+c7wc7u6PztYT+Rs9QDc/F+FQlV3IqphARMVjsQEL3Ln0yohitkhRalGHFcS66WRdaRPWMKr
gkiM7AyLizVCYpncVPODgjGkWxCtKqzgyrTo/QbJbrsA/OkT72Cla0O+j9fAal4hasfCzlWvuS8j
WgTFCpcWZnsa4jReDL178yWd+Dc7fT6PdQKX1JSfCsCPPHTL+vzvhhQCE7Uypvaf0P0aBfIxiKKK
SQqOCjbbO09BzLzqQNSebaCmGv6rPusArANBbRWliO4uDeesiP6huEpfbeqr7zTnOtpWdw7NQOan
de/0KZwTx0MXDzWb+VxssJ6btHGpDHzsbmjLEB+ST48sBwfzkDIIxRB5pb5TIuNKK/Ffmip97Whv
Gl9i9k2n30gez9BBpB/KcLXgv0z8ut0CxiW1pytnLCzvUdd8CGPbGAZuFtTbL+MzKoMqHC/i0DOk
UpI8CADwfcD7KUs2GimdmOR4/iHPyFrIvIyMVqjaCiflmR7G7uvCHp3hAuk/FxNjFdRnBdc+XSF2
Lob1+w7TlhFMxKIsMA3Zyc8IFNXod2Cn3eryaKkeHcXwhWb1eeDiTx7Xy1CuxFWSs3WaXz4nQlbj
U+yyACJrkEGupdGUitRD9+nAEoI5SOCtytrY0QOKKQy62p/xgVfnAY0VsMlf5S8Q+QpjWr5afwyP
dYrkbvo4xC0ccTVn0xCmahA5T9XI8RT5sSKrYu2iIR1qyQ9xWyWv3Ydb3Jm2UOXc8eZa5B0aCrc6
ePg9a7w59lI4Rr48oxu4Hdte2eU1FVpTGgv9C1OO080lKpkpCWdzLaWmKntkpbaCvJIi8RvrtilT
YEK/QoDfnGONv577PlayUZ1FLzeHHITHZ7Xl7nEFqNa5BEy5lRWbdBJOJRf6OmmXzwgZc5cAERHc
7QzrsE3aa0iv9Z/qD/uaXPWGWp0JSsLS7r5V/uIbOr8R9YHyd+CFDW/aGcHtTc924xcsWP/T5hBs
amu0OdF/iEgbju8PFhfbwOwa7HdfBqy/mQmQYm8YZWk/X3+wnbzeX4M5zh10wJTeBezN+WGJiDj9
Mv8rM+j6CeP67vjPf0Xo8JHRFcwjakl/Jrd4SuYq9J3mB2XPl8M9MyyHXWO++6pepV2Xs9oLsRol
1qrY4WLZbkVJDs59IESr/32qkp3c7KlgnD4qyyVlA+uKNQsElKAOwP6MWLqBCwVuyNjhFHd7jdeL
zOMKdMkyQGEbU+1cd2snqGVGflSqcwbxq04k9zYSIxdaTUeSIe6G6jxOt4l4cQvSXVORshVltGkd
qV3YUEC7TqQa15DVxY5hbGYMgL4snviHQdfsQ5T1xGaEgJxd6Bc2CV+t3k4GbENs+DxFo8NUV0ot
voOgj/ndEO5DOctEQMdAagU3Wva/Z3Hq7+/O7GAhI4b7lqkJb5ygKqcHffiRF1izGA/yTZqyr7pU
SWCBbpR1ZsQOl53UEjcwdjm4exvZbjyCjTZMcE2+MH05C8Rv1jmacD1Lq/55TiKLenqffmansT8A
v9PI8BYICgR5PGqRbJkaB+TcK8FS1GdEvGzNwGVbJIdlB+Qz5oW5dPO2MOMl2olvpDA3NOt/DZ1o
G5YX/zxFlpZqXjQ9SRHvYCQDD3+0dEyAy4BBUf66QsRY0O4iGfIEbzFiZVdGhnRlJzJA1NGW8FLa
Je4uI1wFgbdN0dzdhbit6feLe7FSlXR6t7UP7B08kAbo9+qpI8/ANx0hnLWNs1K8M8D3trSysVW5
6S0mo8Ijl2j+ezPV/84fLMqVDkihEtZJLCKxotWDzNldgGc6XvLj1INUlehUWoKXtDOOZFBaQ4mP
CsX+q5nCygl5T6geeWqm6gLn7mrIefTpgkd5YMw8BSiNYjg44Q3MpbsSJaotBmvUgRLnBY0amt3T
YhZH1v4Bg3jrmml9hrZuCtQ7P4oQx/rcN87h/iL0JnwsWzdNJTbgfsy3gKdHDg9qvSH+P7cxpVCT
AAgb4KhewORU08Btbhh6SKNa42hKuzBWyIbKMqreJDHvbrQnM9keDMu85AA+nAUwPHsPkAU/4m4+
rRuwUkBMeBuDiJccrIospmyP1/3ZrNUk8U2rtxNRYp6F28sRXieLTLvnL/kNcny4EK4pE3ITE01p
EVn1bUQWh8NrPBSYR0C1Cm9m8FMxbMNYZH6PToVFUeSsjHl0SRckt8TGnUbUdXc+GoIs/kzd6liL
VTc00Z+ORVfezyVWq0oXI6H4R5j9HowkuzMfI5P3SVZBrESC4RmHOLh32SgDE2rY06/45tza5H4K
guQhnnofwwAdN4P/baHRAeJGAOJaa+J5BJDazo7+CNqddJqesz+FK0ofT+GUXqV7PSpasB/rncfu
8ku1Hcq9PAyTWtKSF2GndYoxFNBxJES7Tmk4csvpKtvn+QFxksqUmP99b5AXgCznwrHi7Jfixgyg
mNB7jI9ETiKgS94kIx2fdor9Qr//6cBvzrCgLt1dGPBG3AIbcj14ku8J6mxZog5ClVNBLo1OdcLT
Ps1QFK59gOjJOaqsJYV8zEk83xU9sPa7VhMYXg0E6wcd8rUzhdMV5E6x9lkhj6xcYJZ3Y5zBSNQX
WZkJ7JtSfW+C9r1GqvniuCgoiGeiHwCE+FMy/B1+/wG6MeeET8e8HczlPyUU/39VLiyk5Gdv2VDP
s/BpF71U5Ch3VuoTqiQ9BOFUkg6BUqnmZJpZQqOSPwiuAotI81356eYDuaxfl+5nG9f5xIQP4xVf
fW+L++etvx/kFeh0DKYYD8+XYASc+dXAeQQ5bISOoC84pMWwalrhRNS0u0MPgaMmwqTDL0OO1oeS
0SrYjxHz9dYVUncBBlA8+cVPXZmVZUCtD4HBTvUjDK2mNAoEek+DapmJyGO4R2hCFxhE9YSf/FQ0
a2I5aDUdwwE3pdVwClulvPz6aWoRz6/FgbJ5UXXZXnBLBbc5rysWK0YHussr0z+iTbat0eoO+0co
uWqW2HucAwawbQ6YcyWFF09qYNkfGeWzoICp2v2qGLWvdG4EhaD/j33HdWgQ6J72asHIccsKNRj3
DsFBmzdeF3ELKG4+83axrQVwd/qIpbk1SAbhcHuUw0SjNUhDsnJA3scm0oRxGhdz0bn94TaGxEPV
1rNB0vbVSgJrgW7XgSn03kIkONB4p9s4f5ZSI81enbT6zPDtkRsqCYZeeApnRCXrCPumYR0c14+7
sYvIZP1HsUSbHNGae5a5f46srvUOpsjj/YRfzaBB1yDLOaUzdJzxDGA4xq8OkIZJuV1hTMSwpaMA
FvCBFBx7IDxsvQI0Z/UavqJFGzAq/xOwqjJanI8QNHWc49M2LC3uzwQ95omwj/WAO2IW4pUZtxbj
Xa1UOBOxR2G8IoVrxGbvmWpGpdaV2q8AkMDoez/M4ZbWxhQ8O1WF+E+RU/eDcahIUTlAGmz1ADDF
ZH48F/EYNwW7lhJUSmHIMOP4ucVx9MVUMwxq/jQlS+s41qRMmhj3Q3yEcLOkZVg/RQIJ4WNPUEsS
1Z3CHTWQVg50IpX3+HB8aznJk/kw9ehl/hMf9AxT+Vd4RG6ZytxHm/qpeZ0uQqQThJsjVgUYOipf
UbKtltG63rekk8xViGJmcgqmAF0RCEieoP7PivOsSt00NhfUmm8EvykItvlpKzxYMOlvw2dV8tcy
h6DIvoq3Gy8f9xHguukS7UsqNk9DFjZgdo63OUUem43p2jeIUostdnH1we6guuyoitYDhn4R9AQ3
lyBky4Z6nqI1ROJT0+/BwG2AfZq36VdYAVEtwFD/xQTISyY671RwMjfNQmhzvdKOWCdqtF8oE8e4
oIH1tIis6pCx3/CKPVWBTqCGgTBk/3GVwRSzW29XoS6//+q/B+BCRTy2WeM8uPPVE39RiMk/hUhf
SzA4L3nLqc2mtr1OgvxarsFy44KDH4VXt5Yp754BNSuGpangraB0fLjXfX82zBuuZf/2HSUbruEz
2tuM8s1bR4nDYpq2xh5zFChHdtE+VnkpumCsByo1ow9KH9gadZJOSlWsZ1kRKPvxemdEO/hE74hh
XSPR4gCctiowapR4NpEna9PZod+s46HZP371gxruka8ALQqLZR5PXBCIp5Kq6wUzjXW3UgpTYb3b
Ep51k1fBAROZpunPc5Kmta5AInddOpVEshrmoME5vZb6X0ol/TdRiO7/FI09jG/OTyf8slDfC/P9
gg2n+ufUvtrRF3wccdQDCcewrNqiH7LUONUIsykBwNg9KXCvVQmOm/eOmvSkasGfLHdvwK6JEjm0
WPpA5KHSzb+r17nK1UrSlys8medc/+2SCh9xZbvv7D8lCWn5ViMvcSb5SSzD8SqkFBdXc9hAjRtH
5NnxpXyM9kseTiNu1Ei+hy+0KAM5gziuP4xE1mh+nD692ZDYo7xkhaNx4JG/owm6BCzl0pfWAHym
CsyQX+jgAfPeJ240EjHN5i1KwHuKFRWbh3NWMKMpV/xeuZCTLw2vVj2DrOcsJSQCAsprql5ZyE/c
jwHTVQv8IV6323eYBJB8ntEo7KrmbewuZnJG9fHtBJ9MiMZhZVQOKiejnVnRhARTqMjgwH1Vl5ky
k09XaHUwbeqVNjOzqLR1pCdtW6I7CwJY+6hcWN563Oe6wEAa6IKIuw1I9efDWSFu8/TRYeMVh2Kx
AcVeoiDrZA4Xe5BI8l32AH9QBxmT852+S6d5m0Ghcbdns6coDGZ7l+5etxVDrornhxa/Wwm+8mly
Ygg8349IMK9Uj29uir43B/oGPc1LVkdGcGSPOqbdh4rWODusKyWCP5CDeUGjyI9tLpwWOe0wLocg
OMs+VJRc7ULHqh9WitcY3/ERPodPJ3tRPh3QqK5TD2Wi6GvUnbI66Jz8SNUAM3FPbb+r1iNovAXb
6GeB28F/I8pqRk5NFgmkfGojJ9sldOgkd7HsiXziy69vkUM11fRFPkn3bP6Umxrp4rjJDfFECX9i
4YA+J0gJ2chWymQwmQLvx4JP17IO8mM/GcNdHVKMGP3RjCMTK5WTndfImQNBV2xsfNMuj3qlBbJI
vv7CFlLUeXd2RG7IX1JlGO3iKK+Z0VlQKk4xb8ELAo6U22hr+OlfpyVkxRwrdBM/IQm9ozy4o5fK
m16n1DHchH23LbSr9q3eix5Z+vma8Zjke15CVXoQb7CX42CJQFfUHX/+jhcdWgUJHRRjlAZXIZ8I
abh3ctiASPlBUaloftiyZXfwiBBfLiPCPWPWPdYeu6WfSpHgfrf33n01bVc5/EZTwGdH5doAw32y
vXtKy31FOzYRFZKoL+aFIPGCMj62b5w9MZeaGOf9mo4JqU3B+8/oqsSN9G1vMfYxR7vBD29v2kVw
iZkgWcgnZGsE2tsFI4RuoE09f2pk7oZz1DsOtTTJP/KQXuZ0GOlYdVyv4MJqFRGPa6zHJ2jgIoFr
2nbRwPcBdnLzJCoUlX6pandpCySnLL/6USCegaIIePyxEtMzuvGjyQLDxOb0JeJVLT2/3wzcq0yG
mg0QOi03ANmhat4ZALPuLpSgwnPdY5ZKxIP8PNGGOn4Qge3rt0gAvMLXj2sHClLDauuiSVRuBmcx
60+oMsZJPUeqRbThAg2bltGvqlbhaSTwvXfEwhtj1Ve5JsuxeTc3OOYWdpDOWSJTV5gT6yC6HYPP
Ku93Vx499muMy1qw6bXc6wfZ5kQf+EmMe98sJQk3kBDH1plNig5hnIjZWM5KOSQ2qpNvqM94c86z
OauS82nqQZBchdNTGHgBG3Hebk2W/R7cMzMz9Hx84bmePG9iIBUkgxlJVwISe/fcpZNuR6hEEd78
nill2A60EzE6aV9tdxyHx9EN45HN0W++Kcv6+XSO39rnsIpld27j8eU911Viu59JpQT1WROF8nWe
CPStBvKIlzNCCGe8Bf1km5HJU6l/zugHF/hUZM+sWXyqfAMdXd2Gl4qyQJe7zqhlZsVAYLiOrplD
AW8Pebea8iv5tHVJLh5iQCU4+zw4vHghCdPGtthVjTdP3YjS0oEtxrMyzkr9bKBURrOW/dttdAYc
fnbz7bB4Zd1OUQKxYPCh+2B/tpzYREwPxhaUWT/fzVctJnsoAvAxDUyJS5pOPPf127o7oAU4RgA7
GBDbmpQ8Aj3QlTHoNaolC1Xp+zDHheXNbcyi49IF57H/HK/Y9NB+9islbCuHPQ4shpeUOXP2IiWY
DeUQQvfPN3j6k0q+eNtmHAvL0VxgcdTuYKQtw0ZDJt/nMf3WOuVCQA0Dvr2HO7kT7LfzDvuHR3NU
PfiU/lseysNt4dy9gUH9YgZzBmJSwMic3FLK6E2qrqfJh6i3Y9aUSCNDe1CYREeuI92kbeeezyRx
Q6HBU0YUsdUuSztcPdEMOZPt8wrtsG3leJDQvIdtSPVHtgdGNR0aFmzt7oMx3BeDebw2fJdFgHcV
LY0BxUOQrEAwFDUY3f9RnCUTjmyKXxXs07jv1qcGa3VIhJV4NEwrEz3IchbuF/IDY08tA3kkiZ4M
Uczvg4J5GEpOFYHOVvcVSG/pqkO35EWnmsFLN8D+T5La5PLcCwwkWOyB/PmsB5DL4IqKmCr69Nq9
ohRzM9ftVF1QP2gzEC+JqUWWPqmEkcWQAC665VOUAWAUhCZL2ng62dUVFWyddSc0m/futUYXoCdN
cQJwz/gmnmRiZDscSpeawQOcpAmKX6T6x6r2Uf+dLCS3SPoZvebbmwadwfEBsna81ds6ypRfgf1i
LWSuXOjXv5RPf1ThLT0/wDHVJ++crXjgRaUoUQS/t1+LatBD7jqAZm3Xpbb7ik0XS27tMo+qXzqv
twaKqBFkVJ6xrJbViv3M+sDwkMn8EfE7aFHK73mGNSaPnIkm0+2KIqkzdaImX8EwFFlvzPIAOD0D
W5OPND6LcLWnH1MkeBq22gXkpToeJcLdYc8pTWJl8Usem2l+37Y0LWYU6vnkAzelhoBYeZwLWrOU
IbOb0lKbivGjnaYYutgF8F1JJRB/Mzb4gPERPuYBsNrXbB14wL0VN35mL0rRq1uaAYfTUkNZ3grF
o1IDZ3LG5alLdzvlhuNmOh3w1/URgUUZ0v3enfMYE6OSpuVrJWQRvJHNGqVrMCK86f7zKOKtfhIe
qhRzj0bfaiBG0eH6OTRHlnWNvqaMsCrYxjVZSvgYwaDKGZdk3YOYPxMW2ANZAa8j5twptpHFMmm/
KUdrxnhsuFwlRFuPGOnvp7vWr6z9XR+czsIBmarUKg/DLzqZXEwNcR16blQBq/zv+g0v8mY9mpn1
svd/45EmPbt+3zezMqxxC4Q7l6pzgWZhefLp5j9nkzMF+tW7F+UN3Ps9lzLYn1iByU3dN1i6Lc0V
1V0F71/OcFhiudDqMmo9aEx4m8SR3IPvx4xxymGzwKSBPgxQr7DwZ9IdNSOmwslBq/6KsCzk3bi2
keMQiKiW8Z+eYvD8SONP74gOLNepGojnsqGlDwOXvcH4jRamEZYX5LJheK1KU8aD7TFSvp+rP2jg
xgWrOADM62P0Uj8wfD3g3hxEgKpUovBXfjvPXtbISUpqSEoiu8OrF/XPyYsqfKl3qt3BOyBq1R9a
xfxr/wBNP++4kRpIMegmniWVcTAzKNWhvE2my+O7+eHHS0o7+8f30em9Y9WuG0v4D1guFZRnk1pp
Thx0VYcnOEj3dlAfUh5QWkc3etCE2mwFUMbn2U4crfOclTLn7BBn/GF0DW2Crv3EBNQSn3l7U4i7
QkxHVLkoFO9p3FGVmkA8kDJkW6tA/dXD0I41dNCa5k2vp9s8CR9SgOnwY3d0FzPLoeIapYKM8TwH
4wHnnQ1vbbVri+KxfkLCEPXLD6fQVKGvANuG+2WylesbIWjvNYmmtb3+qqeibDmaD2iyEvKeb6F7
dH/PuKFYY/S2z9E7vB5C4a7BBtrQqBYS+Sa5mj/RpHp9P0aEe904l7/Tmyoxm+uW2nz29FZkzW4f
Tp5UUsibMBtjYEev+rGtkpw8qOyFuXX9xJzs3xv2Ww4mNgjvWM9vKaVjMY5Q0QkkLQBd79SxjdOQ
Ix7m8OLNbiWa0lFWnTniOKN9NfWAmvA5ty6dTE8lbuc3ouwrF+cPpeJYsiWAecmnlwnQogKkul6s
rlCqS6ljz2zzVsugBO2XLvcWZFNnE3xPpEltxWgh1fILLGGYfNMXXpClTK/nrLv1ZCvPHQ2uf+WH
S8cbdk3niQ389TdRL8P/JFux7Pkx+Oe6Sl2E4bk/YedLmTogNIuwBrhn4+5qCMo/73JFFFcjuNC4
4/kmx6YYoUoq0fHHF15xaq875JWJy6JteKwNpS473LcYFBL+ShtkZbR87JvoFi/GzXaRI2PcX6Ji
E7adX9Wio9wr9gpn7JvG1dJL6LT4VFmh9dfVC59YyNTg/iI0RBRq5SnElDZkpOpJ9MjGx8GVdjrH
I35kn8W03oKMHy1CWYfe+tS5tGIh56fvuhVj1MCIxe1emx5zKNLx/a6ec6lrqywNm6o7MMCMxkPX
T+pQSV/4EmRC0dyXaXMOV3oR543CZznnu6Kk+lDifSnZK/2JkZTXW7U4EKP8Tnj11yrFXhvCfxa0
QhgwoBlae7M7t29H4ORCMv0+rpaod9tLcxNuS2GazdvbvKPyu8hgIzMA06fEHMxzHVl4mwVEmtc0
0k1gVAJJn/a7Yv0rE/nXxdoncje9CU6VxW8ZAzMqQwoEavUvvq81kv64rysSmfU27OA1fwqKvlFN
Di6Ghn35rwqXxlAfPlSg6yTtP1ziQGcAbjvXX9Xrr91lVQ0/5z9uey8RQ2zPP2X+Sm7LkN1Alpkk
BowA0wfNePZBBuOUILTXZd+UI21R7zCh9urbzgYLHiCWUdKMJkPja9JUifFbZz484nyigNOhFUvW
2ngcHOkuyXapR5D3SPrEg9u2t3Wf2G3Nqd3zB93MszX/LI/Eiq+QWiwL87l835HLuCAkoFCqyJRp
y5m8aCkYrWuR9bVGGFu6H28DcoFDHL2sfR7SdUOe/COHpu4briC7dxdngIvytpWjw1pW7JRWvuG4
wWJx4fok9A2IJ8DN9VsnUbvQdQf92cAW9Jl45ut+1bWzNiMbedqxsgk1AcCuFWfBpFzBudxQV2Yk
kZKVSwQMSRX8d6k5FUUf5Yc7BxaiedZf1R1jWRQ39fxpfE1SrhudvqR/QJ0+Gf6fJ51M3Y8fmpBu
qtHBRzU5bsuM5RH2t4J4bLei65+n33UnBeFfeSZQNA6JNerYNvy/sK0R2FfF7DME7zaAuQGGhPYd
z89W90ohaY8i5KEuuW3NNEZjiIHunyqO7zrG3eJUd45tT8KiM5U1roagJsaIuZmK0JhVUNu7afIX
0l6LjWs1zKEsSPRLBWgYi8A3zA3WvhdHiYrF22V4DwjlnkmxoCPhFhm4Pp4aghi16GkN5itIpTeb
rBbGE0Lc+uUtmhxZO3wKqjMQSVjdST7y+i8/Ibz806/EuWpiciDV2OES1BzUQ1SZ33ArywmvbJWm
qaI2gbDP/BbypqCvEej0WkiGFYiyYol3aJvOr8Rjg7nf6cQStCqtoPwu810rHRHq6JfeHS2eReWb
02svCxpAkuppekt+e3k9Re9TT7Ef7OrlgM2hYO9yY+wYh53+ALWXaofUXWmfHQdP1NilPyed60Dd
F3WioozAn1u0LrdTgndKXkLCOyheaV5dZdK6kk+3Z+ClrlvyheYOeu6uIiao+yM2yzhsz1nqcyRo
5JLiBFc1B9gZhd+A1vFAaIPlL3HEz8fDEND6vVnFHvEyA6wEl5p7/j+cjv+4nV8WGvHMOcNpxpkr
nZAFl2RT9dqV90hFwrV96jkwRpgtcy47G91ZBTxGcM5CHTFiRtbZwsGa11CGgQRIzK0NPDmxe8H4
QYJfpguRtA7W9Ych53T6hNt/DgqX0KKCKgvgSp3CB5pXY7BVs9nafrElP1WAQaKscocl0bn2NYZP
ys+qgozkN1Qt6zP4xp+exV2+PVijlnU+PIHqFHrLRweWZr5JuAchhiGFsnVQVRm4pnDF3RzQ0te7
m+hZh1WJOBuVGdDIBvoI8czp0AcNfCGq1tzp/lum4AdwHrcbAAlaMsWIKRN5hgZrsl2B/BF0Bcdl
+fQJAs8hAygKF77RQcOU9dlJ4onyEP4C9SMKL+AD53UhwyH5CD3bBAMeTc/NdmOKPA8RpR6TGY8f
s3CpOCivo59o7NLUsdI6+K+6BEQNVO6jhaWkSJ9LhDsDwIX9jZ0GtGnnvznIFV++HajYycj1hPax
gX//ELaZkczHIZxqyRRQnffu/tPU2+A1P4K9i66Bnphtx3r3VAw7a2EdmNeIk+bjPc4Dh5CcjAtF
tznMuS7SY3KHKSwJyydDY0+B4WUYtSrl4Qx9wHKgyVmgB1SJhVHUaoe5IfI6mVVWT4zIqUjxb9se
r+ocoUdX5ZsBmiOjSJIG2edqFIJb/eD0QgjVZb7cNMyhrNrg/ocTzRqP0saJlZbpf4fnoLF4prVK
j5j1QQv53bvg95xhRuURmXtN656My85S6m6/02k6QtP+jM3gieO/lOY7SH41f8crd3PUJYEwrcB8
MSVWWmAeP7D1gO0RKYqADWU3KDhEg4Juapg5ZlG867E11SJSWXsAFVFO/jb95Uoco6UJ0G1B7xU9
2ZVqSkE2r/d+QbReDBEwEcykTUVbJdO8T/kkTUBaI2hvnvOb8AVNih+8EjciE34n3z7yy/NUJGLm
R+HkVOuUoZ9YQ1tq94L2UE4IrgFsZ3RlOuR2UpVTPFXFyhPrrYZCDdOt+aDUp7K5LtVh5uzlFl3O
NjnQNnUlZnPk6r8Gjbczdw/V4qAsLbA6f58WAciPRV9SUhlrtVYt0hTo5FNqfzQ6lgkZT6rFh5lc
tJPqwum+99rkFHwmdminAvBbTZcVIP+kqoSLE6soiU0Pq9+T7jWgHHr3phfxCZBjqRXLMrFLhcor
w7zweP1jSdBIWVzaoP/4DedMdaPa9QAXzaa4PckoE2ZXItnqfC6QFHgsCe2PGcgFw29AmyDzaGrH
rYkWO9Si/hOYOOwaN8zZ0EKTbC/wJwvANGj6esPl9xU1XHTVKCnlRf5WdIjFdh926CM8hmDEo33X
NQmxn+Vfp3b4xr2iNkNTXVFZo250X4p/sW7quQgmWJNGJQw1ryza0OU+KheJSigevLx9QbH1qNd+
clBBQi0XVin1wG9S88axzA2UIBaob8RnyaBSxDc7KfDht9KMyr2DZHfG6XbSI8GhT+oWAztyk7UD
wSHcGHGoEKkD1AEATmMUF4kUb8ama7AkhxzrbAOKsQHuO6o8cx9ax5SCet3IOkqHhjBj0qSPEiIn
Jm7aIcFmLK0e+f3vNq119u7jCXkvX9cikkeR9EU6X7X9bYdwXnzkTyeh1HbolRweNDVeZEcW4OeJ
FfPHV2GXAXx3dsfUBgoCOSfKbD5bk2HLzzhjq9us+cATEdJv+9BQrDxHMWVz7o+7m8Btq17Twd5p
nm4hVNNunwt8xIqn/mfLSVlibByPEpaLxsrBigh4YXMlnw7obe4eQSbrs2dFuw7CS9AeRpglm+BZ
zBp+faMJbt+9JSRI/xVAX2GfDrCcH5+1/wWrnRPRCJ3q2WTi3lzibRjXuCn4Xj69YOVD+ZFNNl4x
JJ5/2Brc6uXFdtenEtYZDA++BhqICc0tuvWkQEPx7SmzrHDjNq6KR9BEqKaHBOGdMGb+nfRJ6qqv
8vnlqaH4HKfkotpQ2oqrCaxg7AolSl1JZkvN8Ck7mKBQ4egjvMzTxGzpHfPqjeo5K+wHsE49xE+T
iN4kUFHk/zNLUHRlYQ18GtDhKxsb0jALKWejnt3rpZkvFbaAYDh4CB6jzQJx0uOUjGSuXM2FsRAD
FOHqENfQCVYizT5oXK6FCHNZBmV09vSdfLUXV+TpqYKIZem59t/oCM3SvZlWbtDcXc9Tf2ECV3rP
1JBu3cUI1zmuHGchgeJHiaYbbIKftbMW8srLbncnDnwu++YOp8OQd/avaQgxby7vC8Squn+cJlNH
Ne9UaVhPMgtc/Y0n1VtKvnaCAg7lBxu+OgkQSoTL/ncHKRcvg2rqIkxgr/cpRRr7pQV4w2120n3F
Fq1W0G3C02/3JsuogHvNm9Iy4SjlLXMyOOLJxxom7nlOE3YdH9x/TWPe9yJWPWSwkwYEOEc1sFgF
TamsXGzuAwJik6HPelW9VUJX+kfVlRnIj0W58/b/pkTeg2sv4P7GAB/sCDdOMrGJxN0EO73F+PkZ
NC+dRasrQ9FzUJPn+TgEfV43A2W6ZrHD2CyM67UvRh8vTj8Ql/D50TniVJCtZFcNv89mkkz4i9ZF
QT/BUIBxso4GZxDHitdCeQWJ6/cW3rPHgYWDt0dcph23w7IIhJbE3bEQJwQsmuvIoZ7b1PaxzFIP
IK6fI2w8BBlSnd1sbtQ4orpSyXyEHJ9dJdSkAtcMu/CCnCqhRMqDDvRq/cLPN9d2ph9uEPGLwfEk
7xZm7sMKRxqdfKuqRFtQHpcaoXfPMUqVypVLUkB2pqM6pb7r2T0PREEsxodlWi5uIBDuuqczyO5P
IeFPmF4HOArKHpXlzT3MqF3FKlL8geVhTloDFvUhBl7vVa499Pr08SAtXtHBqO/rrpaVdnTSfNij
GQ2XXvwYhzcK2Ktd3zkCiQZVsk1hD5dXFtCdFhfA8+HPQj0uHrNpfLEvpfseSgFykoRAwQ/QFwQ3
x6pSRCyRAyCQuLqvFiNiGvCoY7kD4uj7nR4xG01SuZgo0b3t9L7kVeYAtHtahW9rpGsmyC3DtJN9
Ie7d00xVCNEaUBRtKMDnAgeNwBRpWLYKD+VWZatPwyXGH77RkBSiQRkc3F72saJvch9EiGgWdUbN
H9Rf/DkQuIHtM5nhzIKIP66eRPAIECzfQCLjFEqUMx0NngiYrHhui5Vu2JVVP8nUCLUM7o9BfWVZ
O1+6+o3TWfnj4XCoPASFQZkOVkdSwKLnZfp/jUmLuX8DEFDp3iZieXIfxZ44cHFnRuqRFjGnt0AY
trfx+jUMg00OkpcRDnMsWkrKW6du7KovYDeZXXBOqzuXq0pqrndJzP2w0E0ZJAXPQG6eDjOnrOyN
1JstWHuyioyOY9mZ6Xzyj+hyyfmnVF5yP5R5aMoqzwOOdmaWXK7k3arAwOc7Te3cs7bWpFfLI5op
GIUNmoC3017lD7f4H8cCco6eyi0e7oIuN/To/h4ebse/JxdKr8KYpSiAkKbIKODVP9tSGmOf9uzR
6BVmMe9KLS/WeHI3XXxblso7VSusst27j+20wlQBtruuXuiEmRp9nFTGsjaLGC9VSI6DN9/DdW5i
1ScJBu6SZh/2CX7uGi4jaNBo1D4qNC0e6eLy9SfPjsAaPr60gOnjPJCGFqdwlSZYij//bgk9WTX0
1oLOivL8dOkOpY6O8Zgpy9FyKGKRigoMY6LFnBqDTo5MO0B4SuocJ0tGZZcuZbEU4FF/iItY/Sr5
joyDHe4sZW+xeCpJRnuB6KAD6J9pAlBQEWMvFIk1ovkFTbD6HFoMkkTrroW9nKFrHhS+WukwkJqw
zVEPA8qvoyfLoJYNoLAherBwdfu4G4U7o/dVLab98UNP6oRp41Y1JGPH+FAEFYTQ02hgeof7UJEM
6velP/irTek8tW5ohOr2B7dXoCpAlRnQsrs54PeVDVt7GzHr5ThQR9/DrM/kIdcBbN9Jp5cRZrOC
YYGHa+oIiJWdacOzaGjlNp7nsFHJVj5mjDESiMj+ywp8h0lW96PfhErPyH6/4cokzmVfJPXd7Hyv
qsleDxSDe/uZYdGlxzLx/v0IBwe/M2Ir3WSkjUi+MpoHLJu1X6/Gyr9Tu2U4Bn//wo2pYnrdZuv+
6vPsJFokwoMuLI4X8UPNKDiVBbxTyJKZ9z/BzWi9IaY9LcMZOYZNF2cQSpSwKsErrxx7MPZoZfyr
pe4k5hLnd8b3GfrVTk/IViyDz7F1+qS+UoWKJEqRz65OSrDuRA3rLowTepjXcL40cTJwOKBO5rz5
7wRm0ct+J7zJTEbegeTUMHZ/u5DGCyAi48VnuimFe+f0bf4lUsdBlLF3wld8Imicogk1BYF+Gy8v
9PiuLESea1sB5iiUu1uMj8yFWIfVB9/bzvcDEjpCdeIzK4/VfajHNkt3MNaN7po8LpifWv/h/POw
E9tPr+8YtS3Za4GXqgfkwuFmNlj3bm65pvGgpz97lEB61IcSGgrwRpP0aFDSZv60OGvTcETiTRH2
gUL/SkvJ7M8LwYtmOTmdrNDVc02r2jsSVMW3LccQN8Io6sSUIw5d4wOybV1faT273Unb+4GifCe2
1TOvoNj3HKSCUakSy0i3htya7vwFKHbdvF9P+n7lp1pxz+8c9TIW/m7g1+i4o6DD9XiJeajk6XlW
eonUJzsgS59IRjKCNBVkB7M8z3dnHRm4fzZ8wk3779anMbrgXvhl2DY+3vjR56faz5VjiZ0xIJSI
wJen/Jydxhs8Z9VNGBsdFFB9YoZf++xi+oKYADZHoX/c2q71NoWWDN7K2SK4Eg9qAla9VmQg+sZg
hLUGi3R1lHNi/y0B2A3AeV8OeybrRdZw0QyPaSClvWNzeOrWDTu5sNwXo350vS9lWWu8nZCcnmEp
pX93GTghBaUdrLVwiqVRmRbQABV0Jm5Vh06rIfwnPGeQfZawTyn1VzhOyNvk6m3UDrJgxUaVORBE
lH224uIKbVdtrNNwulizIZanoMKfZZLSTC6Ty0rMn8WPnEhjJuKspdu7+IVBJLZ7RJKusY/QzgRU
+tKoFsOJfCz0x2vET9RY0AHoaynvtuU9UeRDWXDn/mFFeX9bpxByqJJOetp1QomTTFTX+yFXvXPn
juK+oCDSSWzzgFAkpbzrXfn93qkdFj98qWjqytkI7t3gjEKB9iJ7RJpRv5gB+YXwjvZZ5J34T+DH
iLFXD2Kqr4wCuiY6vjyJp3+J213lF8AcUCmACeTNiOP/Bwv8aLgIkCKEg8awYDSYzpQZPnw9FjSn
uIM/2yeSbC4rDJh1dn9vBj/ggVsWmfQd6Ygf2i+1YYTuK4+7lewdJ5lRcMbq3hDxp8eIOVKtWF8+
PYWgfA9GJYFt2c5ZHrEOaC9Z8nCEcUWHe92nuj9b3WaKhlgXrk3lBmGSeKnkdiAOxGZLjmGpBMlA
lZz+HpMIfe1jRKGfbFtCV8fsJCzd9xGdsyq+YySE9/RvejcdqeVXUF/MxHd2b6zm2+tP/9HWHJEl
4zpt+1mVA/LvJJhU+6YokiV8DNkNUijGSb4RNSIdjlSenmIS6kLPM4bL99mZGTvDdzqOzoUrHc/k
WRuJuyx4JCyejuT89ZxYtADmJIvN6GbfM5deUdtXtIA99IC74d2mKRH2Ea1wUfo74LZT/KM2risV
yXCPvsbwMr4iv0cpt0rSNDxL1pYxO80PByeRDGwLkJIrf+pXXIs19QLAiv7qXwcms+yOl95eQJ3O
BVuqX/0U+Q7NlB0X9CfYTMvVHs2i1B3ZhIq7Tt43glWjMtoKLWxaglbl2kOGG5pdtAyH9TuPPNv3
rXqp66uP7D533m3m2N/NdaAF3s6EQ6JEaetzlSFL1MsDYTtfxt4UMuQcbLsaVwMSvKv35qZEgthA
mOzAT4b34CAPjANz+XA02//PdPr4AkzdtAgDq5QK1u/7G6fADcyK7bVj3cabCo4mJYq3IJxzcl/T
rM9VRJ0I72aXkMixLbk0MHy4xyYmhmpF8HLfEsWQC66qBOXMCpCrCKHj9qmPURtUMu3N+j8cqJDP
UlMkwZTvQGKJeGoqvIORfmkczkDwMsByqiTz3vRVXR+A8lzF7GoNAhnYrDmQLe9rCplmu3eDBRYa
ukix55Ebj0SZn0AirqQ1wEJbET7C68RM2K2gTpge3TzD2Joo+JKSD8W+RpkoMYXz+EDgRJUN8uUC
5a4OO+fhZ08Nk+HFjDJ3G+OaqSpmcCaAUyyLu9ofceqOpOZjRhPB31g5gi1V091so6n5MX6m1Bsy
aD5HALbcY55yrimBRq9Awl3vM3MycCIfBQplVNMfsCyrk0cu8J6rnuZ1XMlAyG0TrJzVDJHTDdP3
eCyM248huvHdkpI5ZmqCh8m5sKdnyaVJy7LbzmCOaM4q1CJYpxM+c1O6WUgBrs9jQt0aSz4i/81m
OSaqEuDHmM/g31ONE8EtSbJht7+f3gJV4kVz5/XoCYRTB4RK9vmb4T4n0Pz41GIWZjBkxkd9zoJI
zDieAPHCwwZvuJKFFB5fQw2JSofC3kgN0g7zmJjN5CmQhNIizZ2ded6rrIR3DrcxLhFYLOMJLRPv
SS6UVKC018MzkSwmd1fUMtub5Mkiw55c082Btq0HqWbN3vg+u+6ACxLhoSX17EvBw1gjsqbYuuOY
fkH/TmSfE5IN/se5ZuYhPBc3SuqywfFXQ2BiLchUpXLATlnd9U5JvDgCOjliSK8QdLEhy4YG6TOr
iM4Y0S3Q4C0mYiZekR7c41TLsKSxaUaohdgXHuiAMKWGjevyl/QvYWXL3H2dZcOERG57E2mYFnDn
ZiLWyUiJc52ixnW5u2PWOa4djtr42tAW494byOwBieqI5mM7+SDeE9Bocg7x7gWMUpkJNvLqEbMt
den0kHCqZAJ9DhBjG60gof/SBsqKyrMXYHYGOhW3bICVnPhIyTDElRh0VclMetVdMx5frFMI4rqv
cj/bxJY++LnqHOTwsZ6oAjFBgfsXoSbHIIkrW+MoE597YJQLZ0WVIO/yXZHrB7tYkSlgDr0l8bg9
zhvMYkaRtAev48dog5UeM0/E8GkMOXlirmW4yUsMToH+TTwStyN1vDCQppFJpM9qJOhvh84Qz2H5
4ysjxVRMYSyYnj9TPvBNVLH5oyXgA8V45Nh6G+vSrT2EyFgYuOrZAikAz/dVEqSFePL98aZzZMmO
VSC1dYaoYN48enbWl70//QWZ+DhVAVWhFTqOEN0JTVsoinFRAVga0O811iwgifTlVWaJUGOjoGOl
Ymd4kGQw88XKtT1rPIAB5qnsPXdOYiuLjJBe3+M1YBg1xxMXYhiVxEv/cG8kwdvVUjsaCVSSQY4B
iX6InWcXX4cKphdZIXrS7z28kDsiF23Xz7S8WNeuSdvf6SFyp93WG4taj+NVUTvcB+MTvv60HBRX
31SfoiVT+yoHdNXvffYFf7Ha45iN1ILGN8At76Q9kZJLMH9ETNgImRbmuueGxW56XOXoK6V9yzg3
WMq+Yq4yZZ8JX1vmjudGNOnXpXxH++NWe1UaVZyhgd5U3YoQa+ay57LXei9JnqHvkSNvTdGxR+rB
f4W8QUzincRYPtEqqTfPLRfxSeUucFam2aejAxMApaYJujMH6v4qg5cGtHK9CWYG7zPzdyNjofIc
i0gSA9yNdqSLjxQrhyIKdPQsTMCyelw/d5oCST563/icE4Yttswaml8KZsrXXP9mneIuTMU9vuvH
MMTbZ2NMAs/1EAq7oU2uiCAcL1rmluBKyGqAM8e1KJhqFNXm2AFc3RwBVx4C0hnNJfBWnZLvs+Bt
oQK6UUiBLX3UT3BAjU+X59u7E5Uo9TE5kmNH83URwra+3HC9bXedKhtMLFIealmGlS/l1jLWtw96
2vprYQ+zFQOmUTHzJJj2fXjTm0YQLVof/SHsFpnrIG5qPMej6TwaPe8RkXUuHRgHvpbK4a4uvtr8
eVSoDu/Ywb4bli49UgKFc/fBQIy5wHe04JsDIKFnTpdJ8aHUc/ND6aX4/9zN89gxU/WwTR+QA/VE
CkvsAtB8W2q/7t/ZsZzkms74uUnXYkbiTQM7qKzsaPaLe7OIv/EAf3Chgj76RY6k7iD+X4R8SbMb
NR9egoHhK8dZA1sVssCQASehbj1CcJRZxtb0J4RN5fJbRQBcX8qJMYwROyoYXGXZYc9e84LEroQa
StyOiMAANfW8GDcspNArwdAG7uhje2NHwNNquD2Krv0iEbY7WKuJ/SdFC4AzWYcFP9Ic3jyFl0eD
XiZ0hwqjKz9uFrl1VHEqQvm0WmKtc2x8d361IIx2cF5NJiI2AEru+vt0FKh1CjPxsD/+4+eI1Ivz
k7GfAnJHRJONI2HdaDkHNrGy96dgv1STgWFHpOHZUpL1sOQ4JRpKIAnY80hvHMQJl8UiDqdjUnXO
zcW1p+rBN9G9snmjrDwd8uVAK/QH/htAACIXjZmt9AYfKcUXp5zj1T1rrJhpkqegjsNmMmCYFWm7
anrSmv5FTTICmvV86PYcYrmXDPGcJJc6LC5DE5mqy0j9rtawnEdMoi3IQbWGqnI6fJwSzl4HZsuU
1n+MClQqqNzPgHAAWXgeW09apteudvS2tCDo1uh3F3kjl6lj2dF4dyVOaRysmBEc4ExONu/Kh17B
98nBxaEyfimvBthuAT6mOUPkNAmx/hY7c8sEL+2g2RZOTQ1cVeTfNm/9DEr3X5ih0KSBrLdK1DSn
DoSzGY9daruY8rw6iWZtF8+zNOjCLGmzDOoI5ErXU9aD2Ihs581wx0Fy+3csjarkJNgDJWgc8Bmu
1PCGso714L/2SvFEgSyah95PojPWUO+ecRunDCT02mkBbvvL0hcyK7Turb1rrYUYhtz969Gez6ga
YsvU9cruDblumzHN3x+Af9ZYiPyJ2gDr0t7hi+auu+YUeo4vNiZ5nd0yyDuvXhz2ltu8mYtNq85S
NEWf3nao6Lod/KeZs7U70sI7kgalZrbr6j2WcU5Iawh7sFvD4SrS74/jgPLBJQgVjTJwIhTxXueX
dzHvVswPXf1bf2z6LU/5Ybxvr8Nnfer7AjR3O4xajHZeU4Qi+yz4vwmsBIk6f+AND1rqhheyGwYp
P4r4E0zqu9DC+B/gnTnHk/ED6fz1QvBccu/Er8dkxwMfoNJmK5sV3uiTNHX9DX6/ngT8Lr7bPF72
Nye3ECuPq65MxsSUVBHPe7p60oW1CckuPaG3FFdcWro8GrdGZQ+SbCIRMWark34qG6OiZtXyOuXY
KGx/nlvReRCfkulQG189E8FkgBRnoHee/BUqmRBTfyAA/ZEHzWzVRTt3nEijmCHVc8vnZK/mKPDd
7daxv0s6u+QM3lwihCnA6Q04pLsHQei+U2f2PIeda0+sgF5ekwBK2vu6FCf4e5V2QcY0vq99XJTT
a78a1ukqUo8zuqZHw+CC0b55d7afiCMiofQIm09EYKrRYBe0aWH+ANGC68yvDKeyEh1UToydD7BX
1wWGMg7ydLYNoE5FbqgqB0tZI+fBj/lHsD9pw66zQP9F53OZwFLL9kwUdt/xmgDm/1P/0ksgmd4j
GBv7xZSuazzzJSifB3yU/Wwuw2bEB9DmExMaheR8H9y25fF7/iHd8aLT6zHquUQmsfN1wgyMvw6e
FYaPZHW0OQ5so/EiWvWBafkIqpE4Etw6yIrazydjmqyAmdXE0fr45t7i6fCIoaa1EfL73g1T7DHB
a2yjlCyC7eWg2LEyGscwCI9g/b1sJVyqy3+M+ieyz+ODxq7Q57/EVhNWTJ82jUOPLfNIcZkxGLLk
628AoxXNUtcmHxOhA5/S9H0aPDIdztztIl69AZv+zpZ2FrkTqPuRdRvbsHMa3IphertVOIv65yAF
9c3cxAds5etnKajGYQCqkK/ZDpbJymADJKze3AhnEIjTbbzpoIKAlDIuX3UJ+tSMGYyImghmxQ2D
joOG7nUqrLwXws8W8y6ubQlNdEgOsL0ha/+JQ6q890E1r5VX4pf0dcy1sY7NyvJ7Sfe3ZAymtW8b
wma+R+JhTlWEmodFOi2PWMKXaejGKYWouK73gCr1vvuwF7ScejRj0n2rgDswDG/feb6dTWbb3J6L
xDOLBKOiejxktYpI/jwpPtvBFYXX34/JLJurMepys8uvwSu418Olc+JAhMhOyqHnb5ZIqtuIsATN
JqzjG6bTI0jnJvB78QpuQ3VHxk73rvidrhxEI1a9j3o/+YNti4oNFvko4ErZvNmnyRbXmCUBqg9M
I51FYl63BRj5GAFNX1enigLLBjJf8ignoXRW8iOauqhgBjZeI4++FuEg9WqWtbVM69vPbsGTG3Kw
WgyAO418uDSYSYbOaxk1Gl+y5Kp5nwPYjLZEXXiflvafJAta3A8xlof0K/6U2W9VyHzF/aM9xP/q
ACeE1jjepqjQRINna2xBqSHbQu1Q3qIyMKpLZARCGbCbucJ5AekOjyyaet3uPnHzeDrqD/lr4S23
lTN4R+vV5Bdqr3SKDEWz4eMeC1K1Wmuh9m1JvASRZRWuHa47HyKPoyQ0ZwPPrL4yk9hjn/6rf26G
z2m9CILfg7jZ9mOlQ2iPurI1T3JEgxRvobPsx9sT5///EYs8E/TplxLHCv7vlT3JNb9ce4fcfX3n
gzWK/rKWioCJ3Frvg/G4tH/fDuJMQ+VFjb7i9LbAyXGw9rXdjg2uc6RNsQ6R5ddZkXv+BpI1hZM1
4PV2wbwbBD1GvOqiapueyeCKUq0EdGr6F2gHIWxYZ/OSkmlPfTSfjE0sps4T4u99J28+uT7PblzB
kIrfoLP2dFnk0cpnCaIQI+g19hl/tznJCrSufNmQKsVYNvPAB4tFt4+swS0AM+ykbYbNyapn/oob
kzCg8Jw+nLH1aB0T9MwdOpJV0wcGfGxyuGk2omwDHGumT6K4ph7uaZynkQKaFL/61SSGF3iubEJl
hQeg0LzeDcWItbEo3iRgfyX2y290naMsIeUidAxmT/3bi67iWTmSVn685w8RMSnP504xNxxpwIyc
KrFJZBgKE6EhlhLp1R6xu38TAk8iBDpRc3/T+yUmezRB8Iw6UVN4dY7NYUH29vgjZrhYnxO1wgZh
Zie0+0bUR2bT/8NMjVDZMdxCUDChy+l+5YvKVRvP3odoItzgKUJYDgzNYx0SDkTiOk1oS4dbabHV
ncnpOoQYqrpJMJ9BqoY9CfDXreMyBJfKkuIVIM4hrJxJPxEfvWg5owRFVVy/M0cl1aKwNBL8zLoi
EMHBZJamSNRvUa/BJoxGvMsytmUhqpy/06bPpTcJVlRHD9HVc1YdB0z/b33P263IQYXXTaVy29V5
IHuNM/SD8m5c51ng/exaxRAWLMF+g/BriF8e1gJfWe603bXs3xo2Ovvucec5BJ0hL8YAj3u4aI8a
64fxr5xgusLyQoNRYT/7hZBF2bVwYCUP14FZXE5QWcerzgCJsUAHEU9zzlLHkojsItvf3H0YYrDV
54QXaZC7YSgawmRlPRmRVsIoUThwECuiBO6snRJH9w/H41xeElwZV9YbbGsZyYwFpmwMppqH5gqf
sIxkmg5OrAMcMnPR8mE84VQcZN1vDif/3gwOEVAleVkGGxO4rl6/UUjGoNzCxt7npy/57XIFRuTO
h62ihTyWdmXIotR52LIs3VCgb4yJYMHvOKllPt6fx38TaLp8O9JJrFQdKZLT0FJhUAK6pYKXSKSL
yRJMDcasJ/XybX1elQQqMB+JjxRvQI2z2Lt/uaUYImUdt8XgkfsMXmlTwZXlukdbF1+/LBTeG2AW
zPRfhGf3oPzC681Io+GKJ887FI89MjURC5rSsuCK906Ie5PwyyPrTgDQvDpLHK1I8SV/nrMwmxNr
/mZNW8GL/6mBhjFEtzgnoo1pzGPpUso4b0CB3FtiPw32HxbAcMbP/a7gk3Lihw7Srm7iCL8n6RE4
GZpMPhqRnx8FnGON6lDQajdhcPR8iRfzO4quK7R/NIpVvDLGZcUL4qSYMc91tP4vE47YXw9QIjTk
As3/LVpgxJZ4EByY0YJqxRGrlLS7YXUR/9YyqQidvD0YUA7bCEWYoAEkZjpfESsHtKQg6DNKoppV
dYeGERR5n2mMksFNcX9b4ZRykX/qsQX9rwKmlla+OK0rOuaaOSQNu69Iwrz+MDZgJqP7k46tgjdN
vhbahyJ1kXhDvdq3R65y/jqi5Ag8TfeVzJWvrum/PCg16yAZQlGth/oK2BU6mQjN7XTWKNV5fd7Q
kAtlojdWrBHvp7N8uWCf509lbrJM2d2UDtZ1qaYLd212lIU+1YKLKYWCEqK1zOj/LYbZ6RklcwXP
tI0PEwiXC6Ha6oGLudb9KPTC4DyNn/UtvfL2X2ERQppQO2r5aytrKsVYvXFOfN9/CPAsqB7QTmFE
THXWrFo9UBMZAOC8tVR6r1ezK1BUJDOHne8G0Prr4vfzN5vS5KVsTjPSvgLoz5Xv9LxPXLCkJg5m
AkKy2w29zGzNaXwL7NqeMFbfxHLF90/LD1gRrsGrs0pC3BgEBQNAHzlsaqYAlX1oE8ZJHR56/9Zg
laLlXp+9iRNXgkI52pDN+nYE5za/+ORTgGNWedCc38yYIZ6OXONQquK8KgjFuzDB47GHQpAnQJap
SlX688C9sh04loEsvfx9jqRGoyIW39mCnHkPJiPofSKxlCmMeH9RDb7Ip4Kx6FIq/7UBJHCThLDu
UOYk3pUGhx2BPdE3+Ocbj9On4VaSm4IIAzDJoXZJz5KRW3oELqEiKCE/HNmpptrS/WJUrdjcKCbU
EsniW0lq4sHLQF+TtQzR3UNXMSwp9c4RfzqnsnCSGdl5KwPVLA6Wr5UD89Y0B969rYLfQnr8ANHz
3AKpdRDomGo7Np+8qxV6jzGHdaHqLw4HNy7unHxRMuXLiT+v5JLEAOJcvzaxvCf3gkE8dfASmRMP
SKAW0PG+R92ft+ieqZyTX3pGhFdV0H4sORMuYgVItk5hbTdh5Hn8tc6pE4haTYQLDIc+JwMSm9+E
QdB9yOh+HWYF3XaKeFmWjzhT14rnNa/zEtCn7zyNs7jVcK9KjevTMVa41s5qRrpdeb7oIA+YTrNs
sj8TcBGaMPD7zYoK7LFyjeM/tAn85GZOGPiw3n85E+l7EQTtZDzpHlzMgNBll4efaFx0xoGBrJQa
Dj4POTUV5XbT2sBrFn8YFU8pLxJlERQOc6uAzmW3LkpM0ZSWFlUbyeO/BT7sgEKnIyGCdWPBTeTg
7ZGKxQHeN8DP6UtqPotry+Xc71UHg4bdK62a0+uJiv8q+VuJSuYj6m31C9YbcWxfuqR0TDhuMA75
mYIY0KxZFBem8OK6KO6WtKklEA/l3Aa6vEqGdXXrmD8fgq7K04LK9MO/HRNMIDGEP5Ik77yeBcWW
BeMg/nlMNpBhDFr7DNr+5yjDaDbC4pAumytlJ7/lvSfx2s+SiejXMprtJEor05d/RSgb6SWzjBSQ
b+tfkh0Rx6b64gvoRal32it+BmBdhDq74W+ix/1frBYhqXUwreFZt6zT0LACCcuQt9ENUcIcpzQw
XT22szCRVz/02KFrOlTpjRjUr42z5fPTZFRTdr2E6NFTg8YfvwmpuUSe1pRetLKJn97NJ4Bmnxa6
BOkfNay0cs3Et/pfKnTxwoso9C550TZ0/tPwpbkb4EOg3H8rnIHQclGp/C20BYPJMReW1HelyZnl
pMTiya2HNDWrqxNRE7KocmOaOW8S87REVGa9ZZaMFHHGs9W3TjPRoRIMbCY503s//Yl05dkK//HH
5eOkmUKFU4GZudDsTtps/lE/QSHih4iwqXYTsYgtDACXT/VahrY6ntkrrYp6Jg2TZAdwyIq45qRe
L8MLCTD/AZBQW9tfVEKU4FG/WRtJJkDQt4UEqc2uK1DTMxO9TorJHXHBVpMlKbquD+Ypudq+XdMF
ISJec8cvZN38NJNxnJI+LuiecmBdeW13gx9eJRloWEGJzqSf8Q4FXJYB2eW7cr/q8Xo0z0fPGQS2
636NsPkW5h6SXrDi1dlcX77ClnXphIkVYGegndHUVih5H861czRRqhvznMUKFcv+2L1S1YYBGvNB
jHejIWH0hObwg0NfrMYgmwKTH/JzFgT3zogoVjYF7D/1idQfVLRe0PCsaKqL264uNzFBs5bZOAwI
J7113yzsqt/hEN6UbdAoExYxswax1Di2TxQMytugL8r4Rpe6TblPn2ErCcj6BCA2C9ZiujtiiiOK
+7T2toXSZCE+K87rVVZhl8DgGd/zTlLlEx2u0g5tmJn/oLjUJAgxwVxK3cnVmTr+XF9qXrxTe2nF
YRl6fpF0YYOSLGCUSFxmA1u1FINfuKyVAqwU4ORnpl1DqoLCb+FAf4O8SzzPZs/TwpizU2Z/xUKm
lTm1+h+6jLdywEB6PzjiJ4t8pA6egy1oFNBb2XYjVHueXkPaAChwfMqh42f3BnoT/Q994ewrh1KH
cQ2hC9AAU7cD2EMtmRlO8Cep25lfa3jjyIhqw2EPxmA/ShkXgRGv32jGZe95hMHEZFrTQ7roHz6r
YbJxHp6POuBCAzEwdYqCkeFqLyFENqiBMdMDFzeQBt3w73Dvk1oLX3QaUR4v/R2Xcqc9HdbxcNuf
Y0KUpjkETvMxVGDBGk071y0qEG1emXWMo1sfKnq0Ns7byv7X69mymO6w+lFHae6/JFMYduuSm6Ih
99UXuCzK7Sp6P41hTTjYjg/+qhiVlaEF2n+ujbfG1v/+Zj1I0JnTkQv7H9eOFxoDo5O/G3+zAuOg
zwBLse7fIZ8qNOkWUAirmv34+nkyeX5EzIvFqgden/mGKIiRbv9+TGtnAhQRLgGii04fmnzGIUWX
zYoECL+IJbZsrMhZfHVpLCsc8+LbfvUGyD4dgJsBobT5KZVVJ5DoqlToFuSB9vnr22cyekI5nz1L
f+0FC65nM0Zt1zoQrF7f6II1cSis+x3fx1GyEX3qIm9N7UtSdsKZt3AUQ4gk84L4rX+zbQZZFnUa
hY4WDqEZ7kqiSs1Vpv00whXihgP4LIvcnjmZAtAwXpVYlyxm+s36kCLyKz+Y7IdK8WiM1EF6+cT/
x1t5xIPwDpspat8Vl8kQQb1p31eAskeziGQGGO3Au9BQOluj31IH7vjvMTovzVf+DtLFsFLKIeQ3
6vjp8Dax0deOH7fWPAqOPkBTSa1YaMnIRvbCVR57PNNe+0vgaYKTIbiS/vlXilWM1JpuLH42wbz+
JWZnTwvZAxWu9i6di6kk8SyRetJSvye4IXAEjPB7/hg6aqoqQs2QPGPK98qVfS5TepqmrztyDbAt
5gVIM9eHdJqqki/PM19t/s0ais0AJMprBqokQ+zYbM6jpgzKvurrpIwhw4uYU3V2y3ZYx1+j/mTy
C1ZJv+Tj3U3Fo2Zbtgzq5QmoR2jY+yvgTS5eFFIeE6LSkFx5+C+12fj5gO1cjlUg5tj2SF2Y5xNm
Xs5Ehmo75fso4Hs7nKhbe4PFPEH8ZLS5+pMaC9C1k1r4ILXnZXmeiNnkVk16HL8MMncbhSSh19ws
PvWB/oZbGiJSyodI5+t+ddIgbHZ9JixGuW/bBJmWxXG82D/slvg45e8n3PJOAJPS1JZB17vYDFaB
GX88Uc+rtPuRlTURbKUsmDkfmANawlsHBmUMGzgVewYHL0W30C7xbznOU/tvGNjay0hOBLG9WCwe
mP6fouybpT+KrrO6wCrmq8bL7SfNHctYeV/U/ikRYJmJN96ZJY4nrdhBf+BJm/dvTK0bw1yWJeu3
7UvDcepIkCFtqXxQVIeAcXXvTaQCJqAfX+QPIxxpBQaOKzNOgpwMBuH/VkRJZwK2Xq7QAK5z95r4
QugpnwXiPVTqDrBHqVEQbGrNS9nGFmNWglOaTWDynOhnxvvt6TojzPk3w42WlERfUKasfJfqOow3
UP3aNFoZ3yyF5IqEZCWUZacJsYIhVAzV4pN/5oSUBOFAkbtt3zG4ewcA77R7AYCBj/UUBjUUNUc1
Jg4i+p5uRhH8xV9dcXL/f1mEupRvSpg3qHFEJAtuMCj+JLh9Jkd7WlGVfVm/nuGFzVbTXCKPuYTi
N0s2wjPmAlB8prnQ1KHe92ofSFFds8DChd4rVSfJiQievtnliqLojab8iH5S3EGl75MFT9p6rt3T
gR3oDsALxN3pdRe6GzDYna7u4/krXp4sznYXloSv6E7Y49Bw2hT7CNpZtvJvUds1/nxZa/oCanxO
ipdknMKn/+bgNnKK5lqFzC6kIBgJ2NZZ32uW2QNauIVqlarzPaUEyZ+lksZ2nUoGEHXYvpNJKu7H
I67XvTgxh7AMaIjd2mvW76+pKSE72XqsxFxhjB7vYMn3/wY3dmAsq7pzLbJECUqxn2enQAKR0pON
OiqONLwPLch/+tKwjQ4SkSjcQP4NWkKx1UcT8em5HPQoqplCf7JsvT5dquazqfw2silZ7iGE0anf
ngl7sxOvwvBaJBdQHw0j4PGmAbeMkjo18uUJiq0i9Bi3Julc93JmeXQFvQSudFcY9fxWUn26Z7F8
m8+Xacbhnbx3WGguJme2cun0vdsulwUz1zsGNQmgGvvW2VOIp65yxN+aZM6w4Es0biK/EVbaD/GQ
wkWV/EQSfecLM3dP4jhzG+IBSXamLbHjXuU3I34vRjQ8a4R+wSj9aDFKVNvj7q5mHfduRTJQA+Bk
LUFFRRxFfFXPcvb8jcTbvsrdsy9xYk2o+RRnGJvCYvXa4HhXj7g2u5U6TjTnSFXDCFuzVLj1waV0
NB9UrRiCKJjSo+VGzqubKyKgR5/7FbII9UdSRzrHtggTRcWZeIni8addvRYRxSx3d9th3PwyQtzA
5zH95QilIWjGNnbnSVQxd9rOZvqtsvRaafK7Xv5Ym29tXpyKaYWn0dujcmcPSYpRxZLuv8TkDWrh
PDF/4OdGGT1Za9lOC/RXbYnpA3ynHr6FDsDO0il7pQ2McFThoQobpCZcuG3DfOChrewUxUPmiJxq
qVTIfXhSdlNCKsuTmHl/aQMKgCxuPRsm6Yjjes2rOHlMMUVWtxV9AVcozPGqrLb7b59opDFxbE4M
894TK8NqYKpV1L+iz60n4JN78/WiBrDSJD3UYhpJwONN+hNzgZPEc3efbgNxQqYLh3Pzc8Q6TLeQ
rPBpJ5fv0O7DdK+pv6yuR7I/ki2KBNsaSEf06MrMNOb1F2p/NOJSGen3B+uRiLnfDllYoF1Ac0qm
WuCA9/1V1DCyiFr/l0DpEgEwfiExYOo7LyahUJX7zjVr3fW7Pn3lUqsWoQte7glUWcBbBuXSUcvL
OzDq3uz6Mx0+pvXp00nnonIxIxnChKhHou41RfeDowuSgZIT4c8WSPhCb4J/f2r2WOcsU4XKjpoF
Q5495ZCqDjUB9Yw0oVADkCrmC8PCkymsfUeQu5OUXWMxg27Ikt9pexTMtWhKjddXFMJfCXwWEsVh
DEJGPmd2ctXjpIQdt5JQ4VWa/zNN+pjUQ3UkGMoe/lHYPm61QSQpiEtGYuOSkJzKuIgPpRTZU80w
sVPocqTPc6VFhi63wOCJYtFAiU5ZnV02PBkK5PGaDZtpKcjH7eGdANiOfz+MsFDJ+wTJbHnIlQw4
54e+8YwR6IZkjDTVmNM9qtUGcP2b6Y59KeJSDjxeMWLkaNjZPjy7vgyc6RHA8Z/lppTSlSPZufIB
oVr8DHYPleRQm/MOGAeUBs5AC6F0rSfBaodYx5Bamq9QR0LDOJ3G/7YAjX2tAj/FCEUz+XtvDAuO
yXbMYvhbCvaH2IBsdueM2+cyVMfeVfHZ853MohCOylMds+rGNsxMRmbyMPcTbQE2bYYMnmHUXbDQ
ZCVDoimMK0TWfk0otOA/oN6PVi7XhC+VH1+QB+O8tHjbMIH/G22tAFeWz401lrgMJlIn0hvsA6M5
SIYP13GchNWvEcDh2alrJQzap0zQvI6gcPYOj4E9p2Ua5+xaHm3jp7AcECidSmDd7crrOSlzsB3a
9I8bh+Z0lqVgwJR2F0qX2XKkeJj1v20oBbOmaZ61a+kSksCIQdjtAsRE2auLggl1hCcToOVvc2pu
JKCgrj9+QuRr6DEercySV831i2THHRLBrZ7B2qzk3/OKACR1s8Ro2gLu7iMEyNT44nUndy2s4gCn
qSQWP6hpk+c9g9mEdMVXu0Zxt0nLKtGh2iuZibAL0fZXWKShIUpP94fhZY3+pY6xnRAKvHzOK4xG
nqpxJwO9ocro45H7ZsVxVtad90OmrPzSa2+IUrBu6Xx+Hv6RxhmwUn+tBZQ7lKfVlVNlVRaZPY9v
m/PeN0WGCo/wjHz8oOMxCs2Nd6CsYjWjUVffNlC6qX3VetYX4lZ0fvp8b9ZZVcN5Bqov3ISRJxc/
TmXLk0KAkvD0c8b9S2B/+m/+0mP1IwrSXBkQ1n7vIunR5se+hsprhiptf1yJtqnU1qjaW6oh6W/6
pO6X56GTFX7bGbIXfCuCVy+dASN6za/EH/BCn+6PN1RcipT1vjbVr9l2VbCfuO2ejR3mRIzitLJI
BT7FZfy/CBOwYGxvD7DSqEJ12LJ6KQdrSu+m0ULdOkoXYljhBaweMEXsGgOco3/UAK9P8fip3RcP
0HEpPXYUgCdjlsIZlGsZOoW8rzcMZzBTrDy/SXZke9zPdib2XS4TNtRKPDmCwGk4QS1yO3DSGyR+
/H4nbm/PVwmcdydTtJGPgyzb2kfeBJSbW2Y9XnmUA7q62PwIflAwdWf7rWQPG0hPNfFDNBZsEEkB
XdG230gHfr/tJ7OZUbH1n1wuzQCAQNoy3Li7gEzumG1eVNtK84k3xuBkG552jvjMEQabhJm4HIlu
+SiMGuza0mgnkIzZEMeQT+voHqoVQushOZLQgwxNCaj3k9pdblOvLMuWR/WeSGp2P/PPwoLi5h9E
wjQbzVYlZ4N9bGCQQqfpgpuBxths008hxBjlAQ9XplRicyu4NYLxQABZWv/2qA0xJfYtf0JNtfZ+
u+iVVF0JMhzKurq1MKYX4tmR031fxf2Bb0inkDibyOVr4gKf9cgFGNnA9NpczvL+BQZDNFxOTh3b
JotufFYzyhOGAzfwvgdapYANJ/ZB6SOgbwkvMKQiCM87+HNKASWdv/GbPP6cZc81NhFG3kcWZLyW
LAZP1YzCxJBjC19i3ZYKJmxMS+tzfMcnMGUaRTYF8o3y1InfgLXzDQeKC0ZfuQjQ+T/yQcinB9MQ
kaZuUqlr789SK96iboqfTdJRm/vFRw8bCYzTXdfOH+7rc72kcV7Pxe0dnQGVZjxn3yv2LXpacs2X
u73bkk3pcFNAXsmVO9QWQzuC1HlqsJXe6GuOJVgSE+AdV1VZQJ1RdUtF9jIM2A4BCaJWU7gIXRKw
yAhWgsK3xfRKWvarj66PdW363i871DKjr2ThV3msyRN0RC8Y7Y9O97E709MAc8wrqGdGBmjzR3zF
Z9Ahwjh4vcLiEgtRXoot52ehrlgHwC8AtubFw5ukhqhaDR+vOcUnBAMR4KJeSmC+WA59YcDWGDNV
PRmXWeOJnRh5f4fiNTpvD3Uvgu6+fq8P4N44+ycRBHnb512ird8LdQ2iyDyKxqJkMkc/0RVGZd6d
BEohJSahnfYSC7gbnDVX4MFPzE5fsZa+dS5CPCWO4eYLV+7IX+ZVqdorFbzPT2Hyp8VBhrw3jKA+
WjjgndHMdAFVpydii3EFrx3BTI+5Ux41OPvGCGaZdTfrxQh/ISsm/Ot2NHYLQUR/lyBxkKHi4pBR
1IWNl8LnH4CjDaJa6ugiGMs6L8NQtG/5lAc5o9OOk/Q+eUQBwBKVkyiJl13RMNZSQXRbT2INSJRr
FOBxYeyhJoHw97beOXrvY/0OCgkij3iOvlugZvkQ3YMVCL5RMBT1tagpvI3SmkRWSN9seEWe4dz3
8261rvdEFb4MzzmazwhBze2hsw4dNLKQJsyiZfmtfSuYLRWqITWtMTpO7uo7cstYW1farh7Xx1iC
/MwO3fxQ1nfzEcpldtWq+1GcYk/XI2qz5mrKwfJplRuxx5foKyfCRj4eRs6izbbies9ToOPSRRFS
HdS1huKjvQ693ExlAs6QJKcTp1yLmE6ua1BfcGLUsM4g5tnav94GGJXCT5MtY7dfU13z1vft68Y9
mhv9PbiXbStLgCd50n630HhojbesiWjFPwv1NTuVy27En9mXkbSD7NZXIRtsBPxValCEt1oQXT5D
KbowCc0jvvKVAzeN019PBkjsaF71M4Rmk5gFjMrbexNOVIdCsQEPOtt1KpdsfH5jNlkIoNPt4Bie
ENIw0Q0sohoG9KyQBK0B8a8nLy2sALZoVeBnQyTdNr1JuVewbyBeI+CwNcykD05i125WD422yzAG
6LIECPCECWK6mQHjsVJk+yMhCJq4a8Z35SA7Ol5Z4yhL9NYv00OaioTZfEEjK1XWFtT05whm6701
IaDgz9exWfbSYsgGUKxBAjNQPiQd1MC4zsXQdwgJhi5zMBsKe8AyqFouO1U9t8Lit8Q8WP67VgjW
2dwRsptPFxsmozl26H9CUHKhktxYrcR3E94G7ayKQ+OTtk1FEaYZRxfZcygy4s/OrDXZUulomNbi
+ETfYgMGRucBzHNJXwtB6IKjbbYrVvzelQtG4PgHsDqDrUqc3QLPC3hhYPB7XJncXv9a1U3bjoeE
9+1/fLYYI+8/pV+IkReh03CAz471BZI5yvGTXg4I/I7Sy/k37JXNTXq8EB5MdmjEyXgRGvNJakFq
OKuBiAcMI1UOsl2C0FZPqwpznn283U9RA1UnSXo77uuw93yB14j/VK7s0omvVVrycrm6+70B+DM9
nykSdBDszUYE+1ozB7eAYU3x/uo6IzmnlTHHtExMGbNszBILG2KX88OyYVPFjn84HNk2vwGqmyBH
Nq3ouPFneb+fPqGxVPGcB9NHmnPTH4LV7XnCNQGsWollTtP1zgdCGAw6Sb15Aldlb+gJLtC42ZZ/
NF/bEmosga/C9QzNbiNbu44avhHLEFkpPPtNjQmWLwqSdYZD94bew4hrKxW85qCRiC01knYyfK5+
y+hfM/yjbJQH2GBuA7PVUiPVxb/RJrpGR2m+PQYCEl57NVGWwIIiEvKKb+g8rDF4wJEo0I2dO/rn
vKpxYo3tEdJHL2Pkh4aCofT+zTIuQfnI7+z2BXY6lPQI4M10K+QWbdydu/6pcBA6tn056ceWKOv1
ZuQaVzlR9d+0ivWmCdHVydzppSQgMvVLAw9Mt0BrzGnwrNDwMjMbqo0WQgV8U4KbmKvOdhiLn5GB
quMXhz+r5GCW7sBQfPltgHaNfeSoH3FjbM3TnylOYuFbO7nmRAQPKyl3NsTtjHzrxms/u/+lBAJz
+chUHdAPzjItQizjpRkDtoqn3bbMuPq53G9L8TSxXgtPZp6W2n2WR/h+5hiBzZRSSh7dE7fJ7IIt
vGByqOssgqkDmkJHIwlTyxloDvO9NzzgDRRXh1dDHGy/UmE8T1ROsRd8mIIpsfqGRIEpbFXjRPE2
zlTIkHasBAKaJRKr8Z/oNPHuswflR3m82aYoZUmmjbV3a6qLm1FeIaRmS3ByWtmznRQq9jzt7uKL
62gGnlzYUjZCcoeE/Epoehr/ERXC7TBt4hDWS1CmDToE06Z5pE5QayL+c7ngoKO4tiZNh8CiqUwR
WnG335u4b5EA3wLPrsclY5vTSiBEvieGPff/NWU3zZuH4hsEYCIJxABdm6nypin5bln687nZecQK
+I+Kc09VVtVUGjO4naI4OIrJzjqvqTfLrzv5n9fjma6MVvDwjRp1ijwdUijZbzpCqOdoZ2jvzDtA
IK8ZKjImZk6hG7X60TsAy+Cw09pg9y36nLEQjuhEl7UdYzYagq0k63tN/+VdN9rU9RWutUYcVbSH
yepuBUJTlNgoLQtZmIw14zGSMZ7RKKqp2u/ny7BeEgGYBYudPmc8uEIKwSOmswYBjar7202eqT3/
ug2FYRPluEMUpWvU6k5g4B8EBgGGGQ+qvNq9vD+ukyBEhgmrAxolcd++J+iKd10A1BX4m/RLcJo+
Cj9yIwdWYtTTp0zwBvYLW+UNisNHxT3J9OFu+88tn/Pew8qdAqa8fE5v+0eoUfJptKSXWaaoD5FC
jObgvy3lyFpUQqnfm5xaaNx5a878Y5/znXyWsBQLGfbZ7knqULOeaprysr92ysIPlQjYVgt5/WUx
gyGXECtDEYb2jDljn7OVAwvW/xYRnSsUK3Pbr0K0RmURzsPmYmXcHZ8Nc8bChVgV5fdnVDUi1F50
0ua2r0hpmsdUnps4JZfMFgtZqOfC/1H9Ncde0rw2bhErk3F+s/b36JxHamWeNksFC3yMPbm2G7rL
9EtqPttqV8SCrQDC9n0ZyC66aM+LFO2k5at/XORrWml7gO0AY4RTceSMrzG7b6aaVXMUJWhFMbhB
1hoMIkz11jOBqFOpekJZMv1HxzkRryhxcrSRrjgfiIuP4Um6aPDLkEuiI9HtF9yYrlddtIK6oXkX
WyorFuolyvFsEwNs47jx3iAoSJB4a8hZDjqrGGQ4Q6/ngTKWHoRzvrYw2iAK5YPbYg00JYvdvZpw
hC6FtnLr7/fQCKKE8/8TVy87O6cLLQXS4843/+gwdQ5Va38k0PY8VHtbyRcm33m7uTYHfzvr9V7K
nWPvgUcY2LRIsNka2BfzBA9u+++7edIb5jT9OjSOtkdtK0s35RpXMV+jgrFMRtH/Kps2q1ccefq3
ylua9HjRcC16foiY3dtphWZbNUpdRI9HGS7p9+PLxJwcQq+Tjuxkcv2YMtnm2V5azb3JiAg/gEtJ
D/scCkAfnJOQ4A78iy8dFZVX1S92E5+2LPumQ3/89ormXKyWtExYFVcskmYCVh1EnPalRBplHwzB
oOR+1QRVrWjh03P+DcgnbqgnDrieKkcMdM5PYoxrQrx3RdHQWCpexro9zHWvI+6s6NXcJCfwWnfQ
iiv1WhEXAkH1BnS9hbG7fR6jo/MwNbuxbGzLw200qV0ByvTpxJ2eZS4GDT8hwBQDOMTeExHl4m39
lphLl3Pq8qx+VSbqTCT1sGLhPdzKBD5Rwx9cfUVlSgu5YNYmGfkuLLhA0V3VdZYoX3sdGyatJ+eH
tuAxQU2DxUhfCJlofV8XrSHIOkBAnbwlfkC1AhovJDDMh+izpNDVXWhBJNESdhye6JNqhqc98Bs9
stk1Ay+T9hLoxNu7Dr3flyJXLYcd9pdEZHYmF+MBgAuFEwRxnIL9hvt+e+YHmPW8/6+rxiIwxBaw
iI4SG4eT6MsR9yNe5D4M06d7LJW7Ofx0Ug8JinaLg/poXJdSK5d427QwDw21hBWG1JKTZL0dGjVe
l/mRCZ7wbvMyfkJjETWjt7I8VYLm7SwkuSoX3YGXlw3owbKh2AJFIVbX+TxYi8CdVzHGDII0gvb7
HSLmLFV9nUI2jOSU4wwg90Qp08dC6o0K1D1yLp8WktO6WorP1KhWCXxjI6JCg09HLKe7pB6orPf1
7jy0smd92x9Qk3oIElRegO5N2wAQsRMyeLd41Nhf6QAwZPNFPaH99j0LNSAapUPqjiy3yHuhL9iP
4BeRRiRaqZKiIfQInCvTJAgDp110rwSRTBi5StlxSH9Yo0luQe9sOUOUdAvdJiRnxVrBik9ywkx8
uhopyK6xfyeRyN2JQoRdjisdH4rEq8Ji1K6fi5x+Ah6fsauYayD59D7TC48r50G092tybngUSYWN
SWk1L8qBauEA9AbF1yxEBjjSr8wzeeiHs178p4IDMtXFnVGa/OSFpbimcOWp365dCQ74YgVPyJuO
pIAgeS/1+/52qQfAa/1/SSRBR0C7vna8qY19N6BUEGvYgFRX4lpy3M0LU6OQfUi90buUrTQtXIVz
jQhJ0E0a9qDK7bPKpfmPvmdWPW1q3/YI9LjALjnH6cZMqPpmoTlDZCZZP7i0ThzQf1Aehp9U3t9z
4UkFKDfaRjbRnJdMtEAossW2x0vWTqn6OOzYbtINg0wQuehNS8vPq4z9Zwvq62i4PamIgbJcgQys
AFr3zzdg8kMFbIwDK7zE+lOnOvUjUfywQnR8X7lF6Roz8RcIzJg84EFAZDC2ggUAK8xCPY3mLkGC
AQOI47oR/YwTrIXbfSAXDlZndrd7/NI1npYCMrPq5EtpigN1dRqjHkGhAxjqAdeHOEU+bCJeIfW7
PQmNxA9cfnSADDUXMa9wjf3l4s4BdRhFOcY6tUadAy9+BBnuYolrkfoF0hXkYPr2Xv0ExjK/Zjmu
86wwYQcFOO6QwH+PUn2s6xZcsNcvZAShYe+rdrPTEKZ/esar6Xt9401x4vVFk/i+uY0U6fWLc8kc
sS1nlIV3bQE2BW2ZZ0yvJ7u35a23DJKPJCpL15pZf11jtVUHBcJ8ucYaeyR4Gs8sbk3P4x2xT6BJ
zUgpffV3pA0bU41vMB6i6braGWXzdGH80IJbnn28JieaVPdycpyyv7FRcnX+6tvV2UeQZ3O282W9
UU2ypE4sVqcZVpHV9RZ+gWOUoR7m1p+lhBs6bnDS8FsNca+yNDsE/Mc9hq6Jq4f9mOKhK4R3dHTN
cnr6D3BSmLoSdHzoM52smci30S20RDyDfR+c0HswI6XIN033JduSiC0W+Ukx2liRD4HYyu7GQOZ/
JPkhlQrJ8/xWOjN6X/Zepe9i/5AVBH8hSDfHAOm2YXT98Btr6HAiwKuiPp0nqCbujRr7Tm6I1yuJ
M/kGKqbxF2a1cPNIwqFo86fCzfQeIcJOK08iredGYlih3PP2uVwpZDwNunpCS7Vf0PHhUTOqp6Xn
saYmfAJBEM6LjVQf6KTwQBifgLzKj8gjEvktTcgFXVXBXrbd7o7eq5a7VLj4g/9oDyXZxFuY4TTK
Vd4h9SJJGUOQweae4tu19OzbquhJrHfoj5hiKh1zRvSbqkACB3BrSkfT268K479ZFzH66zyb9xzY
IPodo0O7ShYQcIvALPc+5R7lZAUqYUfOTaJcJqgI52hyLI1u0DORpcIetauaCV38297H1V+5EcHi
7dyaasG2V0fNn3oUjUAjf2hOvv/MSLtZEjMl/vZO8OqpzyS6BJWhot6cq5oPfbpsQfKrLIHr7voW
2MOuesGtvAeWuy8Hj20AvYv8gKNHLfCa3C4mrGdVpiv07B85HL6bfGFZsvnI+IWOqT/77pWNhK0E
k12j0M+A/G3vAj9NqKWopy4Kst0eYTgHvCSBfremuHWLaZeP7NnvdywPt1+7fVMf6uRpGVn5pq36
EN9XomdcSFrrmidAcEVcn310l7j15krIw2KkMwaBpehGgiwd8b4meaTg6VWGg8ddoVWy3pv2tUoY
cFumZ7xfaUyJ9WOPpN4HEY8UJ1OcGwCncJmoXGkmT77v8a6mCLfvw4ZYiZYIobkF3ZASyWovOI8A
28OroXYmHuq0HYbcaLPsxrx9gSqi9dPLz3L/HA9QLywR9WzUvJx+2gw8OYA5gJ1z0diQeUy9RPJk
tXBU8TScOIggNIO8z8rwFP+gTMxxBZoH/iaVYwpxVzVoeHllzfXWTzosTxEhomUYaVS5T9EY4Cv3
IOK0/ie1bD5blwDPVAgujO9EyIkpmBJ93hYSTaILyIy3JLE0bzr0JZKouKj+JE0NN/LZEVKvBduW
UhG2IGaq4lQs2nl6ni1+jUCAl6RmPv+Vl/6esADHmrbaSykIeenldVS215pmpVkPo1aLP/WoBPfH
V4NtUIwOArDq6QAPeB0AXi3rfO+MBMzakRHghYoJsgW2KoPWiECej7tJjTkYks0OnfE8qBJmINOc
XEJb5SlqXC8hv9R0tOY3TgJGn9GpioL0+OOxBauy6a0/oDFHLPznKED8wH0LNoPNC1vQWBk5EZG0
WSlakCMeAr+mY6+yvI7XX7uAXPQx6pOm0pXoRZnXUAY8lYUCXyq6vT0cXeKK6w5V168Nq2ttGrG8
L7V2go7V9fMGK9ZEKn02E1kAle7V3HknGiY25LpzMFv0dekfmJ/R91c+iiX0bLPSLkupiguCSL+k
pDHSzts5NTEwEQNgdRBDBEzX12jsPR+IBlgmUysx5rb1kkxJSejmTxa0bhBh0FGkE4kwicDRMSj3
rM25OGIVTM4iouCWHswp6vvxcHmTIMuZi8y8RMaP+SVOYB1kOu0Bg4rGLlFr3eCFdAqukoFeZJH/
jyFpqca+NZr27k6oVW+nF8k0h6Ihs2CO6xm3Fw2VuI/yBMeTsH92KNwgwP9Q40do8+2jnpSi51U2
sJaFArF/mxmsMZcxQsyE1dFKwnd72sAH6zOtSY3Amnh1ZQlD35q/W16xiGTk88d9s/x2cRCZuc1/
X6kXMZ6tyJSGcA5g1oxp6YbjfYWfDlmjmEF7h3YRJ6BDzlF4t/q0XyWWgxC0Yslqxh4UfuBISRaY
0X3oRixAlM/trdWFkNYIF1Gf7mYc1MtwNQUPoO42joavNzN2JzDag4dKgWK4ABmYO/s4OVVl1/7H
RKw6GZ9pN/iOl3JBwoHiODro+6MVVRn/jX2reXrrMjeJMKn4c66vE62GItMSOG6R+DhYUuf5O/e8
EfVtLFrcsdXDqEDCYd6p1pnEOsR57kJ14R2jxWQw8yhbhWzVO0MV88ttwcBACoFj5dfQdVY3irUX
W4+awJVwhqtGGQgasQ522XpLl9zWxFesaGgsNeJS8GnwV00ZbKRx7P5M0vhPJ/AQM/1Mg02gp6ov
blz2QiK0jKPnst4yb/QzL8oiEuhE3kCbqVto/QeZldIPX2aQuLEXNDXCHCgN0IHTeXGmQAjBzo3j
zj3fcCyQ+gEK0b5T2wvpgaB+b0HnP/XOGzMEkJcYm3vdgupEeKQAgPMo311p/SJHP8GN3pxJ51Na
YwJSXnhSFoEfRekalmLsYRFYsCRIWMwv3GrLQQRRIZBsPpSFiMV92QIqqca+vzUbwR4JryghF0Tt
Ol+RMCHway2a4GIMzcpepYgZJfLB2ubNFESgElKHuVN8RR7lTk4HqEHCTy8gYTx186ljtw8vLv31
KG4vnxFyl6s4Bk0cc9fgc3HKfnlX13+8LZSRcAxCvv/7XE0dgveBfTFnNHiqfSKRZXiqxHTCuQy5
ciNXFqBcdr/HBgSXQoIm0BZ5ECyBDakLpLqSO9gyGbvGEdG6RqmdD0gC6c2dWc5G5MeX3zkJEh8G
KXR0vOXVU9rsT7OlRtuN4XVl81BPscFgP4azR5OW0+Zu3Tf6vevgLu75jBjkXZHenuGE/svjHgCT
gB27XQwcP7bjWv8DuimuoNU+Taq5h4qfPPDEkqEZVskDrfJ2XEzwIwSvWMoOkGvew2cS/45CvIPv
8R3hZFUXh6iDxooARQT9aTRyGXpEElc4ODPjv07MfB5Pqx9UWSxClGSgq0YqzyeXhK2W78c2F2bd
zYXvlpVLBCB0CoQFSQ3tj+89ovWwrK9DMSyuwiJ9QNu+2EPKogY2Vqu2rHo1msf9l8Vp7PrQyrFI
MUzSbLtYLH92/PBaafokqDMbCQT1KHmNABJVLTNLrubvWULUEnXqLrrhWRTo8NewECVNauBr6bkY
r3lTdvqHQVIGvlz6/L9ePC8mX1TOlLaIy4wMYAo3L/2Z8EOwN+c48+H8VcRFPyvE5l+j5a0gW4nx
0vN4thOTlSAVdM7Ck6wx+fLNxextMe70RoYzJWSqYxgoMVu4QqHWSvn6rtAfI9PSjVlyZhepGm3j
6n1qhQUFG4OC82D9GtxVsYNI38E7OWdnP6mCeNJZz9Xyk1HZ76cEcZ0Y9G47mTXCLoAEVGKhZ3xq
BxwINfg1EmSXrb/FY7iBeFsHIaGVW4dbwFXXnqzrym++B/IEMk6Nt2VtEL5xZHk45FaWRjcWXnPr
5vYl8W3iQBlbSbxhLWyOZqB//qzSp4zWYUBU10VoHXN6Bw+O93ZgjW5nbfpMV4xhqVObhpylr/ln
4HQOjZhkQVr49CksfY+ZZmTMYDcwfcIAbPUTjmDOEgj5Lge6S4fNY2TejfXFq7HcUCuTcva8YRyh
WVtKDutbuzwh24FwXME3ldDbUleC2IvQ/G4OqI6Z77CTvZ4LtkQrDcKEJ/t7pxFBM88sa2oE9FP+
/BZlWdxALSVBoVX44zNkZ1oGTJtalCl5I8pQD7Ro10S53w5QjWl9WBMWgUwywtfzVa49pdgxbbgo
hgrHWJG21Wuf87WnRJiqiRDNZjtBNDx8oKS9TxfDeVy35KjC7ERUjNFaKFXa6HoggTkgbXzOZkId
zdRHda2T7LFwuB5eDrqOdu0cx9TizT1ZTFl/DlVryE60FWClEDSlvoyQgznN0y4axiH+g/w3DwS4
Tm0osN13YnyCKaMbzQ9OuCVGTEG12LZkSzSpBdyhf6SJZ/Vppwxl3chOmjtdzIvuUa9pDiuuG27Q
lYEZSfSu2Um3zyJK+GtxHZW2BLv5jaNlevPr3gxkEvC5+A4iQ9pr8hgPIX+z9oRVsvzOeWi79BHH
tlXVg2OpI/eto1rmgijSJN2NJhGcZGhC4SkH+FkOCtNx4YomOA0/TGXpcYmlv52hP/vEp0obUIKY
aHtCO2nPH/sb+QsJ3JmEr7sxv/CgXtk/HfcKSePPWXT2TcK8BCqMV00SPXku2dbWe2zilhyxG4Ly
y2k8FL2YRWQ45z1YrSp8wCgDBExgsMV/W76mDj9TjgF6u04RLxpzxfly4wW2naSe+4g/cu1K99wx
9vfiUnt5wuXeQz5/pcllM3bPsFqBJKX85VZxfWjyegsDxQS5SHsrKvNodlNI9zjHy1lvtNEcdqy7
sC6vnSgJh0qa+bLC5u02AtjVtDBSI/HdUEhFY1VzSB4SqopDXcTpzdFqKqirSJojnt5vkrZ0YE4m
hOxRq+GYwFlCs4rcABwHBec0aTP+mA2/KCixV4CLlSLS98aFsDlOene3IT8foDKdVhYuOm4cZjwC
uRdnmwtBAlZLp03sSt7iatDW3I1CuGnMJ3xxmXDTBxwMulCkpcG03z2KfhDk24JCbzLl1limGQMU
ly/K66CKSvBhV2InvqO3U9KYYHCGckKee1+WpHaudyuUMvj7Q7u+h5YB3RjiWOqtE3JOepqYZ0kP
9WbIoLb4CIsVWIrIhYBm8dRRl5YdPSTPkgWkGIY5rOqmz1q1/ke+1OSe+kTNvSvu6WNGdoHJczRI
vk99X4KKUtu/bbi4KEuPSoB7B2N8II6lSaYeaWUCOTOXrCy0r5tX0hjR4T+7OF7mIjiQq6vHjdor
vb/T60XvsI4klaI441cz7hgeNnU+q8Qt8+oolOjs92BsIDzLpsTvLz9snnuxWA04n3cR9g72H9kU
tWFEW97OoOvSxUFHrF3SdNLcFBbXLLC/ROwYeb1cVSBHI/JwnZil8l4f5yboOOPwx47/Iaj+zXjh
+P/3IWsUnlWGrpHRVpKnQGdZ924evNjlTqh+8+webbnc/3HQeSlx3QY2RojSFV+nfkpXRRmfYut3
uvmuwLwXSihcmEbAJcp1f2rafeCp/bQ7pZByEZdZ6nnv1HbrtUgF2UtlGj2+9guTVCaYhKVvN4ON
0dmBJzsdJrUCnPKqBpugr+c7WmdbqvPygqJ7fwh8rdlQ6vQTP081KO30tzi0T7Y7LGNu1z/Xc8Rq
hiU/XavTYWvQST/11FU1E8e5mSleXE6x3dIYttwaqn9SUFgb/u0NHdUYddjE7P9mUscn6npMJkPH
eOmkcu9Z1pYWWyKq/cXFyWRChoNtIiVPKifoMm3uDBLodzt3aUjbIsGgZBluRz9xLUafaX1IJnRu
h3VCdGpDDr5/U5bANJ4gm639e1PUD0zGKjwnCVD7hnlJjxcDlHUewyRRMILX5LlJn23YYB9A+3Wu
jeZlzNphuuDbBzjGkHU+CzlUiJKufb8WRG03W1DtfFfpe+FrImzM108lFFxzkJ87+OC10Fsp/ql/
xqqv5/NTD8ubPPzUXhf6GfOfmSmeFgzJ9Z4cpiFNCStTUqd1T8FzcJZW0043xSq3MOjIsF6+Lf1z
+HHYno2vZH/BmjJTKuFo5U7REDjHPaiUMBc2tioU6thzUuvmFTH/ve5NUa/5JapwCsjjh4rekyzU
ph1xsVcRBknj7IVCuZxbjuIJrqCbswM3cXu1DcA1pO2KD8HiBYbHMylUVXSzJvgDGHKC1puzSaGL
QhW28QTTqWKooF6MfP8U3+FIVYMQFCUkDHRDe08KRHqw49p0PMgrXc36JSKv8bEpZzeAFMPsmzbB
TyCl1yCDGcoRCzmVk3jy1QDNc/FdEQuS4F3fPadzUCRekHDJeExA9ocNVZ24XHnKdNUhSCskdZYt
atU+/K6WEaCmhWs5hemg9Kscq8YipZZxPUD1lliEKO0HSUY72tKrjlGFsHGV9NfQVnMXFtj7jV2b
0WxZIOIY7DibxB6ZEUOuzqxo1zGEiuruTmg/Oj43PE+ZO5jMrDM75YteWjnqB/JnP69ULbm/Q1z0
uZE/8KWOzIIwHQ0up3WTXb19sB4YaCl35y2eHOrLV1jiuVL8XURdbxGXLIlCLnU7H5rYZcRK4wvW
Q2JDoBJ9Af1Urzq4G3gOvJZjhZhOCMI3/MW8M75Xmnw5gV5icXlNgOqPWI8HMEV869HqG3RlRclf
ZaQqTdS15lWwa5sSDAIYbPK28dvxmxODgH5p22vpL5knjuutFQW/3PULkGO8frQwZ1Cou2QK3IIY
hC1ZNTOAxGvxrZTMGkdH/LDoZ3dqthHuQLUzk+x9qbmkXlX2sNZEK//BDRv+OQ94S99OWj9Jwalw
TXrZ/bp6Fn24ya70ZtvENxlxGjm4H3uFb2JLZ+C3edEdGzIJIDecVioAQBtc/AjF5CDODpdpqLHm
iQryZfWN7sbJnUBNCQhFeugB9G3Z9w51Hlz0w0tZgO3EX4yvK1zeztm6KRFKcaXIADglaGOO356a
iA7SaE6YV3rLGkgfSY8br6Qy26EMiu3ZpVhE1q7vb5MEYSxVDMc1wMFz9g35c+WO6mWEADTmo+ry
mBETDBMByYDnadqtJh1E4ebFEeC1QhnkO13QlUWxaqstFmE7kMOhF+xkn5SKoqs96XJ1C9jOymBH
ZvY4v8xctAR0dGwhzeCprw4EBbVvGtpxsxJBjz2Iv1QXsH/iAe/GxoLxt+SOVaqK1dyyUd514Lnh
7I+bCQ81k5pnNsnEHDiUq7FWkYn2B4mIbaYUZx5zwJJ0Pj/08sAlnNmN/NYV6Tq3HjBrDYKx/4f8
YOwLHlzKit37/zxKlGnMF9CDlatWMintXOmNWLJI+6wzsLelNrDPR7W0yYvQuFNCWSulrFtOKFcm
OgOHbTAOkPm3fLYLaDbYHLDxrg9BIjvCdXvOPr089v9nCOkrt4dsR5WvaqzWJZSFwlngMyUdrOQf
XeZymBKRsNEL/9lGk7TCBKRCOlEWBmaB1E4f58gSCroF5t3H96CYlHQ7RJMXcdYJ7VU0qaTR3JQz
KQHG4yFWM8RWvdsvoDN8kWmztMPXUSz50j4olN0tlidFxhUXtcdbFHrmtrmovjzyK9Yr68Oz6yJ5
3I2lLpNisSzFvikkZy09Wff3qdUGL+c1nr/wEK6CXBw0fejPDhGL19td62s4SE+epvEF5A6j3VSy
xFZczMvrY0YDURcg2NGSKFj8H0WCZAciNuqHvU41NLzwvZRYd60Tm5vh7Ikpoj97GoLfrJF8J2Ly
suwnMPg9tPp2QBG2uI6lUHkXP8ELxoLDdTgDniQfEpLo2egHuAVQMf2ivd3Bfh0qCrEXVYLvoPTh
jkNyvDlIeJLD1Em3LnOdo6BnmNOikKLR/TRkzkulypl6OFud244TCm3+RCwAOFbuqX10beGD/kQG
R+cmTOKj9B7kGIn9zh756f9XvGZYBKbknrd08fe2jKbfyERr0PCizhqTBEsSQAr5Y2PfL1B59t3o
ltisolLhtpXkI8HPtfAeLyIecLZO20GUtPv8f2lu/Ud3VMfYBWWnwnbxC5pPJVqQvMQCwwTzAKXv
uGat/GSQhlTS3ejC8qY8FZ6C26N9iNs9UbVu5YPW5XW7SlQ4M9Zu2gnR07KiS52d/WqjA0Vo5X3H
BuuIDhNg3OGzUAzMJshYswjidTIUoQhv+YI5KBzXE3HSojfYz/mB8UY8UlLj8EAd+3rVcPXHtD7h
6iMcDPf1agM5JcevU+NAImy0xJ7b26QoB3I9rPHt9vx/OL9Am9U0kg4NqQRQwjDYTLjYL1cfHLHx
z5iA+W+IzsUxNRP1Q8gAYAJRjcvpkdEP+Jd4p9mhcrQ6fKw/1nca6Gr2AI2CQKf4dpGz0Dwuzic+
ppwpmAXPwo9dWodnYHhJYFx8qHWaXPp/do2Z7fb8KeOZHSPLsiHZA0cS5db2mSuQN7olUoVNQRah
hahlpVzYeto6oloIaB9Z/ZzQJJhAyMyfTck2A1YPAtTqhmL3r90dQlU0DOvmtCteY7Skadt6XZZA
8ebhEwDEJ2tOhKL81FDbrRmQR57heTUo+LnOkS9RXsZK3ya/J3kLzYlk2vPsQ7wyt5WHSuG9ktCi
8JrnVqefx9BrWX2AR1kda+/hEYWmVvuMwOO0O9L//iCuAYl+JchD310V5X7Vkl/wkhMZ3jslfalq
QMbkXWy8gJ1IL0e+5rElA6L/DwZkh+/8j/JDel/l5f9m7jq8JrEOxZWIZ8nkfSv1emIsLr70y6Ma
N+sDzAXbQBYlda5yZZoWSQKZITy4wvrIPVqm5zHVjZS3eTl4t0COrloa+LREpLZqhkokjazpGW7H
DBDfb9yzS7qXwPRHC/bwRSVknw/Q6UNyfFJjHqKcVII1qMXrVqFEHCT0F8kSvB5CUSTdrwbq5ZAI
qJytD9zGCvZVCP/RZK4FJKKYYRf3vboubm1EEFJcMNLN7sbV5+PJMMoNhHL86Rl1Qx+ESz1qPW1r
/wH+2UX5bbSTu9NYvrTY9ogvVC9eqrFYSZhJ/1hmSdbxARvKYSE7JXgEyUiW9c486WZ/7yA6p7kQ
YXAkvRxztjdaOMaAeVdHDAKZr5BxQqp58cxL2fVnNnSWOA1OX5smaZnvZ4u1eQI+K46djPMK0u32
CaXjXvxqj3hteZtWcLo4DtllO+2CO5RjhcNomzHrQSNzecruRjwvVmk5FeXV6YLqDYo3YNwQCq0Z
/X0h78nC52i0hxY8yQjeRZKv5XZ5XoNRt1I1Laj/+Ocyt7XxfZlzH1gwwow3et53xRO5CWyE6WET
EtxQUvmCv7bN0XaocxBOfKAXYdLvaQwBw5aArJvCNwg6F4EwmiQPhmOLgLy58/o4xGtRFmWBGWr0
+RZxEjFAr3u9D5A0aY95nOtrfTE1sr8ztdbT8tPzke1V2DpyVf2Z38lm/LWB6hYBN9yUPa9rQDPW
zS9ZvQcSRZpqxMIclQ7exieIRrJIC6topTtlSsYNuqt/5S89NaIdVFWmoh7BDX4IbC8QDMhvxOJM
I60aDFUthHVwV7yIC30HBRNefZUHz+nNrucg9JCSne9Q9vnmTELOqtzwm+5afEzVH4Imn5s73wiD
DhJOzofXNTeV11kvQOQznYmzY+sf6sGt0zpEvCSkTDhKtRurFVWqI++QSO1h5BHIFOQ3M7K0MhMi
qdMDZtRXbeAzis+uKgsm4kXYge2UVdyQL6dXe49dvM2nJQfbyD0lIRJoWbooSUd54ysw7g8MGUlg
YHp2GI/pAeTC+Bk+Rpw9UqOKVGQXg8NOumBSJA+2dkN0Ngt6ffFJ/HNSt24ScMcep8CAyb4WcX9g
rzNPn3+OR0UAS4157CnD1kurIoJUctJwNsOshMxiRkmIu95YxF+xjWXjCgUd4xjyQQuIEs03q6YW
aWGBYuuiSDXPRKitMdaVFMCZLranCsqteatBLFa1oJ4SktBK9ylicH4zb8/dbR4iFu+z4QLgwma9
Lw0+QgQnY5w969ytaVCIfbU7xbxi0T+qFTfI+TK1iQKHSpCbSG4bZiisuxMbYXYUj5D+Kv94PflN
QjLwUaQ6rPxMBHWrFIV2MteZH9/qeBe/gLs7VFRrKm60EOchGo1g65omJlVtr3enRCqezhTCXfkg
LrzWbw3aig979Spr5ie0azXLSmkfCcSxft/QBVKGacYCkztaKLYTe55KoVvcjZobMBD31WkPmInl
lj1lFzCF7akcIaT3vmM+5eifvx6O5Z+97F/F+cSPmi3/iQCpkvl103geDzSS880OKAzN0TAIdr3m
3zIrShuMsjvff5B3moq1fTmJtTL44BAPL1NSMA6B/XKTQIQf03XPdtsxyF+6EPadMTG2zYIm0My0
y2vr9TIOLd884SRaK89d7YFdAZs+R2FYVA5jm/gB8hRwshGIkjAM5N5vHoy09wXLQDkU/xuiZwY1
TPtVJ9Dv2mw2Dd+c/DC8yhDK/WI+W4ZecDVE3DzqxVGDVOLDSuQVGqw7IyeJ0DABnBUkPB7ExBqC
WMgLHgRPCLsLzwdweN6SD4WvvlDYSeu2PQS4r/2l5aaXqrQ+Bk9JKPo7dnydL/ULIpEGeh3M/zsl
QcJrholh39e2rDvaAmhxZx16/Zdug3cDu99gFIAaDxw6Kp5gRoJFA8jn7BjdSbNw/NSxlvDkBJan
xhIwbxV47I8AVHGOj7Zl04tIK0ghVyTK+KmF58qH151JrvHkkWl1+OxmA6LisMNG/EDVOCgZoXXn
myn7Q4Z7l3OeARsJSeIIV0TtGsogq05LbX0SPKzQKbfVNpgF69CmrzO59fQKSnNPudCxWnsgZaqh
NQzvx3rEsbssRe8fH5UWEdWCKVnEt8DCJ0+TIplSZey7WKAJJd3tHVpa3C5HBBtHj1HriJeqyXMH
+N3QoYbvzIh91UdJl+5h1uEGvWKZUOXf2lvHf/QbmDiOT3LxvaiViinbAIm/quKFMOfNQAQwcsx/
/0XNGUtsRvRa8Q3+nMQChbXfG8TF/pkBXzGAzmxQyFywsI/bWjuqTGCk/tMPtIv0g2vgxljp9krF
tbm6UtBYdR4mTwgUyElquFwTmicb6GC8MuRyEz0f++wKkFofDSoziv/togq78CJTvpq7n2Y3AHrB
A8YHxtChvsj1aIJzVURwhkrd7Ox/VVlF90NsBH7hcTve8kuAGMW19riei8gyAc98wzLO8LQBQeIi
HC3b1ocAUzhRLQCpwUydRmOd7dh59uEzdSh2uk6RbXHPjRulyaUDpc/5xpDWPk1XJPL///0CDyVH
lXSWNmFnrBMBrxoxv8evGDNwsjEQvmmakkwuCucVRbAvw/04sWas1eB8RgG+SYF1yex6moCt7jcy
aI4K9CaLq8qnHLkT0BUS0lGMBQrmUzwsgzSYe20dgwApTSUE/YN6mRDjL7f251gvUd5N/g/PpcFZ
RNw+R/KMCcSVq6ePtd9UY7sX7Ea1tXkL5HMNZWgCmeuWadi/N7s/da5Fx/uJmGVORyWVxqTnytN5
ckHfOoOHdKns5sa4w+TAAWBBQqZHZDjyE5XrpUKF1+XeZK4dQppPBpI+njC8/0XcjZQ8uKSendhL
uvbC5bhw6DTovrkE3U4yqBGguGX+RtHdfLEsXaZOaNIAV5t0K3LBZT4V5XbcJVPvhl2RTKzqlu21
Ev3eBtdZkVYzWysxbOJGQqorzFF0YwtfNg0gqn6Sc7ug/eQ2Kn8831AKmNYcQqa+en3085xCvP9x
0DIuQ4I273TqwvTUZApd5wVAnWNBpYaalpkMTKFUizgv53qR37dKwc+7xum/iNc1VHGpPPxOAPhW
+xlfILxhsVMlBFGKbWIM5w9ljtzoCQZENQNCuoWAYUSi66gjabi4w7NLjMAh8+JXzfdrAUFrjVSc
cDvva/LnEb9sttkH7s7/bkHQi5CLUT619hjg1kNpdrH+Cht454FGvsrXxg/acaYNrJ0+zjuZ2reX
6v9gbgb8wUQeW284KYmCUSn2Ee/Pl5WxyB6pj/bMtMljblmG2V4l0mD6VrzW7kzABqiOlJiCl4kL
y7VrqU8aDBi9r5CmxEx2jWvXHcA77QBw8BrHoYnQ4kKX7ZO98WO73T7H28vGUsoSnBiptVbZa0sb
+173GZB3N3sF5h3cUWhmMtWi78NsakYxnXHWlFV4iyGVkDSZInQn8e9zPD3L1zQDYrp1ZY0akO1r
HZYMOBRoz0RujrPgaQVNtE0yYWkq6+Y/Ggjwx0xn08q3HEcFec8PWMhOky9QohHbMgd5dI+pEkYk
10W8xQhvJdiXK/6LMquQhP6HJKs6hwnTVZ+Pm/QpGSc974UGeOD8guPef8rS5e3cHLhtQJQOl/4d
3oZJoKP5h3bgnZ+9qgF11wKWI8QZDYLhBIK29yG4D/GyAE0XeFzxzUnHSUSeZ44q1PZbqEC4+fe8
oBL5tk8tEDCU32H2GGkCr0f5d8pfcUu1kx9oEbm0OyTNKPKFphztaL67EgiVM1AQiK72IIQ6C0CN
pr+ZkyrNc2B+ScdJaDY2LHxdjB8SnOfJ6jL3UwfchzRfysJj4qUgGTTCIX/mvvCHOVPp0hn0qXEw
eUkD7EiHcL5qibAb52Zsu3YbLA85Zp1v2345ADgT9krGgInAE7KsPSUma7enIthgP4UiDxr0djHx
zax/YOADcbiTrSeFT6eduDLD/z9+be/pTWvvRCRIPh2NO6X3WLaTADW4zftXbBloxDnzLcqcY0kl
S+hl4Bn+3yfdWXaOgDdQ5zNZvJrPBVHbk46J2iOD7U/a9IWR+gzDxAUGlc4/3frDMW2EjjOUbCVU
aA7HuBBkNjOdUcvo7dtI35ZVX2/Ez+IFfAnEKQ3ZfhT2/XRvuPfFyBzi74kPcxFtttma7U9fbEF5
penIo1QHn0+PlmFE0q4DN6ETAPZVOkcAX5xl3uAH2WTIVBnLnjX/M3WJFqaDKwig/RRGOOdKQinC
ZcUKF0iCoNChM3GyVzup78MeV1ExsZI3skZxvj0jS30GNEJBJ1GC8fHC6wyH5/g61V3uIjiLQ67K
y04Agq3279yAUx4nHoOY2VA1JbHbqgcWIXW+n2qSp7sl4MoDb/laZT2Xo5VPgxjl5hWdp2x1JUQo
k2RQ6ZeFWFHElCAd0QZumEAhTy5YihLzGg6MqeVmd8cJIJ2/hgRUgMwXcbuE4qpQFFMffrB15bF0
mW2L5xsmrgDpEpYtuh9jTHLPODYW+zp75XarUYOx5VAUbsSU0MDGR4EaBnk8mxldqAr+7xpqiHIl
lrc+uIptc7Czp+W/mo6QOjaMOOk16R+rj/o3MZE9/2iHRb7VlgPva1ILfzaPx5d4gPriNDX9U+w4
2OOJ9M/sa8O/6O7Sz3QgdRqMLath0xgU8AD/eXiIVZ0D6ji0h6McMtpXInX11ufz5wkZQJvfCcCj
iSm++HmtpmruVgb6izguQJLIvA6t3RCqEgFuG8rONSNmJeYG79a8M0ccXwSS9AXMz/rc+s7ToLOd
HswuKmxJxXxw4kGvkgr7nARmBsxWkUqPs2s0MTMQ5zKk0NoTOrB6UVYXDS0xLmITeoj7/ccITBf/
X5kJ/CK7RuPdiSyXQqp/PIPUzsiCtsdbIiZB9e1tST9GvAgY4dwyshtZ1a5s+OJSd4eeNlVIfXC4
7BB3NlIyaTD3tSlIT+Knk8j/wX/G1tze1z/wCkt74BLai/AXIpR/2REuJctlgSYhxrOI09LH7+1d
wShMzFLchCrO3zM5lXEx3FuWmO510bFiypF4+/pV8LbHVswpiEo18+s6E5WaZZCQHKr1Da6nWqv2
DBnJ8FJKKWQWBHzkzCWjhvL50ob9uV9ckWjBhi4SdImh9QynS7zkHGhajMJUm171kpybXEbRL5S+
UC7Ho81zc7QhM/JZgfCfiP/umjB4axVVpBPpHqz9Vj0JIofvP53bfVQVMYpzUpIRRMwZSTdfKqOR
rfBO2fc4f/GFDhJRfhD0d2GGTnQg0lku0XPtMiaXDOPbxHHqPJbomOBgtLDaq3031YBTq/SQe+Ed
mhUKlnPobtd8oTzeMD3uTFgrCXHvOuJFgzS3ZcRnL/ro0WmYxWFlIlBwkWxLMn5EtZSLvovOd/ZN
hkTx7Gc1G9vruPm0w494Brbciln17pYiRhg5EIf+iKmERBsy0ZXLUdr2BO770Hc24XCicyKaY6wv
7R02iiK6AhJWAIYioXxurqXgAecVNZswQAFEiBpVp8z8YqjasTkTFyjYruLoNk+LFwl1Xsr/OwPk
rHpMkAbru4VgIYJSec+zZo8SEfpds9Nn5OBx4y5Y9ue0paJkcC7wKiCIQlN9FQe3nKYHqnlvGEaF
mNXLK4nYGjDtOvMyi3IAvDfD9PLusOjS4BKy0lcwVjoYW0XfHXxj7uQ2XCAiAI46Nl6fQ5tbRsVQ
ntYAyqre9pGPHjH51twNw650T+kriLhPZnTkSfTm1AqAWj0FbnfzcH6PodwFkMeEMINntQTTs+b1
nUcYaO/22/Fh1qYIQlRPMb81olOfGdjCJ2UmUmL9PTIBoR3jlVTtliHoUpYvlurpaUgaiu9hA42Y
qCufr4wXGeSOkMPyJFIcZhWUQQp4G0IoIXVXC+3MCxOxh2pmfAcfRqdGmjk/fdKlSctNJNPqy2S5
8EFNgJnSumgr0xmN3MI4YEeWSUtF/f0GzSZHS6aoz4HreH5rrIHA+W/sIVK4KxpYFK5kta4ABvnt
A8XC/bhv9d3Ncu/xUrQTXv0K4kdZsu9lU9bGDheI83pUN4mbnuNmKbTOiIA9xMMbEb2gAIgCnDLc
cBe37OKRf9LTSqFU81gBlqAfGMFlKXMoySGvscK4zltRliSGQecsQq2IbKMHZphvlwcm6gJwPW10
CzfGBzPmojjCjPjqhsRP017WiXvxClvIuit6LfynS5a8WqkZOrbB25RZ5avA8BQq6mQJOtWa0ftU
DQ13UCjETmMb8itElWlVPjt3hzwUcY2HGesItqPxhMWs321QSql8RXTKmj1GylhkOfpfZhwkan3f
z7DQqAILZOs9MnEIHS3TyC0/KmbozddFIT5oe+G6GNkGbm8EnsYGKn1pgsKQ1pyJ2JBqOeyPFg54
b3h9LvX1oWvpn9/eS+i21EyDzbHVkBe7o+qETvASxt7qou2QLHkx8lPMg6jG3+xRCBp85UVsD4LS
D2/7HJDqJ6SC7JFgglVj9nUtEzCj9/iQ5PwUZv4E5TzPRp1xFhpdnzxCmxMZCbxNLsUrrUsbvr1t
nALRkdzhcvlY0gMBYSYkx8/Xho/li5rnrd5c3jAJapaOqV8QuqYsAZ2l5z79GcrbiOMvfcBT7JmU
oIak0GZ7f3XaBSnWSKRM5dM11qPYqwB0AX7KIjogcpAXb27nIgLbNVa3qgaIyYncZ1HjEzNKBrY7
Etr/ytVNLoZ+QiNlIjueYSD7/7qOH8jmcjGlhTWUX/PvbdMw+4g3iJwPgNU7KFu7g/p22PhkSuo3
7WyaZ2wKlygR5GX+wV+RCW2ZUEfs58c0hSUkgzDRrjRovkGgL/Hy01CvUQqQwJg1jlk3k9NoMYkX
JoMeEd0+oZjVggNY1k9EeLYB6QFp/xdKWEQbHSj81TaRInqDN+wE66YhBihsq6xpx9G6HplKEhWl
iJ1dkIJ3OR6cwSQSqAJwx2Sg7hVKXRLijrhdkTPP1kb5CDCNaDh8RGVMt3kJuBihEc9bCO1ZVchk
N696pgwvctddJRkdBclZwQr//dbCeXxuoERbXXy90pSTLDX63oPWPlES5Kk8EgBeV1XyQMfPhmAj
Dlg6xxcBuDwKkT/Zy6EUh53mUuBZtzOE6hfJC/AdqoGPbOZY9uV+/2d8UPa2BLKAs4zGlGzAxfDy
TOp1UIankC/BCCEyA7Wx/Bo/OhBD0Qm4M8WNKnwWkbcFRi+QcBxLj8mrGJR5fj5mYgCnIdo2xBNG
hpxOpJjBxYzUmolIzM1ElL2B8DNFmVTcgCPaBkr44Pk8ZhAuLSJMUSXG1l85aIrCYiiRE0hHoti0
o41syKjGy7BLgON2oZqtBRw7wN8CkRkdyHmMiJyjyLwVM+n4OgPr8dmaXfX+2U4IusAlGOkIo9+H
bI5125V2PMhbPwFwO+ewxBJ7aY/5S/W9L59eRvQuKkj/joHYBVI+E5hUOJZJSztX0Dg1bP8aqldS
1MicUQF4lnS/z3I3Jdp6h9ZWrxW9bmIS1pig4l2p3NTxhMBYF05vRzLSAJuvDECoJdNi3Se4gV35
pGUvKzJYlsSQKspb6QJqVgCS1dhtuCbcSQ6Ikdj3ezsCFT67mlS/EJIk8/zYVNRVuawNqShjglh8
oRycJaGLE/1DZL8pBruoqz4gNffZsWIBX2PffJS6VvFqsb3Pit3TgmLAnMJmRRScVSWy2PlGjLqw
tvxEUmts5jZywlXKskNzH7jIx6yEBdyZa3u4UwXVNxp2TKPungGNNYPouK7sN0OlO8oMDJl/H6j1
xwPFLhFcgWPUstBHvZMHZ5UNDEnJsVL5uR/EJOkI/8B8kLlGLzfQXIXsc2L/1pPL7RHmFuqfYgjs
V1rP6n2axWaWEd+n0ee6kwVh3N6iLu3yaYfzVNku7LouSTFfClT4ZtjXRcQrYGvyaBA3UoVnCw1N
PiC9QCLBAtDfNHp9pIx1DEXZElZgOM93wmv4E0+M5jcTwdVKrLONbh0Ia1ZWmAvSuvjxTfulNvk7
8b5YK9Lzxy92DHs9ZSw5msE1Mpzr9jquxx9iwKpaXnKpU60u7o5BFdyIYbeC1QvZhDVw1v3kVVq0
5ZDLkDiVZAORf2FlA48a33Rrvi99HagSOm8ZfZOh+1yDjejFyUrm0tMuGRBONG1Q0QBJk9E51Dcg
456x19odA8Rok1uDmmoByhq+uMv7tyqfSHHgM69ozc954FujM+tNHEnAPUHrDVgF4xtmjxe0NRdp
2/D1jV7/TE5IVlWOcCygogULkXG9T/dTTVxx731T7YBCn8gcbX5TpX6BGSCYxW4pTrloou+2N28S
CZjT8XlczNhi7CRbNe1lYEgwJ69Fux7zYO7w9CCNY7oY9foXYcTD/DgggIA+wao5CqRvl56fg+5I
HHZwFUSpQsFxViO9DPzkINXsmR5CwtdjCijLD4uVGTvIcrHNZueedBDhsY2mcL9gyvHooxmr39lT
pb1gWZgV91UaAUFGYdiFoS9nDvlkCmCTnXZLwtpG4KYEiB+MMeJnPU0qjrqgwz7dHdAQWISmIh3H
j7jAmMDREtGkqtSj9hOuEMiGkdcaS70oaH6xX9XRTAOH0LBWQnKR8LtOAKWFo2fz7Ek3Guxj/k6r
QRkatQZRPjdHlbzvMrR7MNuaC3cO2/zckpkWEf9igdPu0RtCgv444iuGV6eeKYvWMpk1+1w+Czmx
1xUsrBKJX41gxg/1R96QrvxYP8uPKc7OQyzFRHMCFmtjPi/Y015RWVEEOeSQExtAFk8d/T8pPzME
FCYTVtoIafPPivsIKyNnSKF7WDGQpUHivXrxwhotbrlThN2rC3xEHQdH6KEZBrAtWnrJYHFcWywA
Qc03L61fkSIl1YrAdCqj4aoDnWNFTyS2B1LHY1WhZwtn/Fa82amSKFUjT3ZX1HGUORkNCksGgkXn
EfSDA4QrLZMleBoaA6Vbn6xEPU3MzS1eAfoY3vKo5x4sSwGCtEgJQMxZLwkFCWa19178JgsujvNV
F32F6hz7PbbWk4GbyqOQgWs29cRSOhbdC9iCq6NXSd1Qt0lYhqK7oP5Iyvh7vPBidCx9CPCfcoHs
/MNSbAhOkO3Pn//9HNMJvYa15v7fELHRloLNChjEtl5HRw9S8hauAGl9EoclzEv3DmEnPkKSgiv3
+0rhGS4YrwhhSbJ7NyDQTjsS41cveGarEcHPHtRfsglVj0DFqCa4+xKSXoT0q8VtJ5AAxz5Ez8v8
hPLsc+AVid3Nr94LqTELs41qM/V8TRQdzZZsE4pR3NPuhZZNcUGgoGcctQ2SysDGlT0lsZYBpBxJ
SGYZ9zIWVENB+rFVtLq9+Iok7OURJSMjNOCV07iyPi4WBqE616/X1QPxYsM92sU7mry4sdk45O5t
fxs/lJ4nDQG/4CZb6ILHjAWjhNYFCpQ3KUzP+azyIoD2HgtSQ8pj4L+SXDrqjkrW6xQgBJUoTkmF
MckGChP+2yZwbVoFpWARCKbqfymZAwjU2cIlgm7kwCszGuhq1uYBsziIy1cObYjWWcXuAhHZKjib
q0x+/ZRNjcoymO1dCW9Cs+CeGpqST3+dYGYw/bas5KMCXZJ7ExJurX9z9/twBhGPk8UqijqDq9EG
+w3yvo7CYMAXV1oExIcx0zxLUVmoK53WX+RXN5xzSvqm3KxaOJv1rRzlcnKBcbps9X60a+Z8pup0
spLoZgFOLNzOPaM1aV5XAsIjpZhL6O7n6QBhaVBkcFa5x6ev7NWgcpvIEHL6Wn566wIjoA4px4bK
/HhO0x+jYcfbb1FtGgEmJ1iOP5hV6jS55ZkW9P0f/yXBjudtPJZR/gxgOSM6ar3ZNQJoxZQJhZ2d
8Mpz2ypDK8H29UNldXs/CR6FEtri212uztlqA4iV19GD3wNbnaRGUtVecMboQ9RozmC8ZeCkGAPe
Pi5pxK+3A8nA0fi7NAJF/kI25PSqq//lLp8r+wEww+f14Wemi6RJWSQZiAB8BzSCNAZBnnoOw/dV
TVX8px+7HfWlvXYZKNLgx55oeuMG7FoyjhuZXCT5Qtkosb9dI2rR/T2IBkF5S9feQS7PwJrmvxBd
lkrzmtwNdtxrZX2uX6DQiKPjNTqllPSbTb6IPrLCnGT3peilFxrTcccLF/D34NySzDaBiYKHGfcY
uhCfL8g7JxFRddOQldca4zm9YdRzi/RnutyrUDYCAWQsr7v7ValoY155HEWZooe3w2rYbTjduIta
aJO0zs/HGzCSnlkKDL+IPxeIrra+ZAwQVyCpuaHHnsPtjKMZRO2X3Sfd44IGAQ4oGAAi7f6jUPxx
bjqOzECnHi0BKAkuHSdlorOq2S2/aR0ItJqTEEqkPvjAVkl7yXe+/dLo3rz2ROci0hMIm2AQG6yl
0FajOq5VJcqRaa9g6n0TxCQVcf84F59glLMalSEfUgBD2N7Ah8EeqeiSt8JfDpw840Y3O0lbtClY
ScaD+gyo/4l636Dtf+bE6ztzIci2toPdP+86xhtaKl/uJmIm4NcZMb4DCf1Yholz8a22vqBrESV7
Tb22SjodzZNx45KEP7kV/g2Hxcgefkb41BJpqUrLRN2p8zY64uZGGEq9RBqL825/bD+sINBKNgzR
cRImfPyYv+cLdkfNnxoHBDIMPnqjCONtFF2D59xdZ4PyejI4IsBkhgO4QUxPLvqGUeYvMWYgaLA+
Sgx/dwkKhIn1IW8xghMdD97Qvi8HTDJG3zqhsQR60DV67xtKR10lTfIVTlCdSP1/dn3IULC4d9Ib
Z5hQKYRmReFh8AeB2rw2MofF+iiLwbxx0GPLeuQTxm8OFAIW5TFbH8N5Ub8NXSwyuhFmqvoj13pp
xqznIXRELSGCdXLll/1bVgJoNPoOs2IjbJSehkKc5orDw2cvMvSyib03wp7v9+9psa+xXyMA0f2x
McZ+mPu/fileR/cpxtzqCbXKUfdIahT8NDXOC669Bal9isGNc/g307bE0ZcigR4IeIaBdlEH7Ts8
TNv1iPOOes5oVJBcN7RJGSZNFm15K1iWSinXzskE90HM4TSEY2lb6a0TClyN7+VR/BVv9A3BP6M3
QXq82rNwvjmsiAjthm5VAstAbWAyfs4le7YMI7kwT+CxUUlAl9PYLgX4CU2pTNiEusDrkZj1MrPf
gNpuAH6nKWgzT9TPguYs8mCe9MC0dh3snOFNXwSlGNPQ/7WNm405zDbPAbDdju8Hm/VwkcrFf3b2
N/jiNd7trLxquHGqzlIDCsXryT11HJnklvNhnqSbYALCDH2FhaEFj7VhQ9HlPjJ419p1vn9npsVe
JS4h98CorfOpARzM/iuPzrH6xJBXg+hx3v3kBBx21VGTdhWp2d6q04g9UEqd9poU7zJuBdcheICj
GpS4foz2WkVVOPIoAoXAbTHxkVlXVpphV5W7YXGHf39/UoT4nq9j3+jGWot/sv/+8m8zvq5tuUZa
6PDp7BO3wD4YKlFXY65W7IZwUkaxvdTXkrZha6udUlUYMYZBKIoZijFtEAlzG+QETOngRVbIFhwe
8qMoxPzsMVNf5DO6ZwwqCBZJoRjzeFkixwl6u6xVeHqbOP1gnwcn6bXszTuDxIlrqnrEVI5AXAWw
yynT9DWfzkW0t9X3JEx/Lec1xj95t6gKd2jEs8u19HgDj3XxftKzyQRqPw6oHqx8xjI6UH0+pWB7
N9mJg/SJHMa+UNAE8AfXAy4oO89M6Ypr8+vJx6tF1UNOWPTNhnD4lmsjJ+PXl5Bua2s8Br4CsSL7
mebNtJAr7U/rNfEM3HTvJmWIVfWLeds7NG2njh70l6nHcXaiciboMFTT+7MYiF590vMLBeBQv2rN
RBaqP88MX1qGf+JGPluLBTd8DQLPlOXglZCdR2qjZOTHo4XD3MN1S0z1mxJ2a/M2W3p6jPe6Gx9y
9SkJkPxG3PTq3CDjdEi2FxeyX+2Vb2NteRwT5UsbWd8EzFtL11hKz5rUPXDfHcvz7S6RZKJeBTN8
vwiKLy7+3jh7LEdbu8+dx3J8Mr23QA6K2WhiBIjxoL/q6Cjak3td665Q5nqyrTjXhyoaXsqQ93du
vjmUV76OIXQjVMdMdZeOj0QxHF7hBgGutvVf8stky6jYd5xQYMm4euYPYOQ0M0Bd4e+V/uLTwQbv
k+sPKjETG+eEpyfVOjvjw9oud6yaOBCllin6iTJssAc2W8OwIl0mP0YrvYmNHLOHDf4pTTpqTZeQ
ynMuLlsau2p9JOxJeIdRZEqPZ4zpJlFdMezRmqvNISL+hS9sndIn0cp5U/4W+gq1L3NhO3fUHWIx
P5bu/Gi5Awd6aaa5QIuZrSUQzyXf0E6GNKgPZx7TYMoM7nrrZq8m7mUO07PhtVudLsLs7yJ0lfzA
9Q+lnE1b7otCCo1fg0etENWupCzEqlfpdVgiVaEBofDZVXwo6obsj+34bDz1kxWucZ0/Qy5LPAYf
N90bk/qjD+3vuzHSAFEGZ+dwv9HwETzZUaidwf1UCeaC8m/3p8Q0ykEOo7F7VwTDeVibPHxFUMh4
Q0BQtDTa0rbFqze2JTBO0VzgjICuQGuA1Dk4JQNEeTmQIjXDe2H7CxgiTCq244GBtBm5s9BABY7R
wUVs/MN4JYVJV350/KVXtCdgnZ5oQL0kJktJHwYvZIlc9RG8fulMMibwoZ2+qIhFYiW/r7Q9XEFZ
/3RlWURtmZHy5ff5MHn+PPZEWFsqvmzyZFg8E1oiVtcHgy4RY/IG0mnQA0f9rEVDZ+SRMUTyu+cJ
+0s5BF4n6sRXdN/UR4ooUyZDN3ktD+i7UbY0UkJkKUDwGvoaWCPYTJ5qusm1rn0+zbs2zfEL3wZh
CiDhy2w42eLOy1J8t5LbU9UlmXbzYM57cM6YnzGqfvM2Y74VmXZhT/HUyWCWGEz5acwWrufgVs3u
w+RiELhB5oFeYPz6VS7x1138v7D3PoR6oGsPxWgsFx1XxzhTjNUpnpv0g3J4K7F99/ohbLxz3LHn
vrpyE273bTopJlaaChgq9+kXEASUtUmLLzd040EP/46tvVOoT7lzYC604MEVO5HJXs4Evue0lvD5
1T2j/VgaMKv0POJ/rOiJUfoqP2riGqWAmt8U8eGC6f5vkdgFWFAeUf/hMY3qxY7yEIS/h849InE2
8D0s/hIaDSwN1xeOlgiSLNHAmkLayp+FIS+daY9Ss3/oVMJy5cEu3CIbZ5VUYmId8ZdzO104fQoD
Or0Izqh6MeW72pdnD8ZwbiyFzMMAs+5Jl6+KNE5LxJq9W16piUZT71Cgp/iByezZtYsktkt9bFsy
QAG/cvoUrrnUKLs99FgPakQVAWrG3WnkQU4TEsXSsw05SdIJjjf2ePfv55fKJp620073aKGcGRJX
FM5FwQp3wZewZDjkb98hRrRhSi6cBpxHYHrmjmHhkIEmklJ2gOgl5LGTleOQ3oYlFNd8bqUCgrhD
/Og6lJXfuvasG/ZW1y6eMQ5TR8rZIFVXUVhMCAjdG29EbhE73mAQ+VdHQlt123V/mA83DmVF3sjT
G+kI7FR7883iov+7pg6mvlfZbKeUitDQ/rfj4bkgN+Hn+K/zB1glWntWKRMgZFEhZp0dUFcyGBr4
XUdy+YRLUAIy475JK8y14rOttRN28EBzkdOnE7RGqRd/bZkJ8yMq/04R3dj9qMBRX+a5QcmrK/1s
zrGMhQLTavKD4H5SwMoIjkkPEaAkbYCANnOETKiVSdf7/plCxfciAWeAdtjBm7bcGM40GlmZRnT7
NTAHv2jOXxppYcuZPGkbifclQNOEAA7f8oA5o+m6q/dbVqA5S93nOhnW6Gx+rA9C/4GgtYG/CRwp
1an6rBbplLfqHXBtIbx4WQRFuseSj0mgpFNw4diD2QVO2J9hMwFa0HjsSwYb02Gjs2Y5kZkPnGY5
d5TNoOILfSg/h1KBbTcGO8pjdXxsn3HYSlFbQ5cMOXyPltPMdUQsrLmD/AFj4z2xEgmP22DbcxdH
oExP7rPMGbtF+4CwXoHr1o7rz/C7QFRklGf7atPd2MDl8eu+OEZfCAe14kTqnQkjj6eRoD609qtM
j3tkL30zhZ5/KPW+C53KJtQz3/dy6Q2LElkLDdMGM+VdQimJ528G2m17qx11DQRaMp6zflJwXQNT
0lh48pBmQ1t1S0UGN/yvlDlqtIQ68fVQpJWQqQ3YuLynUhrOPg9wG5h3GPvwRe5mpZmmnhsFgu/5
509gIdTk7Oyp7GFd+Evytop8/bWDPmYKR38Ij7WIxg9v87HotQ6aM/iP5giuhxRK2ynDbFuymk6a
KSbE5UGtuFtB/qV/hXQu8+tSi7zc+iyh43qq/h61N46FNqa1m3Bc77flQ5TjYi958bBV/6iEfm6D
Blf4UHSh0QJDn9MIJNmWaTsJcUN8WQJq7lEAGV4d4tEpOF3vLI+c6qX5gXpYWJ9WW7N9UqvUzHSW
uTqYg+tiBDk+Hj1bheEkbx2zVsOUYdyKdAzucQGsQTDfn5hlWo7fQ4dpcsxkhHtSDdCIlL06TYBh
iTUUEPEgehOlkA6G6MQxg4rFHpVLY+nkeJttnfnMvta6Ct8vFxM43iLLAPlFaw0PUWxEfYLUcNwP
Jk//zcj0fam8njlLB2sooaayCa/Ah9vJIUG1X95fZj15j9duAmnIHzKEyiYL3hA5hMnzUGAge+kt
35rcE2YUxb6twBxSJK3UBeNLTVp9hl6XbfTxnLIi0A3uXWxy1P9jK1ruD4wd3YRu2duDFCGXZMTn
6TsWMKHPb86vFiJ4+FWMwZwinu19H7wz9dxU2KYPYxbpjzCNXHtLJDmr35bpjCitWQlR0pGk1UxX
1v7si/EcADhUUpiltczVSoQWYX4xdY88G7dqvi1tPdBbVoBgsa3v8PHZUQVqR6aKyGTafdzmLd7h
4mpjLr8AdU+eyAg+ZVXNJPdyN8eNZ3N1JUZK5Hab9KHg1dCTjnBAXpxXE27Jg4otG/Xc4jYRXQN9
FJf5Hl57pj9uw1GvhRF5fJWCbspfgwXSiDK99FrPozxQtO5s+lsK4qw4aNoK0vY6dxXkmMAdoImL
Pq+S/CpTnx6ThEN/RKM8TS/ci5wauT7w8hW3sH6sfKmwdl5N88NgOIl6E4suZjJ/UrBYrJUMPAN2
YdHrGM08H0eEvkp+QJZSAM+8KJ9aPJpvpBvivBp49qiTSN63MZwT+c887SRSqvdojVODcolAcqQT
lw4rEQ/+Z3qHf2d921K28QtS2U1Z4/mfeMYUT3PjFgbCd++MsCzZUOxCD6nbh45RZuJ1ywq+SpnH
q7aOQhKUyFClTetu7T8CtehXYlkxhKcwlA083MYcNwqbhSCgrxWYk3aDGIZv44eR7KeppbEdxOvR
UXHbhEvu+FTVBpWjLtyQN2mKq2RPXctZcfybY79LdU8SGdw6BafYKh62oB545ithfNayOi8H/gZn
L3bt7fBLyWdKOfo/8TjOS/Sfg4J77l0/5Sa3cgZI2a9+K+lqYpZQzT6rOKKVTOmEMjjUK4klCVH1
ceI7YpYXsEU0rk8RPY2f0MzdeB06/HVBEG0vYyULvcP3V3zrpXUHh+1Su8RkMRHTjeXiBRw9J56y
sgHTsuT9K+5vAopPNWh676u9hTRAyBo0Klq5B0U9Y84iVR9nMVatbXN4Nd3m6sRwUoBDBFk5+BF+
oqtx7Zt+TatdY+eYB/NMSV8bIbfJoj6MoFQPxaFY9rcDux50AOx94ifWeHErFF5RNAE0fhHjeggz
1V670yjZfJ427Ht5ZUcpCvC5XWwd0ekZONRa1vyup7ssXaqdkF/9ue4LHChYWGugGCkkpW8gP7cp
DqnHPjyxQxlr6AYschS0reSj1z/iattwpwID9VEAMSLUUfKosNFrKUJqEd8+z79K51Ib/nayCP+e
5PoNtxv398FuDeMMjrlnuXaSK2QzM7Z6IXCDJ2csXV8NpcLy6PiXqICQzvcXMSemypWpijgavOnq
aVLTzHuzprMLZ1ZgpYHZFG2ekHL6rTYUi/tjXzRUUfFs+GGwdMlycE7owtYkA6BYF/2NxhqjSkpA
1GKeH/ci6LPJRhKUKj/v7ZNO0bNrTJ7dXezcE7WPCqavFYvooXeRLUpg8xKOSmy4EZ61IfsHhXZG
Bkahh6fUUd3LlM9I4iDqBkf4/Bj5s1MSPTiu1ufQtHOu2TQaafUBBZtTc2dcA300/s69VqFR0Il4
bCj6EIrIpg/ZLiS5y4nvwBeW4oiasZz6e/Eq+zR049Ibfb4/US14ivm/tR1i2+G99dZWMB9VRwFh
WnEmqw0zzjDOch55APlXZuoQmFxuTq2/OLUoPuIr/5LyVnZMo/jwu60gv9JO+x9WFmGpQ6+AbZ6+
ox2GcC8sKzD4bkMmM06ARd14tISIwew8WW/Udak14fGfZeXRieXbiWq+uPM7AIiXT037KBCGdkaq
TgbXBex0/obxunrIK2Hu3hm5A6eWtQRziRbeTZLOQiKMrhyULfdSMrHbiN4gs1PsRIfktcU2oG+A
O93hFhCuWKfiEJpea7T7Gvxd4eXcWQSqtwyXdry/JRkPP/2IIDeqCR1B4YEQwrWfs2Vv5OvMXGfh
jiG6yr6idInR+gXDLzD0Vs39/E5HP6VFgfDHAg5wFA9X/d1kc2ZkdBXCj22CjfQmiVTSt4wv7kPv
ZgXOv7s070JOtVA3FUm2MnsVKi5UfQ6R2YcRDpPktixIeAiMZYYKvjP643e/VsHW+mL/LbJayflN
/yBSzHBqhJEwzPZLsQAOuEblHKQKgK4Y0TFJDbgquYe3oOi85kELs3VofEylDY5QzywHsmIXbGFY
eoz/MQPSxpP+ea8p2ILA4on97Tt+cxHkuII3AdxRhB+C5PkbVVGenPfNsSmyeOFrlWu9q7nlvIiL
Lacfwjys9UNJ+gIkvjH/8CEH27k6BnUlj3lGOSB1dzKdaYSIfz5A9aX0ThDpwSqdVX/XpACEuuAy
/5LRNtlbmnNz1nbZ7dMrSLD8mY8OBUCIOJNRBK+1pbzXPakwaHQYRWDfnRYWMWr3TAi7eUthqzz3
nqEipFl7l8ITrW14O7W6rnEFQi/wn0FdjS72ebcWQuUYQK627yRV8KFPZoC4UHEWIuG8OCt7ytQf
t+qUrHbIgjid5TK8qBYDimKj9B+3UjB47HRKw5pOoTPPRVkHQKoXLXBnotVgJvBUq6nVDaucFKyz
pkvJUAN4PwT/MtlJgB8nFzD5QqGGvduKlOmMUDltUZWVoSOAt0Uwkk+XLAuYkpgkuNLZvjjQO+mZ
rcN8o/OJ1HImxK1jzIL2VcBRKKgOBu+NVqi7nu7XSJw6NzY/9We/jBWW+rcJPImgngk7z5uGFFaP
NV+aN1h5N+gfckfEO3vo2/3VzeYYc3+B29Q/AWT+y1kWinx5zFPRSoYx91clmFPQjjRUfs8ASBrN
6Yg0XUg9zY0LsO0+15X2Iz3VoHah/0TUTL9oiblAFrowng7arhLRGedjrE2ltAKDnjP+ZgmzlkA1
3RlcTTgtrf9tSNtLFc+KW/jDu2EslU9ZJtWmYz25v0/yJ/f4ktAKIqT5L5k0vjgfQ0TZVXnHRxI0
SqyMlvO7Mnhuqd1vWauTX4T9yctBt9IG5faA08HtqoXkN0BHKRFHF6P9jCUU00W3iwPd3Oi0d4VI
AjFXsqqaPFAfahnJ1+PlM3pUc0BkTgA4y1h6CooikbESpg6A3w2O6cUNeKTPka5a6yqvNo/Ig21B
g81YbnQlfgQt34AxzaAEn+PlRFdZfnvg3C89PAvKPYbRgU0ojkFK+EB0Hk7NisAkH+vjQ/suoZbo
aK4PMpE/P5L+whLg2GEZ5fmWkIAT4YM+fSbrlvMqkc8dbVhJjngGnbq4hhTDn5Bm1EOgarjDonqW
exW22IgHd8edTqiaDF7mDlgmw7GQzOj/WnqSWKVTU1oe/8s4YS1uad4/nqb6Gx1q43OxsWWsgPQV
0qo5Wzi8nSXlyBW094+fBCv+wc+6j3m6RayccJwq1ZAtvRCD3R0Z7CkJ0BUupD9ZZ/08A2zX4iMO
eEJarufjKccn0x8FngTypgC0mn5q4Jo6kSqEctcnYRw3Iz5XPSuI9p+YCgWgveqwXt6i5y9iI+XL
EdWE+7u45/aU9Kyk/I9cjE9dXJBGAfI/2wCYIvhzB7VqhWKnTT0C5nVBEhk2OllBggKi+1YRMTDG
G1plOB17iIqXdDHRspgj2nDI/DkFGwzE+HQDp7gqsX5h/77a6qsHDjPOv5Yf9uNMbmKMyuHBINPg
Qu+9xoNpetIF6Gs5zeOh1dQZPlfs1ISifReRTn5jx0n7CFIrGzPbBcBhfoHa1rizTUDANM39kWZu
RLeNXE2Ku8Dkvk2b8XlQ+9TrUDoA74YANXqV1KpZ5sNWcrTYNtGXXrz/xkLmEchEs8J+UQnAovSw
hNfsC01mpzqx9qVZ+2TybkzNBFlnY/2ANPVp2FwjsQh+zbTjbZtqWAETkIxAIDes2SlZquVjdVLF
PQVyuLgZUpEcNCThaybo+ncEc9huqkCd06VxWjf0EX6Lsm7btGUhE7pWdWdjaLQNSoo0uAjDNt3b
dOTOg00STHNosp3lDQWQd0MQKpfXOIYuHzmadwfKNIa3GRPyogHBUsKpTwyDuu5FqjO8YDPMhx5Y
zfyKj4pPZYFjJJMRcj1iq731jVdzkEmhvCvjSJ53CJhZirabUYsJnSnK0yu5fjUVMJPaoIlq1qnz
+alkOU/tAadOM8v20wRoq7XFti7RgbD/rP+ufm8txmHT2Nh3Hfi1KKLylZjWbIWAN3FQDIJ80fp5
5E/1vZRqAs1qNA6jfEHOD9ryX8ByaALYV9TGyyLGY5lcqZxWT2w/AgJ7+r/IPFYgF68xRVg0RrlO
PMjZZbjEt3tA02MlkbrD9iOZo1aTISuBz6BN9Hh+Cz5pdk6xUT4FbIAhtNP/Zxz01k0nq8BrQQMZ
s+U5qlPamPlj2VA7gM6x+tSYhrRBQ06XdCuzIA5ERbuhQ2D7uMCvKEYdX796b+5V491WRZoL17lD
1QxjZzlAvLShnFSAhPD2Mf4SjXDcfHgTKN45RCTM8FOcM2vWP0ow1B5uh6b256PJ2xreUDMm953U
zfiyuabv2hsPv8HrEe81eK83Ibx+b0lIWkV8jNObxD9jNQ+WvZgnNfIyyyA3EXk0TSpZb14qtWto
W7EkhCp4nqJ2NwPoBWC84hKq8JoE0ofwatbkyoxoAPrpG0q0tARr+Kael3OKr3Y714dyifSqZkJZ
rk16jbnmnktw72MxjJayqA2qDQh9NXCx1kdnxA8TXG6EQPo3Oixe2zHpYfW5c9nRC/kmmoBAosS+
EKdfT4Lcf31/dYIAmijYr8puKUPXWRdJ1MRWDuKr7Us8JXSb7/RWj0niN4H1S8rxFwchG1GwEA3Y
2QaQpK6a0MdvYsaLqbpUznZ/IW6hG68K41QyZUk9aKURylWylaubGgzwbXGR2WLg7r0/xJSEro1m
sUEUARf/LpGyaIemdaHh6uqgBHxTbnSh48/JQlEXnzLILxmxU73LezCv3L8bi2RphRfFQfoeNvDz
P7PtF8NefAlNr+nm+CAJxq1cmZPMjJndnYY0RcMnUBtXQYvZE+vMDZGpcXuAw7H8pKpy/AqIuy3D
yk9PQBWDBVZKcDMMHgSZqN/eFEXUdGY3FZuLO0S4MTkl0KUrENjzQ9aiIk/6GjT61dxWPMABJ77n
XYHNn0V5c27yOzOpyQS5/sNqLJDfCFLXmk5yxpZTnLezngWF52juOK+BAMB4PDovMZtXKusZq/7E
mgvOh1WmqflcqmwzP+u3UPMub9Zh5HDhgT2Dp+KzfnpXqMm835PKQBlw4YpatIUW/AxYACgeVeT1
Ew1OVf0PejnNw3nSbxLytboEdP8VtnYQ/ozVfTHajezSiRgKy5v8qaPqpPgtJTjQ2rcn+yStIUog
MrPmQYq0+BppLQCNohwyTZrt4Ryz7+8MLYD7ss5dwMR5C4u8TI6UthDCiwviQOfnCFtsd5ajLxyn
rzR55yzGXJpyJqLHWmjmu56aLTDd+55WY4Qv2qc9pYS8Cs801JZyidFaRKgQnHiiJE39VBLLBlce
cF6lGkt8tBNiNqEqcNsQ49W0Z5B7Pep6lZ6Y/BKtQBuud5QdMmhqzSsmV23iWiRr4XEzqAPIZfNk
kMH3ogK+Omp7fjdP3skpPBDFFvoMf830nqQY+BNQBEISXc1e6/n9cjYkoEXBr8H8wA5jo0TfQRHJ
nwRm/9arlYGZ+nfJFflhg/o8dGleNqVzqRA2iiYNKV0fCkWs1FiAKYm1TjDxndfcT5UXQJRTnWAe
NKjy+cjR3oq1aRR3YANNvq3EimitFxHIM3pexWMjUNvDzvLv1UfYnOW67DFa1ViKsUMtT/dG1V/L
4ocBIzPrx5gzIUeQOWwPfoBX6bigI8kbMy6Q1zC3hR3xTVQ7FJqCkhvc7wd9J96qERCVOl3hblkd
5lSdEXtco3dA6sHupynV99UOSAvQGZjRMe8AHQKuOv6CHkPqN28fp6MJ1uhyXNBztv1b5iTmsp0w
QpIH7ZAnGBxl9EGrL7y8QFzpVD+Qhc3rYex2LfbBjJNxgiNS9HHFmqi2WJLKhtHqfvcmAuf4BpND
t/3gFCOHNAIhT8bpZ/R7BU74Qvibp0FzicmW1P7G+9+3A0jEjf4eQORu1uRiPGSK3CnRJzMLOKGm
1cIBxzoNWW++n5CQQxQjgYMY25yDcIM91gDvpBtzOrcBSGhFt2TRR9HAwbhd7mDEB3Jb8dr5H9qi
MWl8L4g8Zxx3Bsm6nUGcHRSRLp/jn8cLCd8Yptf9zIEflG767BEGe5oq1FXfr/l+0CrqWIvDOBcz
bOstXZtgrPopkTJdjMnCgNUlwlxJEaoIOj6G91fbUGaaOotYHpHy1cxEHO8NB0ETOuRtyQlBguC1
7jkW+tzPJ1wksPMePeE+107lOianYkTi89VraaOTvpCy8uTt6Z8iJXmlxtCiF9YyiMziBPJT77T8
AkR2UwxKBy+FYvhWd8YhoXo1TEHw58Q7QhssezAeuI7XmaJXEp6qOcFYQLvyVDdyHjBzwp16yDiF
KLYv/nV9G4DD9S/N/m4Iud8JzF19q3Kyl634XUA3rPEr7Mv7gFiDK/6CS0Njg9ytYUIH/atmpHRy
56DOnQNSn2t4MjIxLJu1Yz4VL4PgODB+Mv6FhF2zzBuMZYL4RtX5YY1MhGVug+P42PoY8iUbZG6W
RO1xSUafhg5PHNdjVBkgcvhHHv4S9vom4+BQlTBJJJNaLc6TowmpVocSjdDwD3Rcy0m7kMBq7ooR
WVs4sbN72wkd2tBzhlWqbocdU+wR5LKnPzBKT/vzD+xKpmzZyrpb+/rPPGFkxmAuy+nBHOZm1PjW
TEyTfPCLQs5Ir9Sa9ERUncYSwy0FE1m6O+ANGBuPvxm/S6+523+forRsOD+erin7Oanum71V/Sbr
XaSxUnb2WpFvEdf7xin4S34XPgcOh+sU4IKcXYII8yRgwfQiu7U1246g7jqu3skyy46lfdadpsLr
gyyNpvpEU8dxL300KilGqdTl+itAmCwe6U/pZkBwnqTYv0CNiRDBhHsE9ayTZyHXrMezp2J397/S
DHkRXRPP8hB/n7NbVi3shzV+Oa8T96TpoBQRYqk6rZ65ZyEVgFDlZsObWWC/D7b0yg90nA5ING45
RTzI2jqtWUQCPb4yviQumBbBVNVXElM1TVsxjCxq91/KZuWFR6W778WhFRHQDyTYcwTIR3Xpaw4D
tx0zcnC12St/nJRobZuGMp1ASqrgA9AY6MtAH7ZUEN3MbjWhFVwBwtFos2KVkjc0Gf0LMHH3704y
PnXKmPplzAkp8uBgpFD3KMwHbs7MAG46TjpJuV7R5GmWD8qo7+ls0jOAARnDCXymFyZZyhgDqhUX
Ahzhw7PZr4bahD9NH6fD67X3jHmTpfqW2ffpNGcxVgh7t1SDRXFr2gdYqxmPk7sf2RvKyaO69cPk
55QCrVdH+tQarYA/C9qkyWh3SKlX3VePpP2siRFdfmDDwh4kDC4WuCHgeb7udzcc6gNmhoaGVj6R
89OoLMEBvmSZkcLjND1HL13km3xzZGpTfT8ndcI1+mXJNAuB94JulWIvO/5v5fudEOHDSn/PcUGc
bWV4HJrhtNX+C7RaO+rFU9iCsj2xKqyHe4y28kMPdjBRWLU4PfIbQ6ijr5woQGX6Mkldp++57Ljt
wuJ9uVpuIY8D/ZvRIKGd/qvuOlj1njvf6cfy2bFeJoCJjsaIVZ4fGX0omkyNCxCW7I4XmMyVpK3m
XyR0NCjwk095xgndPOB8ztA0tBliU2TFlXDP5H+3oQWMqBFH7SMW0BkznMebF7CCZaE7Z4mMJAot
Y9BVDpkMTYw8f9XccgUnoz+5LOpgprF0iqlslw+5/b22QSRsgg90KHfWuFt5abvUw6vpeQSz30YL
TpMT9fRhzrfXQ8wy9K9C4k1EvLaJpvpLg4xrWb2JA/jJrnAmaztESlIXoB7l7iANdahQk/WBnSpk
sA/ZnB24zgSOfrdPmKzBR9Q5Z/KchyqK+lSfRSNnAaWKpLxU6Wc3NKg67JoqUpp7KgtLVv1nd641
rmIwWX0xIX2+guq5jEh/ahgSWauDs/7Du94/HDCVlnCR2Vi0tg49Qd0lOk8oOxtzC5nk3PGWP7zZ
kZxVxn9eosj1St4BBgk6tXz4/5pHYQlbnXzx/vNWRWyxj1CNZ9cXETwVldJ2uuobfkvblbaFt8YK
F9mvU8LsVDlKphWyNrD8+ua9icxB47IOJMc88jRJXUFGoy6SVJnobS4o9mq1NkgR/Ly9davtd+o4
gTtAZs+pCnPm0atdlva9ejHvTD4hhHrDIePq5/BKnBULq6J41am0cx4nj28piy3Sr8weKRk1/BQp
4bqkuQPOFAcZB5Fkrxw+jUJao1ExO1UuriVNb8364T7okHM+f9xLKe2BswbHfiWA1M9LL+LZAM3b
eMDVPb8xWLLFb65yv9bW2gyLcci5eOwserSSgggivYZyDmUXx+EuPm4Mk89caTBfagBs1Ip0H25B
a8GmoMGzAfRgpyKts6Po/2M40NybCpvx2gPjxI7JAFfn7CdEJYnFYhmk6zXLfuJRPj08CBX15qaz
b7Sv3nlgis3N9oUqsZZFvL/IMpmfScOWJwkW9QzhXaC46NWRH5WAt67LN5gMUU60EdI7qdAHvd/m
FjUyR5qjFfj0T5h3xOqTXe+XeGANOYLe5dUcXBBy6QiWKXHQsVuD6VPQvNCJVPuA1SVv8OjENQXF
FDyqYVtxXXobgKTYJ+OhsEeJ1tkYCu8FXwA09oAHAnhPdN+xZZSIFYHnQDoEdWHKzJ9B8zTUdeAV
yZ+hDBE4UcJXZzLEIBC2HhOw2SQHWMUZfNkwCXX6C/g+hdWdh13iTX+xjWJuPxB5rh+fJQpF1ZvS
XvNUbfhSv3G+njD5jBIAnbNdbdqYiBdSQGGNTFH70LWQfRj5m+VzfAAyN1Zt5HzMziB6jtrmTa7R
PLzzH5J99WbjE/17WY0b/V23O2x0JxjZpZXMqhdytqmbNiQOSNyrtI40uIImLHP7t8F6d86cFKkD
yXFVhA5ZpDY3TmuB6DlG723GcJaCOnKLseNZEsA5OPLz9lUPqWr5Cqb8dbQZrtiGgUF73gnNnkgC
Im75dEZl8H4J82jCiBBSLUx1+JxvOwBSvEf/+6Il2CntDOFNN8PqQ3kDwejVOY20C+Uh8nR+//e1
2ILkoevBvbWAYdinsm9C2rrLdfyaZ6OY7FOY2y7FZmsZfMGpM67ToW6E9T323xCtNkcSZi9PjMKx
nlfbEEsRVl0rCDVg/dsF9/hQfrn6UoXJOOxSdc53vmvGB9BJ9ru69GeY4QvHYga5Lcj8l5rW0Yue
2X2lydP2tgKNNgQRqN60dza2zTtclTGi7+f51PWrOIgD9Sw+SbIYHricgaUFURbJxDIETMnuiusJ
bPFo88SDDACmUsARDx0QLGgZ2vWA5376yRGz2BFAr4a6oK1Hdp1lNKhKpF740AIlmYpqONxLXT+z
gl2y8FvTTosXA+j+xqBsXKhoyrK0pf+JzNAnZof4Ejvx/jOCciUXjtlAEysN1rX2mq5BZbWQrfPR
nTiQZ2eA3uMHBdz/lNCzId1bRs4nk6uh64fLWmoVGLjt9l4Xzc0oPV75zKOHjOMGCFJFyVrwL/Qu
Tc64kZDJTgIfpO8duU23PMijaOPOVp5pzmoOE2At//jfMhR4YoAI/UAY5w97jQf8bP0QzGjm86G7
PA0kuARHQ0sHqQ0jo2PEfFRYek6Es5VLWnRPCvgXrA++xDxpul+NCQ37P9+8lS/SxWVTJEEqmmK7
IAVDd74RfuIMkY6+5I4eZT8h8h9fiuOVeMx2g9um8E9bcVPB0IPfmf5WO+Vc0wEKEmqrgL5HKY1E
YhAz4wJH2pPXvO+CDJyaVGywhDJtiP1GNejaG1cnCCPlfdMixY7L5gz5L3o/kwjOCWZpPtNPBQdr
RgxSHWkDR0c6JaHQq4m1i+avwUkS6ktxt6yqaVE5fOMsSetU/6PrS7V+38tbnCHS7ul0Ed2KMZSK
F/1GXvPKxX0LECiYAd7QpoRpT6dT/l3ISBzwltglvjTljv9sAh330uUgR3tOh7zsUhxwRbII+3+V
X3kb+T6phdHoRX8e5EQLizsvbY8nnsTDA24G+37CffIEfNL4nvdzFXRb5SkzhvSJVOq8MVxOiRCH
AVuQ91w1f+wu0mI6TyjRh1AGF06pfxw6yXpx0pP3H4XD9iQ4v1HvGQVCaKFbQTPNwiTRDjpKXiIE
u6BRFQQRi9Qq1PsYHTVY3+rWLvB8TRY0RMRQiOwZ+1pcT0zUpRGvHCFXAwQyxzI2bYdb4y1TMwH/
3QAuW1Vjfbwcw0m067l0cv5oUiGsjSMGtfYpc+bQgm1QChbsC0xaYMwkDgwQ//VqQPjZrAag6YUb
rXkqSqurXrDBAbbEBlmRwtbFCxSe6bwB2nWV1QpcBQ9zArSYvQSm/0xJdn5EGoFY4NnIo+17RlQw
PysfdBodPCE3XW4k5udBiAqdDLByICarDqCeYv+Vt7p8x3qo0j4AKjXVOipCLILh+3JovXmpiJbq
bfKBtFm/UsRsGXRS76TuMd4xVE/kXQMGouXH6MWxh9LWbBZmYhoeAQoX5YkkUqJMj7SjNf0ZZtiI
Pw7Ws8ZEeQOOUonO8WbsNKyFsrCEndSaXVCz+zTK0f2oYqMYregJ4GCSTVq8SP4xFkzoLRQ2vyN8
0PWWTuftqG0dhQWQjXiMyObP2kyu41rbIOgJdSMp/294lM+qJXADIScH88JYAM9+h6AJ4V1i5sch
n1Mq6fMIyiK171X8txH6fZ3Pxxe9GxSl8jfmoKW0XC1QmhYEwOQ5FQqGaWreRZVBl7InPwHdJAI1
w0kmTFtpEn15l2cRnyvDprW/DpBGe3IAUi85sWjgONyjTWYF77idtv/m/8gDopFEc9SkfTGgvMcH
nxKbQzm7xgcDAOASYG0AWxzvQa6XkeMxfBl8bqCG9v8yxhNJjbvQplBOHDfgh6uVY3lj+CuXhrU1
BZ1XvNkpwzeBJVf/sDRn1HaG52qo/GQrILTVxDpZV2WniHVa6iLxCO6ImKELYvdhboa7PZ6YcdtX
Snbw5Bo7Q4glicZHoiwkzCSxECJ9M9zCBN5XhwaKejYQZFrU7OQuoXfqtCTXzXWiMejscGJCr71j
f5BluQwq4otHmdZ16ASAh1Ot0Ve+3vj4AMoNO0EEhPIyw0BToMuiJEKrr3f0QeUSXgPcl4QQ3hKl
L8jSubqLQJFp/K0Mp/bvk9Nhh136HfeYCd7Xuk3tHjf55vAgMjes/6Ad64ABI2+rfdZ1nJQbnamo
QHTUUCFQnpVkS0igf7GwNqmEWbUKeazRil4QIhECDc91f6sEolBYmNDHXdNr3PWItZbtZpXk7Ac4
veJm6qngu4loKKiHNO/JLSicSmcDLEY4bePgWlZIc+7j8M7ODdI9E8mmxefP/DT+JFLCjvgtZATm
Nu9nhWtw3W2bdphSGyx3fHMF62qIsfCSNWJLaD/uIwE0vwZZa8w/9vVNDgk2zWRb2GHqbzsVAMb3
zSiQBYtrzX5qcm3lIbEYxZjzqwFPhgCTU6ojQXIWH3kPSK3hHZTIYHBS9zv9eu5ALkd4mGxXwza/
vCIaon+qx7gGIxAtJvw6P2rW+QAbAecOxetJ6415MSljGfK/KcQJGgeHH9p/zWVMTBW5EESwSsOs
TRPKfgfOnkPZ8bP44PFVXWqWfOx2FRECY5MbNowvLiFimlBN2gBMxFak8hJMZQuMfkTJGlO2F0ng
K45ylPYCm5OEXFCxcA9ldF/W35t9AbXigHktu4aOW6ywjAlfr00P80d73sW6+YPmZvqGRej73N9X
/ulUSyF2W9Deu/6hotn6FbxYLuM5+t0FNat46vdnSvqlRahCCOCl6wDi5tFFPNA6etseZubUfosp
P0x7bNB609iP/Mnn23Lex/mywpyW/i+3ltvJVwoViuChJ/z4vN3qBKW704Xk6M3whn3wSitkF3wD
bWbExnX1SRVJMe5fYDML/yt3XWqa9UG+u+xzGJZFsZAep3KM2QfbRhEqlthmv21xyAWdBlSifBCG
QDTpOSuPdFtfcMu3jzz7bAaYmEMk+qTFmtJqyHIi4HdV1O9OwWSmQ5zuakNrs9F5AOvHIJJWBETU
wU8S4UX0+d1NM8OUd3pzADDvpcTcOzR/HMEuXWuZPGeAHm/v4JaMz5WMsAoY3tv6cWSF774vtWHg
/Y5CGXm5+pBnkVPePbI8cHq7Y5XV6+wq32HsWWNSjgdQPzCX4ohY/vv20YvYMlFocxjwlH/Ef6E6
Jie/RY4ANV8mUgEHxgI+lw77oNjwGCDDVoElw4WyXSFSFronQccrBPuISvYWfXJ8qBVWotXa7fmQ
MDy9K5DjJKHHg+zhjGvW3ODEmv5N8IeGpQDDfcCIgZ706pDvY8NsV8qy5SJn5wa4/M/JL4zzLQOv
a8wNpgpYMk0fkO0+N4ajyLda8z2RCx3V8/cFSZ0Jc0K9JLtWPuf7KLgCBw9NauMrffgufgSXUJpb
HL3XW+piUsAbQXHcHqC6ARu3xBt3XNY3h88SZ7LDu21pEhRrxaIL5t14g8QDRBBYeUAiofCex6i+
3boFyJHEcwhGDAOfKhKzfF2ZsKr0OLtDeOnNL6KHkyCBh7ZR63mF51gicJd6EhCv6UG/BQbqaTrZ
BASKapYb6kBVxDDKI2JQAYl5CvPvHFlQHdIM/1D79iwx+vLf7FdkODR2Tm94OzBzE+dOBDMGRp55
ZIKISIr6ub9em1hfaUJ5yQjLmSoCEovzcTVLQkB2grhFvMq4RLXaFL5eVtMy7EwVFr/tPKJS435/
GpWlPQxp7yNpiV/gxUL8YeC/ly/1oMz6aOMyhrtEWx87R2VsFbK3d0AYT5Q3ZrosLX3qjy9lOwL8
zuKpr7vFfbRLXYFhLJGVjbi2mMTPIvrWv1j4tiodKPK04GnWtmVIpGdA1WGGSQ4V4YRJGosCmS/K
rz5HeXbOtdGfnwVOLUhzheDeg9p9R4l3xAyNWTpLjIQnzxPQ5v9VmriYPT6Xl41JBeND2HQUsL7u
lW0+oO1/yiDw1AWoqLKt0UuqgOjTAZSXcjOTIcnvz64yJrAhApbtobOSSBOqidTwAIsCQD3GunrV
lueq4arJSsiQMtD+D+RHEIG+Oy7cVdnvNIgEqKbn8dDavgitPuWIUDlPZtnvZZf0UNwxUAaPcv3T
cU5degRnNpgDo0Mu8MZVNQ/KxI/2aVPllRuBVX8qRBKfRaNtNhPCsMnB9MUue8U6tPDT0dEf6mRR
7bac04BePh6TZqHqgFmlu9wQ9DzY7uW+MRVTkekD79NEXCuCqKpkEjtzPGSM8LUCtktszF/MiIyn
a0Z2ZTxO+1wU+mmrL8OaGmhgIlU6Nk6j3F+ql1xWC8Qn63gymkjcU+lpHRoVhprYvk1pWpY8aP4X
KdHhkMHxzBymXDZJnxZrKrPrknHrpjxfyFly4p2+Dse3aNJ9rhjHpNOhpWjuO4x1Sa1UJtDvk9DE
Ns+R18OI6Xs6WEJn8XllAV20i1ctIAlO6LDcKC82Gy1c82lDnIl0PXXAaHm4Qc3XzoJW865IZtei
6HM/tUy5+QbQW0C/HwyxPN5VHO1v3wD6+VsqfjzcHr7lTJ/dRSYaWdbTzeDAv1Y06iWVvtxyn4ap
ALwrmuq+1/8k86sY/QEp9wu0NHyUFlhW5B/IpPWzOxVz8o+BO/oox9Hvc6yGVYRTxtLFgFDr4tbK
IHxS8d07sKFeG3Y6/xH2oKAqCGmewV1/OEsb36f9njYwR8ERcU7RbKmGxgw+sQCW1gQYRsuqxjuC
aPDkUEMcNRZzZPkTwDeAOr14ijzj1TPXCt/A+bgSWs9Rtak+geYCX5jOLEWVRQ+obmOjS+vMA4ak
Aq1ydvcdKCAr9m/M5QCVUDm3w4pumq6jPHOpdYanw8uU/SAYwiOKJVR1TyugEV0B/loFrR9COt09
rn9RPiAQ0ENOXtlQml9q5e6sGblZB2Mjk/5LGhCZpkBgdjabiMVJeTuKHTFElGZkpHcDAbr+kjqk
ljlrFjttJimNRsmtsxbnzKM9C48O0Izzm5GL115z+FxKZmeQhyMOV3w1/a+Q5I1F9IIuO8+6W7mb
u+bJR4KktsA2DbZzgu/LDlANUM0l30z2mtX4e1p4iRl/o3cNpkAVJzreF/2xOCXv2Z7HVJQ6ke07
QtW1etpW9d3sQJP7YbJ2PTt5JDgMoZ95wdkgwVs38LfRCpQPjRFJKuRV8XWJ2NGNb6SdIDgLwW/S
f1xzBJZuoBNT2hXF++8aUCzggyTqpjfUz0jKeUvAjNC/VPUZS5axy4rxcdQwC/8++cZlAmbP1i8K
bKoTxofjGlSG8DHTUltzvWJIdx8nrSW7Tp8/G+lHUvAnX1gH2geV1fKl1bQr4FyEUdi6RshdHhM/
/5WKzSeAqTXKQMbqEy50H+zj6diva6Zyq2Q83culihvdmXY0APqhbMYVFOFNh5bR/i5INgrqt+aE
UWMyxOLQc9qkhBKDyX2fHrEl9bPanVuWDI6TdbIi8xy22jPphvtHe8gKej/hTxGeD0+CVjwHP76o
Z2rUCXvveTlRu6k0AmHFZ+xEej/J4QBpWKBicuxfJiYKV8b2QEq1s2HpEaj0oR0lg2zHtrwnQ5/y
Vqyzu/UC0C7P3afzmq7TryDSI31Cph3iQgBA7ianYopF2mrbiyuRqhLw248mPhZU716GVBhfE8PL
Ra4iuppXT6JDdOyaLY8Y3xM6SGfp+J2o3tV5Xzng3FeLeFsomRm1ISwnmYCDlYRnebcGQJ8VfsCZ
nH/BiqgMVAvpiXcgZ8ovvH+lQwwRZni9ButmoXy3JKnlRi98VvGZCiUNJ8RPRuXyxYeAOkTIp7o9
vsXhr4Iy0WeiOQ+ieTp1wRbSt+v3QQtCqfBPaGZ0c4RRfnw1unOX2EDtpRVQMTNfneryH6WXbfnD
67dG6wgg/6hlD1y40bpauchm6eYvHtDTROP5vkLbI0MK9BqWq5n54Gwm0lC4dgW5xF4kygOIqZzi
SwPI4RxJRAfWx3omP9OrFXAKuobVqWT4MzToGDRHh96j8DHVVobYvbBC+pgOFrUyOzDUo5tEEpp1
Jv99Yv0TX5X67MH5llx57xW/C4tP5cqf5N6xB65kzb5CJNIaj7+yvF6vxBSV0e77FLq6d2zpqS2n
6yCNajW+3HlBway9VETDqaOehcDWCzuBzGyPAQYveS9P1qN1T6s4sO2I9/yLHB82AgL8OKlz7Up8
nwdatdiMvpL3jQyfadJSX1/M7TEX+ba4lS98Ida7NWm8aSev+MZFkT5W8fAu4Ci96ChE0FLz5OfU
7uMgx5XfkN0oEGxYXahxMGXMpt8D6FO3/ER1CcpifOt7sdaCQi/Oi/RfxFZ0vdXAx+2BpxIPVkWs
6r1NSL2wuG3IY1Xe5UOKKaLus0nrcu8dfgSuxr7oe+Zqdut8Ent9i4T+HeMTD/oZGFNtI8ILtchx
tCxWk6pta/nRrFcVwfs26aq7YzhKY5Bj5HX/wQV9SH2I6rpTqYk3GkccXeAdBSNc8/G+aIg1XFu9
2LxEwD74wGg2Ud0rB52gCN9Nd5ql/u2zGxZN07fIt8xsP+CaqJJxrOWrhOZfBRwp8nexGUK3ll5D
GUzcyhkyubMOn+8+8dM5i3xDT/gLttPEISfi0tZCzJfYcgTSi4ggVtVFERmaiIq3hnFZyVULO31e
cbcxM8NskJjPsNaAe+AIjf9Tlb7LN34dQXbLIjVBZleP6fVkibacU58v1gF0tA/H5ZA0DEDoOKZn
y/4IXuDi+HoOeOBEktbn0P2hBQnFHZ635a/5nu1zbt4HaoO8SDfRdo9db+U6gL7CCAvVtYpBlP7W
xL0pNrwz+HZhVorcx4HbSwyhzCGzEh+eFiGjWZOxlL6ubUPQLInFN1N3rZo+FD3mnN9goKywK78J
xh7Su1tk641yzi/YOWbpbOTiquNUvc/59vP/QTAI4mq+tbqH3QpIVXP1UHmTLHVuWU4WZhwKh9fW
rEtOfMttaf9N4DFrMcJ8LLLvQZdwfHihpRQ59ryu/l2J1sAMyjT9tblNP4btgZy5PAjFg27Fp2RO
vAje4hMecl9oAgVII5GD/ARXptIcna4yNtFTleEuAjbghK2xWv5iWc63dqs/5aymAKxdESSr+d6x
WBNdc83jUY99IiE+v7pDqv/mJ0wPb+WK/hiI4F+hwu0tIvIZidvicdAlUYCWpxiL8zHNZJyjRuXc
8s9KpR7kKKVgg9w+UMReyEvkjqIi88qX4JhBdCsOWa4dxYcyWY0no/PagGk15Ks+3O3YE6agNLFh
L4+45Q8eNNXGds/yQDb1jTpmih60l3zTisAYqCLxKFA89OcQfkpy4peliGairPtzh8paOHO6GMH1
ciJXa1g3tjvEThQXytYPZiyKoiV4qvCfMoqX/3qnQMhEvdgEAtEDHnDl68T8WVPWNnnkTip2Q8M8
AEsw3RbDsCYuZYueeb0F5G4/2veAbwj6jfQckeHcUmO9lcOQ3bzUbDSJ8IXUb6T6cpskshv5g3hu
WB2xcP2t6m7Hc2+1ZnwLbsKRU1jo72KOeNhQr+sBrWldwljfUo901e958QZ5fP/qZkU7UiJeR4WY
jb+Gy6SfMewhHsQ48YBZ4AKJ5qdLnX3Kd5v4Jrl+ahrxnjzcNip+wmpAXRoPGGYU9kOtd3XJVR8S
uVHRzNFTjbiEvbGTDk1hzZbRKpTITpyd3QL+4VqReIUacOnMxD52VsytQCmJtOUo8QvPzVQuwitM
LpK1uaFBt05WR3mhEQFUvrPgyWYJgzuq2Me7ONNHr/CMGUBTlXP4yWEUrmBMcl5XSCFo4+CwDCnY
MLnQf4upLAoKBKlwz1xo9TSskhwjFwgrX5omSxnerOAzjevDQnGOx1xilqBaGQRam3u/Ora2myRg
peKgGJH62NfLXSZ8nRWBJLvI/m2qqbUfhUS+W2zUPvxQ6L7y9p+NftcB/+UIP+KI/Hgtz4+tJX83
OJrYoxDqxi6JpWuF+YZjwmPj7le0vKME92KAiVJTyJoqPmPuy69tuqBlI2pvOxTsphzEewZRPT4/
44HYzrwM49cgwagNwdX1hFhELOzXoawvKaZIoIZ+cbhsjZWbLzujtErIp1bOmaxBEpuBg46fEhg2
fT8ZKiz5oXNmLaTdz5SOV0pxuDjPcTLchEHja20CEyFY0woA0WAjYuY5UraBYXm5gMeOanL99bAC
tSLJIJ+6+IqpF7RnLV4clBgChXCM4eh0nMX1aDXoqXfzhLeUm31qaGwnQLekECAUoSxYX1k4qnSu
QtbOxJNG30074Jj13Va1diFb6/xgJQh7YZWx40QQuQ1OuSi+b1fZP61YyqNTUGsW5dgv3Bg2eA1l
7pOsaqcHB2RPxOEte/CUFkuvgXQrAeJLUQv5y8AAUTTPgNHHCk+A7SqqL+ulb8sov+l7uoYQqzax
FkChobFPrAcfNneScg2ebmtiXwT1pYdz4WUFrCyM7Kgo5m+qJdljBnxydYGWgRZPEeaPLFjr+KgI
zxs8i19aoY9MHDknhDOa0a+QsNLyvvkU5iScSlh5Adc/khJ5vyJE+i3pAQqqCFfF8hk8NeCTQJox
LJwhR3N1E8kCw15xzoE9gTrMksfGVnV3rmmHWoOZdFF7YAkEsxhbIGYxLLIXp2TZi9hirqdHoz0B
PWf9oCUJNYWyD1L9YgTIJZlaUfusPWVHrwgyTn4hvWdmPDcgfvS+4DDLTjj0pNp5KYBMWPNuTkxT
O/3aI234GMUIewaj9Q9z4MaJAYDaf/D5RTX2BloKz/OKunUYKoa7pyFGR0U3lqpJnUB94DnNxWOx
nwlVuL6f78/joYlUaF2Us++SxRji/NSzpfW5rJ+8UcfcRgX+5YhbRwfutMIVAuUAwZqRgQVGc4TY
stvW1m+SVsC9tD4jHe7H08ZHtTuj5MBrDHZTHZSofm+HCMbBrVXnNLJC+JWoVbOKfvXVN0k5KuHy
LLAfzhGqW9kCfXqwYflLdiR0pxbmPrUZ3i6DfixVKDtISHKmJjcGOuW4BbrEb5lO9pcpmaG8nwRN
Ww0DKVTX93N9KqzLos/2Adsg9A8cusqmuV+lggE7+p96SfXalOohcj+PW+2aJyjkmoOXQm3Qo0Ea
ZeohkgCaSO391T+AHZUPGOcncd47iBVb0RMHgoVBeplh7CEH11FsL9HGoO9y90Kz1SnhmXKyDDZ8
BOJumZSw7x5Q1TGs8VQU0FiOm0wnL417CF5KdiNCnQ7Z1RROyFV8O7cIs7AYVveKbmuafZ91up1W
KpAGz8rMBXtZKHnEatDmIIAxDSvWPNqEdW2Fpmu40RQyBgOshT898dybogd0AV5HbeOUyY74WjHo
KdKuHdVvsfcD/jTSQbucNtoeVH/h0DJZBJSJ6prjje3eRAFq3mrbGbUSrWOgYiZ28B/kGWV9xX80
0UAZ49DiA3vabJ45iiFRAEvx/1ukvCKtc/uaTY7b4MSLZ9JwTeCus+Z2HbJWpvqukdX/21rIyD08
CPsm1Z/mONOi0gsiAB1QKTHbNwpOHiIfzsKMPZyjKpYrfgv8JJk7ca6ehBdf7u74MHRgdVuC7AIY
e+ODzjBh1xXEuMAIvc3d/XHPhdirAvmU7acuyHbXW+g+N8KJrE5oxtQeSdkjwP+YVLB95PZSPgxX
XNx+8i1zFwn8HloPoXElJz7EKt207ZMyJ2UQskkFcYMnejVVUfHgFXQ2kMQ3qvskcAW8j/ikx8Wz
gwO7ma2anCkuB1zsLwy7q2/MP2XqIlaDHkxri0MKTRDcvJXeU4BMYbX8E5m+sODKXxypzNGK3ELr
vOFTmObDexYjh7Q3LITEmBZ6HidCxeSIzJ6eGWYsXk3bkByLQJZDGWtdqIMcsOXZEtjo4etNzmb8
AZoU6n3L1pl4df+ZYDYiqy2/6ORh7V85Dmy0PaPjx6bcVK/racWapl6z+E7UBBN1qXXJ5OtoGmaG
/xmlEmGlYcQW/XwXDSdyZXXOEXas9S4nOlmFPrbEFB+VRt6RCBoaSTy8/MXZlBT9x8Ud8Ntirype
4TCgk19D7gR2/gSwvj26XHGJOg2Xvi1BVB6zPqrbPB3xTQvqaDex7WJW5i6Y/73kD7F+94plILa/
VFYGH69XSu5kdfjlNcjFQPb5IuWKIzoriQJrXtkpHzKfkkIQtnPPbDaabbFG/HfQ1RCYPNOnbHQV
6kQtVJNP/Wc0rFNo7xbVlr4J/p4oN2XxbROTiKOQDqYYYeCf3RUqlHS4CTlr1xbV5UUQBi94b3Iv
QZ+77ir4JZzOFTCkDm4Xvckng56+P5vJUfXU23d0A2JRyZl3Wpc3VF69VqOkocvFrfe9fdmUKiOL
QAKg6/jGVKVUWGIA98e4xqFoARzVsymMQxoRSXifsyf1rt6L6FE6Mhl0BXmFGshS/y5e7f0PoTTv
jeJx7gjKnkBSNG0E///BKtd1LYT36apVYctsb+rkpuDfh4yKCqYmZAJmyKLPpEeNLLf4nnVPIilr
v3JGGc7uLO0FMkawI9njXUe+63B8wwD+0cKPMk9xxS1WeuLshcdoFb1XA21eZ8gdU2xmcFItavTg
K8f/EO8/LkjQniOL/06g8S4XPx4NZ/0PoGpePKfob3Pmbjf7qr6z95cHQKElSy+xxIC064c2O6vF
cD3K4nYVc2ASAguDF6ZwGL3YV/x0EFiAQfyEUwl9CY33LCwEeVI16MxRj4vNYzJF2iXTlO3PEkjh
3aOfDa/hVuJhACZEzhxBKhf/plV3SAfdIXw4jSdO9KKKuwZ9io42/PJPqQf5g7UB4oZfDWy/Gucx
WcEuqisfvqTQQ7qW8gCxyWzMIHrJlryr6qDkd5Dy2xWQXdHGFJZ79uSPlTOe+MZOFZE2P3MgFTCd
3xqkwnf4o6JYf/ZlEi54v6iH8ReV/dMpTEcjFPtFedUjRq97LHZ+3lB5Hbq877Rfre2h6jxkOrt8
9TmqkzHW6ccuh6eQGCJ951fAAGHq0obOND5O4tBOdFZ66UfEyU5gNVxJmY1M5Cne4CFa9b7JiLz5
aZXIYOxieK2i7vJkC6cbX3IFTIcpaPJoVCpFeh2znK+nechemq2zuwVsbtKHz/btviFMiwSIWoxj
lX296RkiU/rzfub9X65J9JdfZT3ExRNBvws6M4UuH88N8Xi++T05BQvroSUe2b+Ia9PmHKrxlmSx
DQh63RGvsQXcfvPacGN9kQh92SwvpFLNfhIhdnI786VVsgIlDuEO0z66EQyI22BZjiX7KhO2mMXK
O0uP7EnSyL34b1zjL2dJjelt/Tg1V29Wd7IRJSeQ6zlTbTVsya8kmgP1OatikDITMr3thkUcAKrU
r+T0JvE2AuKPxErH+14pFe4ZAl38QNg9syepxd8iKgMU2GKon2iHLRb+gOWC43fRkyYWx1xTEi9x
z6Tzkge1hnZTQjTwyEcnEUycUwNMgzXT004AyHnOdmOZk3/Bfleq9Zc+8+dtEO4BrVcnv6bFSYEc
OTryu20DYwiCAdbD3QW/2ouk3MxG/XDyC2CJ5bU3dOdmwt8wxcc9dsRPPbaXsqkAl267ze+66O5L
qAZJ/4h5/Y8lfozRteIPKL4ME7+y6KZ/G4kniVEkSuYeKCPH1TVq7fvi/lUYagab9+vU1ghpeNtx
OKOryHJFwV/yM/8a1eKBMKxuIBuNy7M0csmzNI0nw5IOBOMBmYm2VN2H/RMVCUwLuZXzrl6uMiqI
mSr/tFnlJmfJQIOj4XOtSs1Jgk0+I1f4JnwR7XpKIbZQs4kfhcbfROtc/IQfpZamqe6RZnLE/xhQ
52blr55CXDbm8Nkf23PH8jHsTfzSpxdNo+r9qVPm5CSsC/CUqSSIcf1GN246isrELJeajQRjmLCq
YcusH5qg9Yi+ajzxQOLF3xpOTUs4RatGuWqzLTuv7sTTX0wt0MJH05Et5eKUL3pjOXGwVXURFLCt
UQwgx/KZaW40RR4O01DpC3cYiCIONRX/pNZ4RuQe5RUXPmM/UwsrzWKup4ofOP5iZ6oA2xcvw4FB
AUyEg1EmpCVgaF4b0Wjl5mINndJrNybi8uSQ4qO6L8JTQgAa9hq2Sukkg8jj1H2beq9kD58xyglA
bnilPRST5f5aA8Go/DgpJdgY5zaMW4Ckdrv+J2He30uMeUp2HuliOt37vnHMBDhfN4U0xoaCVtAP
hvnZB5KqKK6Gbn5XG91GWX2/bx+ma2j1MobIpO0AP8rUxJ1a94A0ehvHM21QeyH676uk1/0Ui0S0
xGEPgyR/op7gHRRPZmLHlZu0Ep8Oe2XrS7F39haGjsH8nAI13JVYStRl18KlXTWwOqkKBbeG2FoC
rMWeFb/L7shTfkhAoWTquqW7222s1VTHxiL5k6lpAvqCvb6GcKuH1YPGoYsCetZgvpdD2j3F0r31
mHCd2UGAiAKGDBRmeRl26MXFwl4U7+vWhaPOd76YiRts5K9rQHWWpSqXRiMg4IEnJVg/mZHJB/sf
OB3gPLZlG7ZTeDlE27XqyHT9DJ++vJPLixQ4YTSVfZMG+C58btpCyMesLbJSfbC3YN8xv+RrOWup
DXcYakfsK+fm0JxZp+k8fOcATn5G3jwIHH0IhlhN8XNs6B5OPkKJIDTcUaY6fyXpuueFVlm+9akm
MBVRkDqU2OzWnz3VzfO5kUHwMdkiY0PPilbMxQrxVWW3cNTsqtLKwws+gNEQom/zFMNdrax8FBtZ
VrtmpmzcFqA/b3amd2XbOOP/eagwAClM65dz3ADxN4RfCAUz5iJ2hiqTKYG6e8gx6lciALIjlEmX
fowxu+Db4UiNNyTswpwO6tK3qkIswfz0yd/2ZjBOjjZpWLTAoAZvUskNLBZQFyPo9RgfPa6h+v/j
mE5J4DyX3P++LU3tbrvhI/LWwCuoOfXMaVrCMs2MJSV0qlhXJDVw/MyPy7Eq9pmeO5x5kdtzWTUG
Yt5C85XXlgkDY+AUkHxXyFepJll7IBB6Qr9MbSSw+tEo+gtDeTTgvlK4/+fdy+xCyR64lfZyXONH
OENe2YyRNyHc0sR1AiqWBZW3q4+tv34zYKal0e6P83ZgU74PfpmY3E7ib2FVymjseAkh7segAy/6
05jAYCJUnam2dtMox+xOZJQvY03f2BcFvPNRtlybWkjp8YfuB2X7wnAd8Qe1Z7j5FMxsQRzgJOlu
4Tf/gk+Tq+SIJbvyxCBy5YEoU6/wn4lG/qAaft9wJVFz5lxs/0HL07/sXvgjzrhjLuykrjllO78R
lq42Iy7MYKqV7NvUIiLumdMr4z3stLiP2mkVkgTa0TKdkvu2HqleD8t3HTM/4fGjU1QqxQKbn1ZB
WkMtfnFzCMhkiN39Ia2zvrRPw0679+dsrFYZZsL5eyWvWSovbItWc4qFJjVKim3O49n4xZRXNGnY
7KRtDbhFnIdFkoMLQHLzvq4UUgNo0vjW5IgD+a0FSG/ydgngj/aoEDJAwvmiF74Dct49iT2QYJGg
J1ZXHBn+pZVzakdwCHZjpOK4w3WphWRKwJI4W6rfiQOHX/LF1AkORPUBqYSDMvPsBEh16J54wXXo
m5x7F444iuV2TTs58R3pTuGpXlj4FvEpRGE6B+BZBmsficasBkEE5Ek6uHHx9+Jkr5G2i/LZsao5
nZgFkGZhbqHZEmOzv5JNvfjriVVXEMeqwzVc+pW9qQlCjdaywy/XLzfayjUicoRMHbFiTGLDg8IT
8UTCaRupJFxvORCxvL67gDShhuDqdcrn+x+untJ22insEjwKYZnPHzSgyP9NGzxA/MgwoUhkh2GI
VrSLJyPjXA+tu4krEq/9zbz1X8KkEooA77onE733m3/sQnLXpVUPJ7k76mV+xS0u2Heo6TacQimq
M1DlPlQcHodO/K732vr8QzCbWikC26Ln68oW/gIBCnm0Lp2/k9mqWkfpWvZrZ2pmIaGNPDll1C4a
I3Nk84K4DKVbQ2RnPcDCpGvedcnIQ4i1uzhEqkQllkrzB0/eVH0kiaphsvwAfdwhz8jfugmMKu+1
H7xUZ3Tw6igjCXCWGB5az/P6BBT899wcRwP9dbczYqh9rH+QCkqw9UoO7xTMzybNSqy3/VYlm7jj
/6qaa/jNsItcBYsbqI+cFurMQmuBuwmkx88DmVC6DxCmVzt7bbOu+Y3QW/2qPF2y3CbEuqkwP3uw
6iWLE2sDHMO9FwQSo1j8wNgwYdZKP1my1jgYDxusrO6MWWt1XgCdypPfRZfY06UhJpJTlsaqXnlD
m9i0MH1dEXMi0QGBPXI7DuuhRk/uN0f098eT2+QR+g43mJs03eD8rsEld6EP9+ckmrig+oMV2FG6
f5jIb7CpflIu7kEGfUGTVgBbDu/bJh4pvHuh7ZQfEMhXL0c9aKSNe7nBFvzN0hDUcAIm9xfK0gaB
G/8i6oHfSTzrWL70eDswXgyI2tp8tCnDjqyhhOhDoE+lFSI+VHAzRO/tlDm7L0msYH5NS4d57TwH
dVNWgLLVgAY/OPH/OSQAYVo+Sj72XmetX0x5nqoypdQW3JHLW9wDFCfD/YL4g/fPiBASiVhu9S3Y
V3f2sXrrbx/M3wO4PpFEkjxOYeJoFvj7vNCqwUWwih5QLtctW5aYAAOoIDoWp0orTsk9GhiVN0ia
DuOebPodsnZBBoa0Kp75oSYAW7rGPw6GAyM7GwyM9SodjkZqjtwAimXKX4WTdJedxsDhQfqHE5HM
HgI6/99aJsf7VYimgpiZK/aIy2ekwWrfF4vWslsjjaCEBpqz6GOnXFBAQ0WWqsSWlTMM41lNuNv7
kEpQ2amizOfrfMLAVcEjJF1AwBTHwfMPAxg37cKNteKNfzuoeKBNvFyJKxR4qm5IS+fjk2t34H77
w2ylwS6x7G53U/uhI8J3c/C4sxPYy838gWfkeo/3PFIp/lu7F33xmAmjDhIGkBtNDF+GFUHDlWpc
q5taMeDuw3i0iro39SVDzULbVW/tk/8ehX+02nJfbz+GN+Fz7q4OF8wmrEhA8d7LGD66B06UhEQQ
dPrkhZpcxutRvE6A3zYAau6WEn+YmBGI/eDi1ibcH7G0rmcVKXDEffJE3uRifoXWcz/0l/q9oPmg
SgcF0LavPs79NgGMzrHASVFL7yNf381XBwgWT5qL0R6uEk1W9tZLI2OGr1bsrRKJIyv/9pMMq3vX
uBRw6uDQEYq5NCif5tLx04pUh/XVzi6raFsMHtrb/MGUwoN8EMONVwYigEfEgqr344SNQZFagd+g
9dY/VpQYfKJ+QrRza7OTxmHX4hUGJOSIUVXRENtZBMb1G8/D2qSdkinuVONjf7M8s5OlbIvwZdwJ
mWibK4BxnY+5iCrhCrix+eOmGPUgwzM4nRQrzVzGskvpdE9UOKYb2zDzMrMGvaR0LuRVOxj4+yh5
ezR6JxUzDSbXB06xKbHgeEwif6sbMinyvuh8Y0RhknSdBWYakMVaFmBZnIf0h4upbdCtOigwRCdo
w808tYtmIK8XlZYrzKoifA/++oilLSffZdurO6cDW6dKx97SmxLk8iNrleCsC0uqUh7FJ/9P9nJm
oqzxWBIMmK/Sia/tPYWJMuImZS475actJCpMKoCVcv/pK3AJujA0CaLQM3F6vOf/sa770ZNwQSQj
JiN+EsX3wCD6kXjB8obqKi9n7hFGWk6GBrfNJnm1P4zMEEKQ54C06Ao58Nbkbhw73jYbkPTNO4Ud
7IGxLzo0EZc+Bb31EPwjmI0STuEyciwQLMWA4W2m+dXsGTrbBcRQtfmKBaECUJQXpoafP59xu4W9
JCv3taE5Ak0qHkiA8tTgUlUEL3UG4Uz72tVlsWcB8eGyagu/NAFAgiSn/NPiSUutuqRhGwSsglF4
xyFHmtOJrdjDkWOA6IMNkSqpITkumtsPBpYhPTP9OBWwh8fqSDl08ln/KYVmpbCB7Z/t9Ju+m3Gx
ePaJfNL0END4cKtd82HJ82LUyZ67HZFTya5gzGTnZvopKqO5RYE7QLBGizVWDtAL9i7vHWxFzmbf
GEIetXDaDeMVtS6KBEoagO5zz4wFOHr1bPWzZ1MJ9n3m2AYf6O1j5DeKJbq+z9AklaqOAh/Xd5s6
ufNx/+FgW85Rcg612wfmmfZpmp7JVBtPBbkabOV8sszZi2lwqcsrg1BcrLX9gy6NNYX9b1sAyzaM
liFW88PHf1qjGPPoI4Pr4o6pAk14SmTNfNvx2v/Y6bChWzMcUUsTCWqAAK6uPuDVh0bJb96pTgxZ
LTPkq4oAkvwXeue05abRYcR40bxYj+5UA8x1huVlmPjyNIAesvK1EzlDIaEXjI3ebbT974+55o5H
Ova3KO7+DHW1eywzLxfJtfhmP/fI8XoqePvWgMCGld0V9Dlzgsjl/HBw2IGDRvCaOzjgdEcTdpHg
I7jwwYEaE8nqe7T45j088EdPElJ2rNs0QTSzNny9WO/x1/+AxsXD7pXeDc7tsK8qH0oJETptsahi
ovZSnhYVoYPibxZ8kEYtTyNoELcwZGFyvP87rjFRXgs/z9tDEMsNFONIXompAQ8yWQWS6m6d4+ZQ
L/gXKLULguvAUSBWMDPxQzrtpW7r7VNqORj1kLudt5h0CDar6pwI9e4H+OApj/5ucU75vgasBxCw
jdAZ2XuchkuCEtu7KiKCRaulZq2+SaeAtUkA2i33E7pPyhb85JiG9S6+cobFpWKxugY0HeTulkJE
TPzv21/9aT1lwJetDQeThJ6hWAuy0T+U2YycPfrpWvE26QxMZNg29iFjT2lzlDBGnzWNLDJkwy5e
6gynlqmtdZBTjLzys7+bcD++cKNngWxC0VF58mujtQuFnl/wJKHdPo6we0hOKqTkef6ih+SDDyP+
PNnmgUqU9b646d2dlZnlSCRv1bJ3VrblyXXsWNk4e/2MOcMlELqcOFQ7tSpBzawnQ6G55ea27Dpa
Ba3jOCXPKNcAmefi94B2fYMbm6K3tsM6SMnv50sxgwwPN2axQzNOZcBAi/bZBrBcqWm84xk6+eHF
vzB4Pvbl+YlTcJ9+L8iXARy6xA0JVcR/Sken3nMOCOBiioG28JGJuh8CsXRuIdfQkt+XJhUYjuqM
oOYzcys6zFWvw4OcDXGYdsu9to2/Dm1J8OHBM7jqcQUVKDGMxGqwSPN+Mb/3Ce0P+/cTPsCtT3Bi
jLrPKNhXS+aK8lP7kwWq68H1JEwnwiOxPCKYd2msprIOsiQ2uJXOGkuF+2u5g4ONOLIVN6Ma9/wK
ea45DwZR7tPU4tzRLTucLmIL7Nt3xmjVZ/01lW2kD4dCL4J7hd/gZErFY5s01z0yVgNKUbRHNlQa
KqMeoPxQ5TAhY6w/r3ss8O4LrfEJ6/6SNXKWQlPTQSCXEoKVuWU3poJQhfo5T4oAuQfkg9BlKnzR
6P8La9ReDgvZFDqJFhJVKHD5ecZjHhokfYeM/szjdkjWfK2MrG2FVLzVIhfASWjrjO4AeMBUB2qn
8DDU0FitSAN/PAJJmrnvP8+NPpou9TIsfYMjsrAgOlMqa8qAJ6cfbJIf6qOES5IfOh0XhEViEAWL
jpaWPA0I92U2upH6fFdeD9CfjJuE6089h8vVa/oDVvZLQQpC7PNS9fjJaNh/fn99Wb02xxl3q9Qq
ZSCV2HZqM8tmZgBWnPwH4dHUWwshc8pdZimnx0IHaQv0Sy48Pf+IwEiqMHeGzV+xeaiGyvY0RIpE
KZaj6yhVccv8a99890DXFfJjT34YU5OpNrzDkYDMQoW0bq07UMjXkmLa0aAZqZ3E7VwqafRNxfbf
nHLWPxCtqQASq1PVNePhsLwFrL3VD+ut/2GtAsVFCg3S2cHtxbarEDKjTDyN46pjykX4VoqD3qE/
FVLt/829AqQgxsdkSo6XiOz+eyesaiLYxEVjJq7xvM11oj7xZIUt49iencoPzd/u+tEf3uHHaF9F
j3NaO+bMPArILC6PrPI/EsZ4XQj2pyVw0LpQMVQp6v4E/pLlag81gbF7ZMpVIcOcfGqosxN7VI9k
mEhmbF73HnFIDGLKKf33vTQi4Jb0XQ38C5Qji3fqW+rr21ino9vnK7kz5lUL+bIt/Mx+dd2TJT4S
G4AJ4b1MkYfJ9teUFD9vzuCHF2qL+fpFPA4S7pUASffCgDJhjwaS15g4eEj+aw5IxqkLJoKYqPUI
AK7nz62GJO0UadJHoePueTKnwk5TkdulUYp4mwcQ5rfwdP3larsxTzJtu3lx3qwv65UPlvW/cGsg
cCEdPhIN9RzrxVxBWE5KTkB5uA4fJh7gNn9e9aJd9As1IIlXK0eFhoWlmbT6T0IQ8ucoCl2ou52S
cCzmTx5zcs3Ww0y4fWl7N/qsR3jAb6KHRfLhhXDi1a9sgLT5zhyqJNhQFEllqnpPR3nHgQOszMEy
OwicoQj2Gi0Ou2+C6PqWwgF1JhXZnBLMH3D40nI4sLb9z6SRp1jqi8ZpOOc8J5YhGzWNLItsFB4h
9eYgvCqwtMLDNm7deqGTrJoH1o319f/TOEIpgZXJml4dcfzjEacmxQ27DCyVk8dGhCnB1N+hNtMq
JEGxf7ELAqB8XTfKaWrKkTSOWrm4JX0TRp4KqwX+G2E+ypODgGBUvf4dMMKE6TIGXUQY8x2D1Y/T
c3QwOCmV5D02bMLfFeyv4BxR0iIV1wGPe79UEy5QULw9ZWa7t6DdOuip55OqfTdkAOZDyBaBRb6Y
2ps0rCoQoKhFt9F6UavNLDbazGyfIBAb2sZRJszQeNqbmBYUQ5wXVEz81UdTN3NawZJzFC0PREkR
HUJy/rluMDBvRHHPRCsKL9gwR8/L/wbt2aLtVl6Q/DlzS9SEGZw3aD8/NplFUMb0wxVA2JTHjbCo
r6bDmmz0zvWnDOBOCV6UqnlkL/T/OJt2ps61LGAt5sY1Q89tAoQXLI2K8dxHzrjBvRbIcK08QYdp
49gbpfab+R0ZJRpu4/PszLIRgIFSw3ijAyvmq6R4zxb9twcbzl6OzkjAAh6OIcls+aRMHagwPs6z
UDakP6R/cDZqElHvEbr1qtHhkx37acGpqye6Z8kTR16oAslsNSdpjdTCXYfB1VpBRAlqOB1s2jps
cM8tzIASX3URdDcV96/bJ3ygu9Agi73+9OnKUOAozXsNVIKet/4+8FX9qSaT2RRDLXAw+L0jU4ps
EjbSzbGVhTPW1wKtC0IHPXmi57mECa/Jnn9Bm6DcV2yEqgMLFwea+iBsSNyfff8ZigSSwct0pjLd
HwKdPfPUm4vRRVkiFYe0DhETx9J2QkBeXr2aFJqxII5omPQ8A4vIjfmmpNxwUFSY8EZ12c5a8iSm
Sd+LEJJh7ClsnEqaiuHVuQj+oC+on8q/ITOzzsOjbqKBK04Tapm1Y9wk5capt43Os24Cj8E9ccYX
1PnFH9OC+MmBup/lyXgTrnDFMGZBh5qufVf6ffbBeVTPnwsicAkCCQSlL6wiXV1GnHPeSJsX8BqD
VtyGutOzWsWZWtiydwJLcFRWyJiLKPoe5lCNNRFVEPbzmUKq+ihk7jo+PcnP3P+2vUTtHPPT41et
9PL0LcTntMNgccv4xUCjpZONhVqL2mBYGhWON5RunvvPwL25nRZVzYvj4uM4XoXUxXsms93+LnSM
Pu2riSGnqap9SPqLonXAkMHgQ/qruT+N/GX3z8wLf4gzp470u4YLs/JouIC4Mg699N+xRDrnLuPD
ggYJiPqUIYIBCL3lYV5XPmS1X216JmcwY19F+Chf/zKNeprphDIymePoy8Sb1uoJV5/nzlo36mzT
Aea3qPSztMZtc74JRKUzjufZQSs0dfyVCIcUUzwheAqL+aLFKHrRpk7MQ7fMlWdGU8IdwzXuM6Hf
4jtLk5lObNBUY1WiE/KDIF2ohBbewaZNcbd8uVvUPxR0PWt2Ovb3Sl3KbACUdOpZZ6C37XIgWF3e
a0NzS1Xajq9z4H4DDG0AsU0gK7KQhPfu0JDjcNeZ1DpuUvqTr2CteLbmd/ceTDU7YjDKP8RMnIlY
x0D39URKots4qurAEvkLzFVEUa1SWJXERl9uztVBFQHzac7bT02E6iY7E5dfY6glIwq+gdgim1+s
YZpDXax1Na8AOPdnGSVWLTKcTJo/TX9ILW/w5U03k13CjSLrjmNIk3Qn79hZAQhzHHVKLYVZOu82
34iCzDxbOrFLNJtM+4kV52FFLBd2+djt4tx7I4OiccMcqx4vzPCLHfFWb+66sr3EZXiuLTAZnBy2
c9ql5b0QrYpYxObsRPQbmFaQboXzaqZKUfnQkluAtR4TxrPv3Qgue137AC+ZczmEcRkEKa1rOzLK
Yc0E2t9qFjkv1aJj7UZPpuZtPgdQaU6/bSAREd9BJji8GptJ/gYEIz+spoh8bjGspIuAmAkC0xRR
n2PYkterVNHvqlvTO4PUlhMFZoJHDAbN8MgTPN8iSshvU9di59yhpCdx2rOQwlD0azYx42JQbN50
Jh0ZnF2VlopfhXE0XZiJX2Y7uJQvDMb+iyyWVGOZm3uDlsZgNJqvMMIDHtL7WJQsDsUuq0lgQcUj
3IdBm5s05fMlNumFtNv2jskF8Qr7l857VWfrFh9u/ABaOS+zHLmkRoNBVylWWKP4pNPWhJ2NEkb6
RI7IOzxthborg0qPx79fTGDBP+gUUd8kC/v3RvG7S2Qx6H1z5Gq/hYOEKyiXqFKq4JTLrC4kPGYR
ZBYH0yrvMI3jzMUTIOU/y9FIRx4JO0Fp3W1e57mCKiZkEOTfGyCZ6IxDasvcOYl6OD/mVSOfY5pi
B4K2XRNbiIRfGJ/KmNQIfMDprwJ7CYi/LHqEBPifLzYwhWp8J6DBdZenTmaPgjeoBXLjjN7ClLK9
hvQL7w4mR5hvJxKE3Sif7YD2amm0/Tc13ajE4o6vYobMnwcVc6kh8zKl286dR+nAZ9sbWWad95O9
o4xI3XMoV3QALUzwqvGdWrrpevFCbxW+yiOMdrfM0YC+iOTU+v4i42ifNOAdfctxg/bTztg9h0Iv
s5IvGlYDgPMpQq0+JBjf4wgFONEjw2jC2bZNB1ldkLztBE+6db95fqF3uFgx+4BkDB9nVVfoUG2+
hmamSES7uI7Hhlnmov/ttOuc2oHapqTRx5+inKqtv+mfyDjwWw0UBVtWx7GNIHahhQO/GzL/UQ7h
IPubyAFgM5sTE9HhHGcNAQuRinqm6FSIyFu6vzGy+kaw1GHlO70I7wfNL7PQMn6/ay22iC0X3z3p
RvMBxzSC1Q9yvbnF4OCrQ8K/P/u5oMLkG39yvkcIGWJv/uwOjmLCO8u/7uMiZZeIsAa9o0VT/faF
yea4YlqTmdmXhquodXgSBUWYjhnvUjns+441SSp3zvCdKglSLN5FWvjlujgoeZIXbc2ISHcW8nGU
CVy43rzVIRMpyESo6+rW6aO1PPKtVGYE6wzNelmrvVUjM2WaUEN1pD2RRVT+OZxIWvSO0NiimVeQ
09uWglfqdTxJOk4EpB8lIPysxo8NFSf9sq+JbE6ROci1EtzZ6V/+gi427ydGO6yaYLXvFGNqzuoi
fV95psuHVFVkWOwIctMJ348axDk2PMUFCxckVW09wJ0fBwdadoKPLzdiZdoztrsdtiyyjp4w59YC
5t/C5txZmuH/deW4r6TY2eLjLb2H71G0wZRPAf1e6J7WwufRLI/p9RUdsUrsgVSDBT6UNqtlnXmI
sbFcsecFWrtHQcKhkWs11gZdjaFXvOp5VA2abnSohXNv1SFFuHQmXzI8MDrIvyySYoVo9xrgkp50
dZvSD/3c3TSyZw7IBLQWcv8d+sYu3FVS52wJupG4BA5I8ymaxDAe9/sDEB6nUIagz66a/Mc46dmu
O6MqTEdGn6BPuSDsLdnkVxM9Yh3UvQMAb3kQAJ7NHHX00LVZjtjY/+6A9jEoNF/mLXz/o5QRxlWJ
7MjsK/RICQbXlOrRkUmijYGd2rpesHkVFuC3SRYOuRGCtvLWM8ddPLFTNacwT06XQvNQbHwEBmzu
nSDgnOZjDWNMCOerKsBALLJqhxCRoMpRGpmoT4D//rVGcqob3KeXkMChRZNtuURPSN8SQ4yUSjuF
eM9VP0SlfTF9EI2y9BRaL96R+ouNOhpwPYB8IK9YXUSrq3iaj0fgvbQnHznN/xdkIRPYp8PRKL6C
bndfOqxqCw3oYGKasAuX39YZoFimAhYLWTxR/+VtnfOt7oTLa2g60LcDA+L+LD0uC2YOw4/abt4Q
ESXUwPPF8LE4Vc7IpkrAiWRD4oO9sVSD/YmTvZ7nMZuQOEftTVTQXVV3bRQFr/0wFd24OrTFvoPK
xJ/j6Chi22VYeFI8KVrcEgjaxjC3Ns3anyz+NxS+p2AvTUaZgnBJjzWvgDB2pgpJsAvoxaqpGg25
gTfL9v+9ZLHYTTsUnYEx8E8m3pgloFgLaV8lVjkdDP5w6wWPEljYDzjczThYQOFBem9UNMjKEk2p
fHc1PsO/wL1yTF8peyEcuICzXxYzC8rMNA0CH7QOkBi2UcI5SZ/A7ccJdRdkvh+W6yXMe+Xbgkbs
PmaNiBuo9IEDG89rlg0r82/zMaxPL3PUk979vLrrp0AMobviTMpbi+4ETIqKjEF8GmsuGO8cFPaC
vhnMazI6WcdCoaV8R2ujzrqt/eJgFAHH/yZywDJOKLGXz6cuuzer8dus3OpxcDpRaOoB0MumtMcO
qOigb6PXl8beYe3SEZQOdinFS+FF/ARrwavR+yUh7eLMamnOgg5b2V6V6sXyw/SZFgZDhbt1zDjj
/cG7iB9Mm452wEO/0c1gxunZHcZrPOq/DD8eCwCqN6iKZrEDBdYam2xjJ+DyU3nUHqJwYTjeaqvJ
F6tIbKzHSkdrzAHNOBC71LZ7bWN84ghAVAynEyIqvlpiQ+0pvK8Ru2UqJSysF6kg8QF7Mqwj0E5t
Xz+miXMe1psYp1t6AI1ggspkL/IVvlbXvxfFp5Ho5pBKaXTn/7mP5ORh69Cd0AJaYRmvgqNXfVag
uh+oh7lnCM0cB3hIJJ5XH8AZNzLOM3zCSIbZQceHzUjRIjlk2Bpri/oVtQ9T2WfC7mmMS0UGv0CA
BY0pqtBiKjTLgP1RdruQS/f0RcSW5+2C08dHT7TfZn98UEnGR+TOmgTcyt0egWPl9dnJxQisMOIf
Fx6LT7F0bLJ4hsUXhS6MTieQKxarsBBN4ergyKGIiywyuCornms8b9IyO4aue16/YsjZzAE6K5mF
Zh+khVF/04O7a6AJsJ3/E2vKixWOYNd5sVQnx2ceqUc4Xy6uW75eOy8I6/CZPbZ2p1BPXxU1FrWD
A2lstdG7gWOSQn86fBDX2JqvlJczfTmBWH/tcZclrJrZlMgtJ/chdGjRpLVFs0wV7FBGmsbNLAAk
sAs/pIWf++KsMCBB8sINdMfdT0igXhCNqc7LoirGiqRHTu7vPLQZawxoHtHKnTsKK2aWVa5dydie
aHrli22qsqVY3s7w9t6ogGqA4VCnQ8j35JgpU1O1QN9Ta4XzD/4HdDNKR/hzd9O44F/gL085pyic
N+ACTb3fB7400XLh+hY2/d9lEWf2iAVdvz3PJ0etRuesqWnJ3vF85Sgax/7701BFWxd1dKm1oeb+
inqnDyjEDcFEnxOSeysGiuDugOnI5pSWdyOC9v1skls5kQWZ0rTH/voMMeAMqzlnt56KkEj8baUs
ppPYi5orJWOMdfQ3lYAC5+iUlTm9O45l+0Zgnv4tgD0MbSblY7JoRir8MLzt+6JeKku76Aqe80sY
54X3x8Et1Mesg/qZWfl+GOPbw+rSgNlpeteVAguLhKoAFPN8IkCyL4d95hOhY8cy7ra5Z7JxkGrx
Hib1/75i+mOydxG4+86Kwhag/6YjehsddD2EMhcvgNoBTuFmTnxg/lDoA0fBOMsGveZHHdcrvZaa
qBmUzFkZuMqr6nI7sUIVXdi01qZMT6Pn9oiUyekKcuf6eybFIpdYqUBcDWQwFhIVNU4Soml9Jzqq
RGYuyCpwRSIpFeyvydmsqvHbts/M7KDwDT0aoJPhVjIpQPLvBVkdcKG2s9bWa1CL50IODU3D3KpH
CW1qaQGcshsaTauqj718M8gBproLqpyWc9tj516mFb5OYdZ2qZBEeU7O8p6GJT1EnPTZrvjrVQy2
3vn9oXqEHL3TDG6D1lPUXNFM1HURSVjBaDjqQIVYyeGBCyIUT4mZt2LodCrK3UwzKYWYcG7yvMVt
K+tufzbLh4eViDz+LqlnpAFzny1Tb1MxcE9kNql8TT1KjgkUPmDgwnce2737d1AI2S0669sKSLcZ
EvYyByALTaThdO4Ur0vqPWHJ3rNAy1T3/fWICvYHvC1tCL2/z5P7tasTurU8Lsrc5GGNuRLOC2Sh
Kf2WS0+aM9DF4Xa7oONx+nXSjPqe5Nbb1E+mt98V+h9pU2GAoaVCaSfy3w/WACnnAIkn6SoqmAiE
qZ9xFAohYmHykooOUDYd1Gg/Cgu8yMS24Ly659qWaJLEDYjk/q6k4gfivA2Dsraferg2iehTgBTO
FiX8rRvj3ouXEz0E//cfwdCM6wrAveh0Y5fwkQAs+xZIBYRrj4qxVYPFPKvdAvei33YpFUu7E6Se
m08mEEdM75pu1NYUk6m6CEDGkLgMFUoZlYz2kzMfQNKuht+iT1R9cHJB1qDeOWv+m5X6SCbDWDfG
Wax+atzDwYPQqe3Q5SXM6NtOcVRzg5Ua4Lb1+kk1UZAOh9NKuiFrbLe//9qBZG/0f9fJYAvHJYdr
ls74gnpWQnglAn7yC0WsUBFOH7bonRbGkzGkVbBaMDUSWSu0f/fLdI/raRA+76EUBMRezfU/DARP
9v17ja7BlvCukSVAJn6HPSlmQ5TTpuHTU9n3wcxFz9MwNl29sfiwG195M/HUTBiva++sU8gr9C48
E6XDhGnscG6XGOTxZZZksv1jCmSpb0K6nfpZiCk0go6mGS+ayqAaMpZjc++3KqIptA0vIvT7PByk
cVP/FJDC0u708/rd3vEYXjzhyF9ChI08RtzAiwl86uaxnTOVpil7XvFjphzHgincldOqIKD9xDA+
8dgTSaS5r1Mp78QHuL7kaovPp6Z9s37pBYlHzyIzNhQuPBKeifYHsbd+wNjPNoJkMgtBOCQ54pJD
GsoI18EUMi12G4dAc8PzZu9A38EpKDacar5QWeX9V5LL9D8yXuxzN813ZNZqQtvttfDUxfBuxVYm
qiZzS79MIrnA95DA8LdPyvroL+oloyp/OTI16revsqp/mIYtqRy02FQ+MdOrLoRqkVomszKKtL2N
K7DOyjyXM3DjzdP0D1w4cFNp5PAX1+QwvfRl6oDjj5CrL9qq97zAEieWBjLldno34GVN5OwWR2WX
O2DZ3Vu6VgwWU8NEq74EqewNWVD3lI8+ERtsv+Al+y0piAYlW7mrJReeuNmAJeBdBDTpWgzQYJ9x
tLhxtiJV8tUI5fgGI1QEy1erfIFD45r1Ho7zXaTtFcCJgssPRH5zXmuGPTVjakB5Hr09dMIyvAw3
Io+Wm6Mg67JVVVc/4CY2KiGeOBxiLXDx7s+6944H+lAljdDwSA5MIHEN0YiuFNfLTWWqN+NMIX3+
DYqw82NxsP9COQ/5FFUFn7F8/aWKJ887UuLrF/kCaaHRMUFWz/hmPxZWEVwmi5tO3PsyR4dpgSDd
74Mx7hjRYYc4w2gxDIhl7CmjmnyfGk2BTciWN1hn1KNqdnELpnF00bmB/y9hN02+04l15iNrA+NF
HrHwtgue9kzkp+tsfbZS5i6LajTNX2vK34tg3FlidZ36W3nVFT9PiwYSpg0edHH8CPGvI2FR/nKH
zotq1PbfMTRO3xHekc2yJzL+j8hINeaNK+tglAzjT3RPHfoC/HXmWWWQa9IuNAXMgmCSkDl88EzE
tZ8U4vbDjN4/tN3zMKfY4nTnIB5ht//lldfqHojh25SngOmfKUEQESQDluTx80GI1zoSEOOWc74q
swCFHXnP5GxQlKDRI5hiybbvhyNu0RWQeuX++vwn5t0JWyfSWl57s+14kWf46boUy1If4ja8Syqt
4kMzLVmQp8n7mT8ahWzPMKrr/QbngoPRCwTOg3uy/12YP/MbPR8k5L7qnS//ChAU/wovVA2AChbs
ATMYE37g+qy9ZTg2nQXazYo91dRJIMb8zCLAM86GDr3szT64Ai+BMc4bQqxQF3Ub1tBG/8voGms5
vMw/5VcUNS/ZjWYJvKJpBt/6Vl0JOFOiI/qg5TCnsCMD+V4FahmPpAnRCowsNxHBJqlvbKeSm0PT
Bwp/sPHFgQh+dzkWvLX1k7Me5v3oTMbj8wkxHn2IkaVoSFzS/ajWE2qynlf6EXqb5kIR0i+gSQGD
HWgk2p9OVi3L0KP95OshJkUS1Fde/GvIbkGdOsiZYtjUc+YYcexbK6q1eMa2MyhPSJPvYFgl8YGR
looiIV6ow6dOUkPLAWPrJukFOnKUZWqWt2sYhrUCQvWLR5vIPYQkeRq0I4Qd8ncyAoD+ch0KC0SS
+AtNKw8c0IH0qlntUyx8Y3YjpYyuFNrkOr5cxXNMQgT9ThsIEk86HLMWrzyeez017N05CmhQOrgp
dl3MPek/AAjfvmAsa/mi1f9+gonytWnZ2T4xfwYgOaRbBnlJlJMIuGOehwVCaH48T54XyGf6Xmpl
KFGrWEZW2Om/u+KWyaILHeDeRHR8HM26d+FD9So5lcRpi2Whp/LXDSjRzUAl6BxtHhfrU8r6M7Rz
+nL9FXtMgxPA28SVrVnxDaOEhCRTXtr15hJtSADdms1W+K66wSJLAcX10yZH69YhGtWPhYTR8CwO
aA6FoC0r1+gvjRmnrSC95yxrepXP3UUm6pGT4MlArSiQgBjXZCb0ELEwEuz58pFnwIC2cRZK+G2T
8W0VgrbaJilaJE+h7kpHumamPanAkgI/a+rEXJe473ztodqEcvRD9pfm1ryruIKpPQOyX8uVezAd
WkbG+8KRmbSC32DyUQERxGcu1kdsK//c0vbe6oJlU7oUiosBzBUBQf5sZZ3HZOwlj5zhPVhaVWZ5
3DLO/k1GxBnzzi3u7LeQ/1rf7ycNTk/c6StSBrDs7MLH8YSB4J2QkM9/wOFLX1sv8GiAOJjH4f68
SKBdy9rD9vxOTrVb4W3gJISM/P+lqjVZra0A4BTlxC1oTjs2QMHQJ9j722zDeHg3M9QUbsvSdrDm
fBrShssqAMYkwsp18CTx9oD1wifS3yXhl04D5mL/ELLwHoJLLVSDQeGNvm3yfOctRTEmgafUh9Wf
Csw2ABwJAy4NgI6OxDtPNO0EhIIF7uitaGasK54c0Zv/6xSwYv1YG4K3rSTLuspp/vOYmZKzbKyk
IgkLZJmzkV2nO8Q1q8mqaEhe2++KnJswWBd6NZYsNk88yC06Gtlg8oDzig2YsCYFf2ZvKp8CJDDx
L7GkZ3sWJ2wX7IuJRNCbu11kEYqd5d4todNQfJIZXiN5il3m/aGqc++Ri/A/DcJTaj+CDClB/1+u
GyzvxyE4LzhgUC7tVgdEdQDjE+COXAnFO0x1gBn4jCv5KtQuMIeQG2kth1hm+xF2UWTug//Ob3lM
HsP1GQjGeXk8euo4/WU+rk1ZVnwf+9nNuTGnOYNRr13fwBWNZp1X1axk6PKdqd0HrTdMkDH4gqp9
9Gf8rtowB0SRLiN4Pe/x+2KeIR6aaWA1CEMw5SCBlbVVHtW2BYKSkb4GXKnxfospOgmvUe0oMqGP
uQX+1Q+JqJoXgkUZ1BQcOVACpsYDGYtFr5d1RISJm8WA+T3X5EEWB8MT4PkI1wOr6OaPfeJHDDs5
9bT3r+RORZ6l+9VggOWNt0HT4gSKv9Vhits7R62iSzz3o6iRJK/3c258WQgBmFSQ1eHfJIHkZXXw
JxTlf2Md4T9Rb0yvHzXvW3sHHtZQ4sDyQZUuvBoleq9DuC6ra4q1O5g6WEiUmuDqEHdXtdpTdg7R
mtnbMKwaztOoMig7tHl+CWaLBk1zMDa6yxMb6ZLkzRYeVNMsaSMHNmfPPIs9N2uO1EIPj/FYh07C
fVe3iOd8IXYEWPWLIiIGh96sTHKxNbWm1msA04NDW84It+PgaK5R67k8k6LZST3zUpjZ8S0phFYK
Ts2qL4XGJfm0qrULUiLxDU4rXKMeGtmC4c/PSWvF/KZHs1saaXh9Q0D7lBfdu6AQB26waxHM9+/e
OfbvUo7yn8r6PqCbW/H85sYgJiAEkCG+B3YWp4zWxkLTw2X5IRX3pgWDQn65/uwXuiUxvDWEYr02
jHO5d/E52NB1ABL0Ne2EO1807uPe51PAjI3v3chiW6S8M9pqp3TPD72HNRyhwzDZdOqT+2C2zlji
BixsnLoAFk0dBvd+GpCM7rKv6YvWWqu7R8WHMGkO5sPPDmQbNwncklPo2755360PmHdijWlcQzCw
sdSDKD1zeoBzJfSfqMOjUjOHicemIqV/L0ad+OaqMfZOFbAR+qM4fsToQvYLT7lZ3DBLA6UzvQ/M
bA3vRbb5WR0f4bJG5hswBToH1XysCdDHaePnX+WZdR0roDCruB+thAs4u0aq+vIdhMPAzcY2LJQb
mnmYJ4qXukmyYhO3zhWcATxQJM+5wg/C3KKslh1hgMSJDzfE73Gns4bfCW9B3/NC6X28+6zaBPg8
7pG7B23SoCvkhFbB9LMcpCzIHVSRmNEu6TzNYlg5L0HQ6RAqsesA0gZAp83se7U1LPhL/7nq0Heb
BohejK7yk8NY4kRt8sbznzEKGGNZCsFvKji/W+mThkVcF7ouEVOA+PUZUwhYHEGyGS/QTF0klzQN
WXoVmgJmpTCDwMRWM+my2uaDCAFf6Jbhek8S8m7Gtd+yWREEpwW6cvj3Ze+kUcp4wTLppkqIsRdI
S/kqnsmS5IWVPjx2/r+LINIB/snzOADtONJKpe91g9rgNJR/EQ+rwR+O1wD0sYbRz28MGpTxS4Xe
XXyXCyqOOX7znBSzO8iei40YN0plRy9blEJKnfLshE3ruKwIWssCDosvCEhMvxQDKgM73+8exW8J
yON6VvJpbLb16laAT9ULwCY//3ghV5wSEw1SWMBK3oYJzKaffv2BaHW1/9z9dnEZlQv0v+XkUIhh
NL0VdnO5HybbDfHNpgCmsfQFDiiPYsHmBn1p9oliB6du02RRWZsma+INI05VHupQXpLPO1oBLLXi
5Q+r+QhKTmZngwraKpVYyTwLS97upsFVNgo8onHfoIad0zJeRgMh7dxblfpEJ0cE8KA1dIwCcyeL
rJv1+70/74r5RsXSismPZZrM537acuQuqb3+kyYA0CMWP9DSYw/pt/QVLVp8/0xUzM8ZZE/ECqMW
o/mCB+Mw2EyUFojHP+c/OGrCrAdFd9LS0q0+t7W7oxQvb3utNugxvKAwdX+8mw6rs7rHD2xxM9YG
FeSQnZqbIMSBsBFZp9lf7sSFLNNCUShGI0Bp0ePx21GCBHK1U4LS/bXK7UVj1x4abo9VH4xCMPTV
lqRhAFFgL2WRWDizYIxyibcsRLxi+DKW6XB53Cz5iSMjS9C09Ovdemfe8ixhq9DRxwlmjHzqaHKW
4qqfvhfKqUeravdgHN2bRt/DW3gZ9gptwkLk+uHIK8XsqRfBB+vB1Zx3UHpju16DRVGQv0V6AaDR
gEltbrxrYvkdjW7QH33bswMgoNgqGW8aWZSfRFSICBpt7xEw4BRnaaKN2TS5+SWCBmWy1u4o38y4
zSZgIn0ZdT7lgL0wD7JEOlTahV//bXtX9AI4C9wJboJ5oijjpZquRDg5MjHdphuAyOp5583JpnpR
P5qxqnDD+5irmiwv7E1sVv8oRozEGKg/Ttln+f9zuPxb1+Mi9zm6vp4O87dGervNrGRPYSYzfrL5
fRyz4uqt9UEuzt9Gv30QBTTx6/oFPSE1UIahdxWSznq9xpQY2/WLKxRahRMmJ2QzAer2yOCqF+4a
g/4XWuLMMe96kjcJ+kmyeXvfEvoJT7oqJR5msTUVKy7PDzhJUUTquBkEusiRe+RrzX0cnQpaJLcQ
OzAnD8WS8yq5m7u5SHof2UmaRw8a0rBRGrrqN0MFHj1SxNaNjUgFZuh+2ib4kzZYa16SdJWTXzNf
HpxWZCdCNm07ymL/eUq8YyQU9BAlE7w1iGatVBqe/Fp8eY7Hd5mJoqMoi7lzBhPbj7z12IOsFnrZ
Ul0y8bZhhwyNjtuDfYj1PE7y1i0p/9EpKpTsWVfL9jqc6oeXQczxaxvxcVtG5GNuU5GSYPxEUiUw
L0oO8/KdrSqUUK7ip+c1GqsenX+HWQMIwo5tsmu5QXTkPQ57kg5F+r7C8kP0o+X+iaos86C8E59b
s9En1xdRZnf3Ns6j3C0qU+3w/zSHb0QGADE7q4K6IHR7+i7zNf6CVF3S8ttH03XYfkxJmT2Ya0ga
wFmLlqkotGXqOY2ww9Ke3OXRX6FKvBNEBLb8/0KlaVqcxF2d6UcgHEfNbn3pHD1blm9om6MySE8Y
LbKKSXHEFldaQJ8Ws/hV93I9hndCn3n4KDdDEEWh1qaXdjLoC/GZZ8Kvsqiezi4zN4Dka7IY2wju
RmXL1OjsKIE2AwXOAbMc3NIo7rXdDqr/eJdYVUQRclLM/iY3yMLZGS4xL5/ZQHhlUuwKJdX4jCll
Kb7c+3FSGuOFsmcyh3XWz0Z6mz67yvS6IWycDXGSOlO3WZlxcEncFAKDMT7ctw3xC+WsVRxbSISl
UbZu4nTJA129KHGwmfmJVS1vWAAvGL9kFcB6gVnUGfgwi+UJ9xge/x71mNumV1rRoBglK4SbC2bh
4WYQ7l2FXefCNjCmN1/aBdpE8TKuiv9yh+3X2x6XZm5mBkzwVE2HFRnTBBQbTUf0eCxZHEhOTw7Q
pPHjSVijaZA1IgokePh2n6+jVNv6vsYLypzSTE6s64bIcLQjXWOXTayNCiKQ5Acu/urjALbJF78u
Y6QTqesd6UcU+isTOWkHcNKDxPYd7DzWbUfGKtr2g5LmgqQ0fnsdtkArrEIc6l+danSJn+yUVB3Y
m/bHJ1yEIA7YiWvtnCPXyW1Zn2EY+wMTG3yMmgD6yL4e0wP6wbA2tDjG1cy+5F2CsKIhfI/+8Nou
+vM8fRfn/8hkeqDYDc+PWkgOVTwJ6qiDrhzLylztt/3XuG451f4+++JuvWue8UOGMCHYO1pky36I
u/YYKMvWQNuQc9w5MD7xjdlDibWKUtFZRbzxCRYyDGUDrg9WJnOB3YGrDSYTEJoVs9E/5xEO5Q1P
kZp3CyYdD/CGyZLc87sdOVlWuISqp8Z7KS6rU+W9+S5TUNGHu+V41wrZEd4MImYU9Hmr5VLRBsKP
dad8AHMibWG6hxf4rA2ewWNocxXwcCBLyJBKipHzO+rFtrhk07Pe7p756D+b2FQJPcfIxcv5JK/4
R10C70JtMIxTKHekAvS/5EL/r8bkC1gGoD8ALodixpdH8+sOsRUkVq52TXnHIdazsdLbOQUpr7H9
fJNvccfJxpoXxIC/jaKuK2XvQJjXxm1UEeYGCh0JFxnAEso+DMn3O478LmpyPPEqjQBAzldNull9
GO6ywRXBb5aa7LJvGcbN8iolo1WJ2PF7tW63pPf6DgcenOJwDImSQG3OuHWyw/bw1GlhxBHDUiuc
hW4HpFj+zGEFPjjIz0hYc0jaCfTsqJZiLQtr0T6C44kbAkhx7y47X5LoIQ7or3J2ZYg7dkexrlmH
iL1DAQHNsDopcYKR3M8bJos7/9nuyeDLMzSPpZI0k+iLC/mKclm+xN/fDYpwJa1YDsJNEyZXc+XR
CZc3FqycvznSa78G7dMu0PgeUtPqN1H4raB3NqfWvkZlZgMJca+trK74r+A74j9VeWEm7SSAs4MT
nzzSnuwKUlrBVVyoGDmi8eMV7xjdWosL7PMp//tcAX5zxpx9mZBUxwP/0M7pnBIhFnXKGMC4Bowj
ICQbTxm/h28QZ9JrSvA1JtGsjdkb2eEpg4BRj4nFRmQtphPBesT4eXYn5+wgxKW/PC5wHP6Oijaz
QpmHpaXtrk1/r/GBWb24m51RVenltqnNpzm6A20dp3AtUwvaDCTlVyAcjuuL44fzfKNdjAyp4hxk
IMbo60spKP+drff/2tYLC2524eOHXN375hXGsQlX4jHAvl7x8jehxBPEZU10AzAxcwURIxBEE5iE
EbyB37ni2e9dB/SQB+wng23FToZW2BQnWpqaEkPQkurJrIomHNi8H5tYm5LN3nfDceTnwY2PgTjf
81u9vM3PiedaXsfSshCyE+6SOm75nBvJeIKnU1IPz+1HsjTFMBAdYgC6Z10ANnuo6guFAVzdhzfX
7QIrvP2xz47hj4lZaxHW+IBi9hYa5eYM2ucTs9opIrjn2Gxyy2ZMTOOeDQ1UKdsMBDr1V6Fs9+kr
fI1K6DmQKCmgyVQe/FCU9ag/qV5Wmv6YnvAU4nsUk9Z5b6jrFMcYtefmkDBNAnniGDmfJ9Fql7mk
0O8XKPKVirCvJfI9ThC0XfU7kgUOiKhMB+8zfe31LuhhQWn+VudSiGUKBklGuZuzIXQ1GmOJyFY+
VXh+v0JGhcKsGODK2f5CB0jlJ6G14Alg4y0ByGJtFpzTfmuI6KsK1DmOLFroo8MdXlvpASt1I5/4
vexL/+a2M9z+nsNhFNNdafFvuX3MctE4lI5YayWseOHH87ILymvRA90XosYGr5egkTh8ZJHSYgoI
LOT6JDXCqYS4Yj6nCf/UUpWn42nt+GO/qWo6luZ6JfhRN9aoH7dwRrVTI8y71D9++h/WCMxWCeiF
VXDZB8cGQ1Wj02UBX9ROtNm1SrktGtLrxyGTfvqCiMUcvyItbWEpm0JIlbZgKlKi9NatfNw03Rw2
4ISR4w8c9HPhP0S36kOFMf3Jwf7zYRPnlLiBWTHlZT+kQ0Z26m92VxiXvaBH/g1QY3o8tFpobzvk
oWjncHj+E5Gkh1rh3vhW0NYFrf7LHma8ZOh6tLT2ju+qeDV/U3q+al35ukI7G21NAnH5QLMbc8Tk
qFOqh2rNkgaGSapIP6KG5qiNwzpM3g7Bdt/d1821pJ2MHxszg02t1XskpYBUwkWFojkDmgVChtu/
Nmcgg/QkJaqVhY+7RPxAIpxcFnGK9ijP19/cQ9FoCVAGn/dOn0rMUQsB94lugYrYbWyTRMAPteoR
my+GkdfKShY2rjvMrKNK+5kQjweT4r5Hpj8eARfzdd/bdvTzSuC3y1KFsmVZ8rr3cMnqzJb2J4/Z
jJcDd0NzHZdnNAY3+rXNadi3yop79eB7RCxeF5QFQh5ZWyPqTD37epOh5guGgjmno03ixmZyEtCT
o6az3s8U+SRxKPfaOuaDQOmtm5tleMZWQNI6JGcE4ef/iyckU3DjTbAtevj4vRfA2Q2e9i5fZQQk
ujvChuhyVtbaCXHihXzFVjRqM1Bxd/HihPpW2/1toLyu+ZWkDKvquwPZPkEShy7rHP1B9jIZgkRn
UBWVQraycVM0jR/1mXYBzZrPJ/q5Qmd46FpAyn0m2XjDAeP4+tkRkpScGbeQMtJSgdCAIaOga2Z6
5KTVRfdl5OJ4tdwjPY3KQuC2yaFEVDJ3vvUuods2wkr4uF12Cb+tH5+cbwPQ2BS4hkVf9nkrwOqh
kGE4N0//RmKoYjonwNxWS8do7ZRjI3xUv0iUBEL9vwkGJTQdoujgPXWHTy3uiTj+uhvVDI9nCbs8
q54Z4VDfAd/afnN+br76O8ycVDsEFVzRi8d0znb8xgubLPVr+SPGSGEYxKgZso162wymjPxSfX1Q
w4B4SBb2YTOHrBhEr/l/kjR+e2UTIB6RgnlsY/aafvHuC2x72lotYr39xxBepxq3fQUblTH5a6WL
XRIqz70ozzNVwfWbwmRFvoYlh9VslbchT0Evk8ok4mgej/8KFMsbG3ivnkRvw4TMxKHNFcXIkSYq
0r294CTP13zq6S84VRLJg/DmIRNgYzS488OFjuupu59Jqub9yBrOvLn0dyB+7/RwV/B+9h92+KP9
KUMXieH78OVawBUm5VM3m8VijatF2c8Hlg+4YlEDM2fH0OO7hkeV/WWN7DvLoMt8+7vud6avkv+Y
/mqZHgh/Y3zRlbXA9Xa16ZYieC1BojlyAw0Q6VgZm40NCATqd7gNLSA1adA1RVN8ELJVtz/rbayQ
6W5qkhR9KciCbVD4JB7jO6lqHVnx4oyUwIQ4GtE9QscKNE5F1L/2U4Hk/cEv3WCqonF5hG43HohA
skSjaATbHrLlqYQw8/4NZ51AZ+F/Do7885NTMEN3a6ca0QVmeYxkCRggCFNr1enZdN3GR20V96qF
7r/Fa5coLH+MUVMkkyFJ4HeItUHkVzHTIg+OD7AZKyD4REthZgWPV79KwRgoqtPoqxAxUJuNZ8Ia
GdOsXfdxjiKn8ukqu53duA6VBb4Er3VpOctvGutIRgMDxj5++zbUFQE+anh/6jJtGK5MMQuW5Yw1
cu6oq3eoUQteXKafdVJywD23Otx1bzNP64AOWJCQvjDBSss+wAWNUXQUsP8SOwIkhxrmokxC0f6J
kClBJ3jlwaX4kyIwxIVilOrKQcpMpxg0C2+ZR5Gf9v+zpScTfXdjNH1sXCVVppV9ytqoDbouoI1z
CJLyvZQ1qFVC7tTCVo9U2UjOmCQO5d4zXpgT1HVL1N37xWb32deCtJU9jNemggzM6UafNEAs481e
ec3sK7ZYH6rDg0uRwVzZqJeRze68GXe5aw+shZSnoNxZAH1wEtkeUDVpNGEQgIjgms8JEfGPTXrm
zWCSSNlrro3VxjemCJzEZMDkw4N1GFolkKdRXGb/bW3BtddCgFR2d9wxQCTHAG+w46Jndam1zER7
Tg4F8dVC7ZJu7ScPPbQx91OWfsda++t0nK7dsIqn/wfsbXjK+x2VjeTNn16xHb/gVGdpxtCF/Ybv
yXz+0IBcclTNFiGprpzDqRhXKhoaR03LschVTjVdrd1TssuNgN9gyzP1mEclC1RMidefntGDK6CQ
k7VdVI87V9ERJ+HlE1MDw8014zaEi5XosBdQPEuXc2Sydgwl8wtR4ZWxzbx7xQRu32rDGoWZAMTz
vYT5y7OMdg7B8KbXm0PORyPZTpugA7SgOnTKgtC0uWPVnJDi4CkpJCbl4c/cVAitNb3ZzKHZg7yr
ARtonh3Q+/yb5/LaehsKdmpL7YBhHwpe87iTzhwCT4LrRuhNrHMRz669ZLrwoXHjpAcveA7Atezu
/8NJyze7/a9cdTXGVtDdhOfM8ncr+3C8Ior3PHRP7HjSDcgVESjclC1JrBtzw8iIticw2ogh5Vll
5aG/RolP9UtxO+oBJD5FBORV4WgwVZQ4P5GPRjTC8P5S+EbmLi9hl9JEqs8Q8lVLpwIYHERW7HfF
oaa+SOVF0Ed1T/p3Qqj8APHW5tIdOuWyIvTTsNQol55N7ZPscNHcx9z5jakfJ7mSHHmQB/JQlAdf
FW/iQPfyXPvUrfoggqnwou/V3xZAUS3PghyYRcjK1+ZNeeoAAqh7Z8PtEvd3GH/D/e40ofg62jKo
YBaEVnkJzU9WSgArzJYss7HlvuYHuovNcHqLw9eVKKUI68fgLfA8ot/KgGT/gon2pah0YSDTgM1H
oCmLrKm1FkUvP2AoV+/uDM3j0t1zIPnG7xi3ANVVdVtZUhuwKjjKObeKIdKgMAuWZvCa3DBZoY5H
VS0n3YmoOehc3AvRychea/pKkJXHuehASIKeuFxIuFllK03PVoh2McgTzfig+/O88FyngDlQt+YT
iEXb/0YjyW/9nKOAo7x5PELlvVkGvphNoY+j/jHig5oP6OnscjG/sRl+QQUG8mkmQRliiiq9mHSm
UIucoVh8xoZaLwdARnz8VoUmLsIpLFF67x2yRBQS1lQwu7KYMX1twWRDcCgRsi1htb3t3x9nfHIE
CmXc5fnzw+c6OGcDCuee6j+iur9wrVI13ENwQJEBVBhreNTah/PrPODdva21+FS4KjiHaJmRaeog
rQIYPUKDNjhCCBv/+dFhWdf4C0Rlw5CfpiqR82WOqjRbYKFxh3UNahl2NzOlx+3dhGiCQIO7LyVQ
iYy1c585eEDB+cc6E5hVfslF1vTgvAkmnzXHvreCqsRLHRjDS2lIL7L1mo6KMV9H9LpOIiFPHCuT
7jW/ijW2w2K1z2Nc0yPmcsfGGhNbJ0uuB3rlxtdho/+gbr27DQr3rQf2r6ybpiX4Mvep0tyxPQbf
HW+7nHefQGIklIgEYmN3JeuNPalOZPHo49x+SBsLYw2vCxqgiFVzys2vF0EEhZeH95kWkuAbd1ZE
0TBf9Uiys7deL5FA0Wc/mHu8XJf2KgetKJVyInak1v/CgyhWkSlBULuWszv6mJClNiYs8o4Y5P92
QBPvAkV5BtEWXEFZSDsu1rxJyWKydcEPU3j0LnkPVCqgDXwFEflLmtFkeOvvLcJg1CKS/5dma/Fd
QCA4R32R38lnrbO8ueVrxkMDTG09Drhz5ZzqE/Q3Zl8aCNcSou1sSi5YdPpyCN1O79Naz/fRpfxk
72Gab0BpshhaO2iJqoLZROiBfpqHwJvSuueEIrKA7rPPCCIiGeafp0nXiY9eOAINtEVdOMMkkE5s
m3X3fVUaU+LbI8ul4+0I+J68Kw9cF/AYkzsAp8SlyKd+qMagk/3duAaqRB1fyfawOvn7ozKe4JB5
lmt1Mbqwoxk0jhMkZGXW2KvvSGoYPZ/62opLKW+aMneon3rbDxuXbWRoHwtanRcLH2ouinXiOJLN
SMai2tsqvEHy3TB5Jz03eLgVwFeO1Il+niLJxMw1ONkZF+7ws5TBEhn+/fCESleea14MqrZeg7k3
wHktwXuw62my8useQSTg+rrwpcf7tPtSqQtGvVyv/sf9o5+hQCkLRDxLQyoTKNbZ7Xq0MMUYMJWa
dvewCOU8JX5WoN6+w1VkYVbf3WdH78TPLbHjDxRzmEXfVw5Vcgi/0oMErZgdQVZ2BWpCq9Qhwq/C
KAJSvw/SJY3xdqEaekpEbkcfBlLruR0alS2yl7WIwh0uMTj8a8eKdL5UYgU4CJP0qNCn+xxFodk/
z752v0kB5Zl4XB/B+xIb0SEjp+K6Ip790gp9liMaL+qKYcY4r+l8Q3WfjIh4nAboBl8V4pH1ILWc
ntmdsWFfDrvnMpDdcZ4kKIpxO5aphLlQbhkqe1tFt6YWlp1iTd+/rdLanI7qwK4fiYITeCPGv/6c
TFJvrdcgqbgjtGGFsj+Qplm5Zn58OWiP/gvTVsxLZng9q6FZylS4eeOd3kJJHnXha1nLMdgVXCR1
hPM2yPrfKJZqYjM3gVlwQtSNj5Xec7r0+cgtdYAltgBNlGWFRNm3Apnzhb17V2VVdI+5kz/7fPAg
76tqQ0kYbSSr8jB6e8gZL/0hcxAa4TobfVIota7WGge6rPx37z9Sf4wSw2zijyoDgWnQcDL8+9UY
ldOzQCa+PqmBQY6xXfxlfCKSFajixIzqgL0gpKsBOHsAW0hw+8DLJEdal+BdphGb/F387c0iSdwu
htximwgzb4Zt8RYAj4Zja/WivvgpOhF9hshFDD2juMOvm0I5Ur+zxCfZ69IszTIqnd0LS9a34jDz
OqjESxVsJeQ9xcrwBthORZUJboQS3rNwW9N/ZqYMG8wBlrFaslNCQZ11Y7Q3qiyUzOuH1w0NqYYJ
DvG3K+k6xBLtPV9kawo6o0RGQje60aci9o8snC7Vto+2z1JKFn8wmZYA6vkWlBf5x95YQxY5YuTV
ORLKMd+YQd1Zenlqe2upFtlysgdWNskIc08xCic52MzXYBZDMIhWBtB741QOk9I37pAb3HfEwCQ5
1P21TvI09MjLLWNzSbDNNBpITIKyQ2S8c7odLuksJZJjeQHEpRWIS/Ye2DkKG7u/kr3S23ySVCTV
adJ09VI38OCKqB7bP/Y1TEToUMsOB4tVQfkuot6KzOe/ftweHlGsfeNQ42+bqPVbULRnPTsHTXI1
cgXaKpouKfKBAv+cNop67CJuTJ5l7VcDiTyruCxphsLgxB3hbqQJiL8dTv3i2D3EMw3V0SuEqyJC
7RmNHKisjc9DvQNO9m4ag88xY9jRzOnpzQD8jmHV3gFkSrMVzAoNoZPQYovsfjAKyaeITCqQ0d72
8NWJK2YwUoO2A6ezgifci2EqOz9tZh/r7MnvFGjKbe2Hja932BPa71e/Ees4wxPXM+sB++Zl9fQj
3IG/naVQZ6o5cJeBHBqFiJPLPPzk7T1DXeLzpmaqhDoDy+sRroo51HpSlgL7WsKBFCRy1btV7+NK
gJlmPxooeArQJoXFnL+M6XwiL9p6H98NEII70eL+D2+fIqd1uQ3HgQtxNbSIgJXkXkLgRr7fKsTN
SQEjzpM+wQZO5nrK7Gj1GCxKiYXbDyuet+h3CvYyzmP3Vmhfm1LtOPWEynWFDbN4/el6tFKS6slp
6bFtmWKHE6NeLcPMg5e4wZ4QVyMs63O5nwQsCaM7Vr2G/Fz6ddVz9SBVC0L0CFpPWanRVP6AV0FX
dL54XuLcOoqXyXSontocwgIB3N8YWLhqlqvSidaaKo28d8Oqy+DN85GztMi2jiaOM34fk5hyUQaD
knDTzaKxASTHJ341mhZyyy5qaUFDfZehli8BXn3HZPWAYZoUo6F9xo7yqIFuYq7Ccs8LOvH53pRd
OADeCVoSVBYI6rqBysCMXhjex+BDOtbrboiXa9MhIkAQHOXZBtw8wVxOGXkPp0Pz6C4lbqiWKKan
1e86LDxx5os+gRBr/jF+qjvFyM5oJnM2fk0JVQF68p9jOgDznvHgQ4P861jHytUd+k6NN2M1q+Q8
fQPjrYvkHDbtutWMAIlCi+e19KUuxxGESBwqEyoThP6edYNlcaW4VYuarTDJVid+pYtDkfdJxjla
f/l1oXZnKJuvZ0bF2ZaZVs2nVmYu+N0qta1K34bYFvC6UOVJr2pTvJQMNsQRO1DrFh2o884J4Pg9
YhFGHr4eOKoXqsQjjYA6rxVSmpenkmsL0KB2jNOD3h8xEtJ6HhZU4l851M2JUmaegDBozcZ3IXRZ
Kc9upBXax7j2k1RJ7oLbnbmyYdsf+Qk2HeVkGc6rLNBALm/f/zN8/DoRaSZ2R9GIxyAq9AUlMK+e
RyqXuL4hOYalcUZMmdOHcIVqLgXy1gy05Df6Q38fFtWwvchtQ3Pm2xODF6ERaxMfLrm1z6GR/FNz
C4jyv7DgRudnK0F88YoJmIFAcRjiyM4S8S9+chWr+ptmuqEWiAvjRHoNULdtgHLR1xsDdj+S7AJs
qgZH/Wk9kHZ3NtpyYHq8LPovRvtrj7w2DVPloEA2p1OnuhdS08t7tWcsYydMi9WKJcu4uTYuGc8N
mdklv54fXIU2U5377dsj85ERtc+kZMggSy/3tCiUMIvz5pvEkvOWoZGof01mmF2n3G/bkXUU840Z
p1pQYhRQ8fRrenso4ZMbuwjtIyFrN57ropDnx8ce1s9I2TYmbQKF1SXXo+RwsPOIn19+hbxpylOz
2FcAmG0zINPIKX7Gl4px59uFteK6Def6ZL2QaScFJ+c4iou6IEoND7cbI4XxTGkzWwl8b/7kEY9a
hZ/yBsiAF50YY7gLv7SEtnhyNDuA6dRyIsdWlaPkgjpOFpiwY/EwXMYnGy+MQHoziCAdxSno4l8d
afU+MvS/HaEBvGUO6Wmsx8XEoUUGcSL+uq13czlQV/d4i5l/tqFff618nbIc3wHTHLFcD2DQ4+cg
4O4AERP/hQ1DOLqL/A6Am+9oq+X8eTAUFFSUJmhLzIXdl8gQL5czWlbYR5pAJvrR951Kbyo3IEDl
l3HcAyZXInjVPjWNhudZ7g4/RxnVwyOcduDMj9iFX42olnDARDI7xWiRR5UALM7w4jEWX+f1Th+L
sCkC10EK9XefLds94vs32sZfog3TzFcRBUmMyO5jVheluUT2bBWqPAQBt/0ShO8Txh0Vu5yaqbXL
mtBVHAgPA2UK1+xazQ4ZDMKAY3xIasfFSeGfGEqab8yTbSDycBeeiaKKLboSLL/UxxN3DzKa+NeQ
X2QioCwr9kQ5sXlBSqAUj9kpvDi3+XXaiO7iWiQ29AyWrTg6ZvZqmZVsPQKQ/X/u0kR7BTrHeu09
RcKvaQ1oSvjILgJDqyu1NktNzXXQ61R/7hitom6yPbc06AvS9WRml1Tydgwob0QQG0T4v713jYrC
WoGZJIJOGXhG1D5qpQ8+TSaIgpyrlIpzaUv+eRfO6aJF9mX9SLVckT1H/UQUi0VYAvVYyaEoG8/X
gJkNZPESZdsiPh8SnX8Cu3CWGQkawtD8EVnY+pJledmpCTjPUHk3luS4alaQtXZNjwYBVA792ri1
1XrXnUixm7oRUp6vIn2KWbakwP49IKduq704kU+OUyfTzhY8oFpJIx/p8gjNUxoOA/g3Dter3zTN
cTNZfdRhXcK86cD3QRfB5JzyzjsdU/sth5n38MctEZGW8EQkxNK0t1OBX9ZR+ev/q1xNp7ikesCF
fraSivZDlOt6FL6bfzQMUnX50gZ3FD5mKk2UsddreKT2u5RVIA+2qp2q1E9wp1zfuCoWAG+gGb+t
EEULJPYPvG2wqmO+R/BCTJAcsXlLT8uZQWAHTVzwSybHF3/3hspiwbokzy9MHNlVnnhxLU6QCtjc
TtboWoXNXek0lm90ZEKm+9SmF3VPI+n4RNClZAwEfBwI+bPgba28To4jom2J07+m360q4KTPzbkA
3alk4Ez8LVdgccLc4OjtoXXfG6VVC3lG9zP+E7gzsJIDdu2SKisLqj7f5nVY9PMCmSBG++0f8Upc
IkLfy/Am/iPV3M+ALqfaFS5anuJU/0hUThZPG3klUr6k+cCyOALtMEv75PRSwE0o6DQGvFNqVX+Z
8D81+Jfik17ww1tTuC7KdSy2XLahSboXEjERZhy29chgOQ+R8HeiaM0HndFWoYeE4XVKKJ6BgohV
Kgfe9rGuxgB+qtdIoBZ/h2v2MZgL0Hnran5UahkHV6nKJM/QV23UIQ7O+akJm/WY3kgGUsTFZitU
pXrqnpItuVv4yo6e9spLbKmAwJ9q3CO+FG5SlDoVKfh6n8YgyDBGryzfbXanWxPl9DatyDviYZzs
2Da0L2eh3fhY7G5UZ/7mFuKoNjllopQQppOXWn1Ou3Ld313mJ2pvkYYu3BDHfqpzpavqxTX3i4u4
s3bcicNg0YNt5XfG/qkfH205K2Hxo40jhaTtNL5mRiNpL8kPgJX8ERGOWHMRvyuwN76w4r2TbFRD
SuZaXNyZm+DS80flaQoc34Hw3D1CwMOD3Goo10Ck+J/QiJEGF7SaW077Ard09EjsikYjahYVAEuF
442Eu8c0sOsMi4+hOogPCOSqclUT9GFSD1xM3+GwwItSv/RgszngVLyjXtGPiWMjZDF7TdCb8XDq
dAjR34qriZtut/U6PLGSf16WUFAVCLxmdTRepjjjRvn7tV+bd9wZFdvPFbzB6mhzHP/w79HrQBeA
lFnQtz9LiFYwlO38NKC3/JQnc7KU5UwL9bjx4RGdWrYW+GALIVSQq+V21IB2OHUkWcrWJ2BosqC7
ouh/EGkqqRKFeOGKsdoxTp/dK0kSEgN4AiSVb0abLPJFojicjwJVuN0tBCPCkYKvUyYNjS+2MrUI
r/RyB85dR1wdU/WintUaTbBORLY6IY70aBZJvupQg0FlhPyqhcNP5GrFEwYjtKSVxWWf5v0R7Krq
UlBNyj87Hy0TslPsd7FGQB2725cGopIRiDiKEX0BRCtkviLIjSG59Js1e0qOPBkrZ0ogSESXu0we
D5BuBNhvmBkf4kIDPu+sXP16h61nZLrP4CrE080o16cpTa/OR0TbDowVugI4wGcxx4g1kFbHzy0v
WXLx3WKuTzV7wIjdb7jnPbgL7l5LjGK0VN684C4Dc7A1G7Sjl9VNWxw/rbPQa5UOkCM9kCf42UHB
QlsC7QrPlpr/JOyBbnMztXZOIcnbOS/mlDdSlEann6uuyd0O+V2xINSaEwpTx8EG6sl+IQ8Pmh08
sAucSgIX/3aqip24TiAtxm6jCzG2g2a3wITMzaqF2vC/ucrJ0cLUpigl2tFbBGlfkKNXmmzHXzRH
XbhD8TL9YT4WHPZRoKgOls5avfdf839nTEcdpgsOUMPOcYN70/1ErtfligcoqafxLETwXdPu1JQI
AAYXxJj/y/CkuhuIB9Ntx5y8cz18azP+a8HmwBSsJPkPAGjlD8oglZTgRCCDaHS6LCacJZdFqajW
ZjTEqex3YFTOGz8kLI/US0cd6sRITGt5tsOlV1P90psus9CZ9KxSQaESQmOwrRlSKLOJYg5EQ9Gv
7T/LFVkP8+yzG/veO1s90Z6HvfPrxXubMnmhxYhYCpG3JS/ivr+tCy2B//l+UWB+op7leR0Eo3nq
jZpVEH/tITb7NhX504RriJAaSwgKbW/hhATfvCm+vIT7EVerSwdntd8uBI97rO7ffUXWsTIcohv+
1nLpGpPszue1WcX7BSvfUccPe3uekv+WLIwkrlBgefgVca4wRRa3WGFd+DbS+HZTVlZiEyS1itKm
ogBJqy98teVPrgd0hVVQWsS4NVrmgXUCvdNop3rOV3T2rUOkos9fq1cT+pjzCRfVDsRWkio2vqRv
KNJ8FZ9Nxguj7c3tVQMqYi2SM7Nxj1E94PUbn0Yy4RSh5W1yO/UmfiYyDi2xIyL22tdEr4SFPYaZ
xtc2MeBTbgjoUsRLvuNKuaLOfAiJrZjrJudk9N2KdL1vf/odnJVjoBB9MxMPXbV20nFVJpfqQqlH
fA1YRkOrqytnhU6FdJhoGmiU2P5mI7+rqM6Qj28nNBKmeQ3MeV1qpUs/AX0EeMAQgoIZwjdzA4ug
w2zW8eH2tshl8vu6xIXogAC1SAj/I5GLPT0hO0ydO+UvPwTDM5qg5yGLY/HSq4MzUaCq7xLc4L8D
v6nK6pCDdWnTzm8dWIEDhf0B4McAiv4V7HPOFuR5FBFMOokpKZgfJm/uZawd1aXFheK7Seu/UZRX
CzQ4zU3POg6VLpGl84dO9u2+KnpsC0QG4oj5M/VZyDvmZ+VEW7rCNHMg25FQNC0hC9skRqahJWof
VUqaCfJWBS1tRm+BGPbzxHPM+FSavfWK8+0iCb/Vp5m/x8cFoePmEJjCRTtn5b4SLB4ZUlDxxkuk
JOiq4OZWhhJPkH7hV2n6hvt7fnI62NwFgwTi1JEXYkTjP3z12Q4um6QiCaE8Y8rWGfwvHXBR3OLs
4H6N7uo4/HYol5X/MuzDpXQMbgPY1sYVGgwriIX3xDyRKicS8h0M2ZyC4F3NXSOMSboeCQcz0Men
oodG+qnetlttMYT4L7ouAYezkx1anGXt62JoVPlIcRoc/hQnjndNeHDDbuZIBFThxAKFSnr87dKU
nmOwJE1Bg761ZxGP/dbxuiaSp77LEgzYq5C2kiZcK3ApjbbEb5wr0359SDYFgkUGemZzNAySmwbd
7z7sbsx3tz0cJk6bZ1nCl3Z7r8DDqwNFCkoT/+acB6VnIlNBoCMWejyHu1rGl26Wh77dHwoUdhD3
XOFvQHLimTTBZFxJIYxHprXj3WluEpzLzZYXgfWI/aiuGvHkFDzZRAy0fkJTWeBKzmbHJv5bJVNy
WQCIETzk4ZqVDIM7Y7d83wc7e+ouXWASp8JikYOjBu/18C3Wx5KYjPwKRkEDcwfiQAq9v1T78pXI
W6ezvJtSgD47EdcggrqG8yg4blLgM59mpKe62g/JrIBGZTS96yY/R6FmGGtXQuWoENnQP2/pJ+9O
DUxSE/5vxhO2gZtAIGSGv4W6C4c8rAqn2j27ycFiEhXLu679I63t6BTuYPIc4o05b4duXBxpgeUE
sNxKytGW4SDABCpGlSRcVcKiTLfTdN03GZMLhPdef0Tbi7qLPr16nY6wXjt6x0flDqkG/V0M9ZoK
dfEX4a7e4hdat7uU3P2T9q5qGBNJvuYduXBolclnhyazzFeVO0OabzTYOeBRDc4arryM/L9w+Zf4
OzPGjoUcH1gjpgc6zw4kRi4lnN89IpXouqRTx15exoeqqMyfFfyJqqhg6Gl9S3IrwQvA0nvNh3yR
Y2nf7NnU9lZIDbf48yUvotYWt6krGJnKyi90dugl0DAgjx3W3Bgv6rlEO3RmCijsMfAzhZW7b6jk
l//uFEAokoFObTidEwftwuGppG4m3NUc71YSxlc4k5PAo1oBPWZz9iS5CYFA/642KOFxlMFXWc5A
U4wLG5JDOPqbGcMK3TDSfvtBohgCWarHb+NKSSzkdkPlkqTiOY9GEnBb3qwDVXKUR3wSyuXsg/PI
SIwAj/UXUKw4eYa8teiMwqoocrN2eDg0NBi+jS9JNdyjVinPMVMMpDlgAlZLC0BUj7ke6rXE77tE
8KowhV5ovjSsK/CoiJ/ETp+RRzzqG+9PcFp4QhgbiFitGl5F6CN+YQEgTN3eXTWAI0FfO5S+oGeU
srb+yXVloUXk2MFkNZhOwSRBdndM2oqnQ42AqHtNHzvHbyLQ1SFr/wJaRmwvoxo3YOtY1+oxLjHq
/uB3wmR/jcP15/gmhevTQ1WCJKhge7HCCxWVzsT7qFUIsa9kWx8KQHQxfjllhU/N6YXFDHabNEAH
3d5gUhqfDx+jCS3Xsq/fmxYcw1osldPzOsZEdrBf3F+COfLdTHGxz2SSbnpJVBg8r1u+I0m2rXms
RFBO+g26/wMUyPLLoCBafv3bDujdl488eH8uuefZA7OXWmwRC2/dyhirvQeErYh+myCnU9+z+ka1
BI/ZwH/SKwX5V0ANN0q9Bfei//4yXl+HOFdYBaxWpc2NlHovD0CHh5yrgHoEHpRajmd9w5TnO+Oa
DmmHgDH3VsYvFsbNfA1r6qYXOMTqIM/t3t7+NYcghPpbNVJ+O9vKhrSY+Mte3sk0RGc5+ZVsSk+8
TygM/ekDkQhxBXglxBOUnc8joODcNzNJjwkPXQaMu0A+XrA7LCRi1AOoCYCuZXcxGarelKdcDpHs
xbpXzziqY//5vK3RB00KAa3KiM/RUwfTksiCmpO6VIIqUkcyYwp0YP8EaWzM/8mDYsyS2/r1UkBD
9xKIBKcHpyxdM3yBA57BLd+9ZbwLzKuku7lBaxvw65imxDyGI7RiCL+Tw0uX3XSsiwpIBrhw0JBH
n259dDuSiqwq6n/u5csbKKzZsJDnPBFPF7BYTAV5GKnBtkBqFa/8psLkTmk9Wy+iHHzYblKEVYu4
aoj8mKJ1edHVaKfbCBR1G2B5YMenA6tubGU8BciyJ/eU22icXwAK84RNbdTVvb7Mp9adD75vB1hS
Tgy4imQBaA5xic3Z4b5S84w+Wx6TUrGziaoYpEIbM6qEjwqZuhYK0bK5Px5rUB7Mqpb76UKglhgP
0Nbm3A59ZvjzPgPHjtpzkIPzDOAZF9ldiqbzXtYzD9WFUNeU6Ww5240kQiwPfW6Ksod/RdSUiJZV
wP5sSz8uYqgplAabCdc4S1N7sP6UEdI/uynw28MbX+CZGYoDKyZKFD2jUOyvUVZBYEQdSaEN5Kiu
zDuiMcVvhYceR9imh3q8yqUPvg1G/YDTMO8JOaWjtS8YPHfLYCG1WaoCkBvRCfgLtxMZX67+u1wA
iEy95SCCNldcd2Nx3V2r0ID5ESdE7L3ziLat+BwyGd1EfECy61qSYYkrMu42STxwcKIOtbW4L+JW
M8L3gQwMiMBQ22fsJrX6lRHM+VMhKmqTvlL1H4FrQAAqpJGXSvJs39Et4HcNxOl5HsddO9uZo69P
V5oYP16tcbyHFTxWHjyf4HJG88b4D6/JfZGIe1nqoy6IjhYSyI8bozniH86dRvOBXg9bD6cgnDlQ
iGZOqHIKTPHa4hf+6cFC+sd4ymWzBkNXk2OAuEsgTEOaNpDALCr0f3Cc69mcSnX/fhHOcPEc0G96
yr+vc8pmRRah/BZdA/KBzgT00lqrsfu+BxSK4zm4tJWQ4GiYXqg7vgIzAPv7NRm4CHSZk6IX9Vlh
EgaMcRRb4QmL9PXHuCV4zMaPhKEVfkSmQbgrOKQDB1MkcJw+lMs0JBZwIVQ6fbIVs61sEPT4JT+7
72mOstUlnu3JpfTNx6O14UQDsYbOYRCl1Ln8VgB0Voz2Unnalw6bTFgc7oPc6WfB9HAWyef13QPg
/nwI3b7/U1u2MI8tVyORXdPdaVGUBgMAEw+T9bFsvz45NHWDmflq6qjIzWBVofdgfNBx/try2qhu
N6FXMVWcIojAhVRpG8+6KsmRNUgVcdyuUMkSWIjhOFdsl+L4TYIMAB1qqTAeUVPExV1OfamYW0JX
54cvlTTLKK/HPSggQuZrCQ/L/nldZP2Tl/KjUzaUtFpLCqYWcGMd1UnyMdYk/AsoYsoSMySFgKVz
HKkJJlWMD//UyUmokLxpt3XYtXtOvLmyc5P6legXgf+jrPOWZNsHIfUyi7d9o9CWVa/Knslh9HsB
Hfl6gA7LNAoEdOoAU3R8YSykcg2dGKVtobTYDjLzstMK0TTAXedeJ3ObVputGIzhvNUrDkPPUMSS
qERpqYZeRBO0p9RlKpMk4MB6eUSFjeuHQAmAbQJumIooPKV29qGJ7L0tmN3PE9asTEby4VypnDxT
SBZe9hliEsoONd1U/C2GHdzsYh25NlQo+aHT7nUSyktMM8pgmV1JH38YVnSJo3WOKUsgszuemuZv
XcrgTHo5e4wzFx3Nrq8K6+9iY3WPldJBoEKzrokU8lcdEoW5nOQxnrK1t877zX4vvoLfRbQmpfB4
/ksyqGpDGvC/6Qf2kp61pZDJ9HZrUPjHin2DE2V3r0dCt2/tlaPdpMbPjU9Ek3vt0orLaVtAZMBp
s9qq5oGtCXfLJ+OyurHsrgR4jhp68MNSgYop9lTn+u9/lvOnmXY5VhQn8jxX6yTHZnIyepS/64Gt
wbP/PCl2I5rco0IZPR3w5d5eA47ULr2dTPB2mrLzH0W0EDgb5QmZmBj7ZmyHCKjWhB97mijHq8Tn
a1yP9HgVdgHDvFiXOSeLKRxtW+UhlR61gTfw3m0I1a6MVK6FvhcJSfzHpAbcY8G4XVfRwnllEHww
kvtb6YgLzhQGlIL5+VdDiyBkomnz+Adtq3779lMXWsHqJebnpvKzoOm2INIQf1Y5vTTdMGa/hv58
LWrhLcrN13MxcivSZpUQJAOijhbWoYlHuWGwcN7Pa7DyVImdA/T84Qk0CxY/wQBDp4MA2VILRuGd
oqn8me+caDArhdCK8b8Bb395L7Tz/YMmQrGHSAQzMLk9d68AV7Mp49TgHtAKlyNXcQxRokFhZQ/z
KsCeuFe+9YQIjwFfjnoYOb7T5EMRCqReiuMYxnOdWBdFylPrIlGkLFSp4U5KjvTaRdC5I/GCNQHO
oCbqSe1k5qHxkdvZwZm5A4PQ1VJucNh9lQGCmS74kYsGNSpLLywZFgk9pt5Z3JXKMvF2AjKI33W1
vcaWE3nOxtaooyjCyv14/ySQ7lJdbr+/dbZiR8YJuskM6A5SjVYpZbIKBG01RpstE2dNr7hCcwlL
/Y6jfIkBevWkWCnp6AR88I5QXXeL1dbr7bqXuBFjtHLRqnm8ST6jQ4HtqvB5tPo2Mn67Hp8HDkG6
XqkRgCtIo/xWucVmwRUOLr66WGnfTj3wTdk+TTjBASdityxQG08jiVYNHMhdDYezLvvjJk1BdjHh
qjEHczHK8maQ/hr8B65ldgiYw6v4p4fVgOy0JVRiRi0Ou7gzHdbLSdI4WTnWFSLXc9y2QHBs5btc
CH7bdIYeapNzEr/s+HZCrqGUc3Wuk004BJTwH57TkvjYzaqm/cDcM36DMlx+CJKbxQlAOdtzypHL
tGhiW70lgjQrXUYJ0h8AIZkxmQpdqnZXBIPcDMxfiVEBlx4naSjKr+YRjlyC4F9m64VvI6m83tDQ
37KaSpBcgHlr6XRWRxsRDtTVL+Qwzb9pdePHnWtQW2T+BTUpl3klOqb51RgbE8FqQpPmdBfVFHIU
oeN67L1+66wPlFWrUYbMQMbrcoUuVpsJgiIEFtkwsL20Irx8NmkegeOqL8xJoPnPqJidqhCKeLKU
FqFcScUEE+WFkiF/wOSAv4Q7NBGmLC/b/72vJmmVAU0CqSClp/g4941pzcV/1K2qsiDQDBwMsuE2
quJMsqjpketBsjaVZOzhoTVdi70cuqNX8wqyFXZxpVF7xDbS/3ABYN+np9Jzs48eG8Snj1NkuT2V
TjgrxxoyVqzOnrvRx5xRQF3745cza6LstTDTGAVjgYkQ8TUrBKFdw3SG8/BR9w3L3fEYyO9IOM0T
3n/zW9ODiMqymlWCWIipOR99RldDgP9cSVB7i5siFVutMDaDU1HRLjHBPzDq0TkbAJiUc+pxAO33
1GGiIOPuPg9DgtVk/iiHeuC223X7hhYoYOsDYgC+56Hj28ESiZ/qIYeh6H4PYqAvR5EhT0cAIkvY
4XGZnMRqO3W4jtUYPbstfcHa3gIvH9lkQ+F3GDbRmRWcBo1C2XXYuPwUSJaaqD3ACmM/Y9R4w7qM
2xbnTNgQGJMXGhkeicFhjmVWfbFmKjR2wg3RXb8WZrMbUO+qmDIR9OKuvjpANRZX4/rftSDsoWcr
iyDogihokCVKhOc5V/7a84MqHbcOl4M/VJ6wtbCKOGziyyz0hVC80ZH1fIpR3TKSJiqUtMruX2oJ
db/FzthUCRZ1CzZobWx6vMceDFPakqBJNN+2flJMZOHqPdspUp8cwrExrO0ndGYpnG8HM01IE7FO
4tJ0VMwqv1G2Iq/iYxOAZoJZEpuPeD+cF9gPNpVwUpIHVu5170gUkzLMIBrasKEjM41tw3VgBq1A
zoecB30YkbzvBE4NMD/0+Ql3s2p1Y+uJ6qC+wCKWrgdPnCt1GpcSSK8pzvX3dzzEc6At1/65T5hQ
rvnyas22Sm2qYWMeZoMw2HN2gOEW5ETbu18qiW6doKuRJCp9l3y/EjUC5tPdZagEqBDHMZbZ6VVE
1qjTw129xRivMVJSY+aEKwK/l0eFQrYhOeJ40YxnEK/OOnh6XjvXTdyUm5PkWfdAsnBImlHxAqtF
t+so/1BDcGHNUUS0wKgHh5BKn9mUbrGMdZTUjteJBEEp2WvJIhKxro0YTtL53yJjPzsMnDt0mWpK
/AOqTGkZrj/XQr6wRlA1ZbAa4EcBdoXjplKJOAGJTVyVvkbuYrDbRq46jNqlR4p0zVqIdLVMi1wB
sy/mkQ+bUEXF2kMWipCkDgygu3mbsU5LFC2i/9xUlUtexq4USTffM0N7QRrUFk0SQusDAUiWwuZu
xHU6tX7OstcnkogDH0vvBtC2aNKj+YZ8bUdGbgADT+AAaJnnNrz10MG/OkCsgQZ/+EFLoSzgJwsp
7srE6BMHDPSQsBah4K4qG7tlOUe2o6+2DXlwgayS7yjaxIZPSB48DSvMlduOhI4F8FF1DD3aTJud
FyewJFPsvU2ZyBHkxjVnEBzumuVwCOFcdeGV2sYYCp/boNdGth67ex7R9JGoRUH4zQcj7nA4U/wJ
UFy0eWvyXLmPzepyad1meDMKSdrw3kvj7mWxQy8DHOQ6VgKt9DQhZwPYNjakRhTirLpFgs3gk93d
dhmqYV0YIDw/uibU0+jgzuGmlhTXO9PXrd5oAXDCrTdmKGYSPLKj18Qo6pWOTjkwEMlTAKh9bDSG
j8cgwj8uQjqq9zFS7fhttzH6RHmBB7odrF2q5AF0L5jqWVETf3QaHRmO6DKY78/agAnl/eDMdY+a
2+nXm4JeKbtDdlHDJ7dZbu9oVkL4pVBn3d9U5AnIUkZWkQXVIuwI5xWAiQhDWavKFWNVCoT6zynU
iCQaYQMSW6yKq1h/f+oZcKmYYHxCBoFS0BO0hdmWu3M9Nhtqb60ezvbqYEgSYnLYO/p1iVJ8SOqn
y7CKEdeoos1f4c8LgZOqn8OxjugdTpBsSf0fur57vlhDu6aQqNj2O5V09ueLmsiLyOu+cJb6fHdP
uo3lpkjuTEpofG5SOCuRF0qIrIgdyPC9YULeGHBIeG5FUwvK+oBM/blLOsldEyAYKFEW9E6Zi1fS
v0aOaU+Im4rXTFxDTS5wn9hfX9yK8oVtetNoWxAsIY2rtJ645p3gmOb1/IjrOFu5y2WlLnPzFhw0
89HYDqwXv3lgpxQgKXDGhMdCNAHVkemUnbo1hUkHkVuoyQSQTrt82UuaVPQHpev4+3ZMXHVYfMG0
aTrlvv8n23rnWvVeTydpViga19dy0X6t13OY9wuYoxNadjOF0VAUGCrG1MMvjaKdv5aZgQoW9/Al
7TNKOml9qYtkIrGQmQ4mfpSkIpL+OYLfa/pFbT11ZmFYtkN3pXE3HGtPxC29PlXK6/nCJJUdtgfh
ZmLSUzon18D5zUdNQ1fgjVIqnPbpl1bdrBQqZ9EjGs8QTEGyUwJhzzkJYkADi/68AUJUmY+aKJQD
7xn+GWE0dwN2Jh/GQtp9Vj2AS2AOsqMtpw1oqLhModuVRtQ235AsLi28Cvy6AVw/m5l9akMvphKB
/eKY4JW0dboASi2x2O7RouH4QFoS3GAuRHs4c9gclghpQEPz+6ZCDGb8d8Vmm2HkvERlfBrXZWU6
eKqypFEgjPgdF1pTybAQrH1MriX7huaoFdVGC+PlCoinHpL4046qK2eVga+3wJM401K6u4GCG4Dp
W4N96/3+1rZ8VM3NYXZYsU4RTfz4mvMWUpt6DOHlnmoLVB1YwBkyvdlyD0bp82cEKNcAGWCMrYxa
YeTM0Ufz6P5mWS6c0Kggny0KfQhWPyysBpziihVvi5sAyg/hAIBsAK+vj6cUNoD5pwr0szlJ89j1
zMHs2e/fjFOiBjCBNac6PD+0JrAjjF2Rne6xAKGS07ZcwOIkN/m6pcJ+RdH1aTi0pJPzWFQNCC/X
7/Z1M1tNFxbIioUt80odwEfCZAGp8RVI4ujnzBMfnSuqpnPLn2H5Qxs1Pr/TpTm3WEe6b/5yYOo5
Ttc/N4d0oqu0WkekWDH1VecE57Vgf7xNMLJoRcnIrAF3ptklX//PrIn37jiA7aMYVCELQf4+/9or
777euwklO+B+nmhQ/Z0lAgjM4NsSBo+EDaGYJhf2rmKKAgDp4MA1lxEG/acZb5Jgj4ji2koBWuQt
NhiX3yRoLaT/AoYwUMMh6XHe9HNZ/HwEBUka2qqEOp4nzbVc3h3rM8Og1jLs+1hQ+jBCZi24hxdd
ccutrHbFpr/oD20yvxWJbLadxusRY0AqZ2HXLHnRy4OUKhGvB/fYMdS0stCK+IQ438oX3YBy5yb7
Wl9chIMASMnMmuII/Jcl2q5CYmhZ9S4CMNKJ3QECi5a3Mc5bte/6RQ2VozuglpJM41yOoomKAJ34
yZuIF+oRSt5yXnS/+d8Fw5UXV1kHUemLRmuul5McPzt8ubhI2SGbOxirHdngHlJ0C8QlgW2Sa3AW
AsAAfXbosTdCik6b8ei5yE0omRig005PCOoG75hY5/86+Vq29Ck1fx3TpMPoS3xk+8MQtTZN6b0h
U5AQZcccJUr/wJrlbM6dWq1hyI5D22waxH/sErcCTnEpvSkKaqC9zAzhX3Oy8o7zcIQclBL+rQzA
U3GUEdCujIe/v5tDrMZmr0nhDKKCZQs/xBvL27RNqBY6P7Eh1G1eKRfjc4wDYMR7fcO2WuThiser
/qXU0jwC8wek9SzWLv5hIb+u0TUZS6DEq5DzVW6DVqJiJ4gCUT/4E4txmuqu6e5H5LZ2hrAmjuyc
F/ifFqOdJ+FrAPrWBrBxrq/P5KPg/uZ/EihxiglVRg/F2l2OXJgks7fRqrGLBSLvWfFLSEgwH+/9
Le86iBzPeUbJFk6uBPYYvo2PljgyVWQFSaoBo8GYkknj+hMb7qpt/3b8oKjS+rLIOUiEMQX3cLc8
f/SY6W+jGuL6p08ruzycKR/5TIY57Ko9szoaNIL51OQZFsQekCds/wK4okIt8N11dZnP/4jcLHCL
yAdJimQUMTg17droHNrp9zHDO9jmNz1phZKa0a53n7nGQr3rY85iHWWPnyo9PrOi+PTtqi+MgYgH
AXf9Jk2pCiHsXXXS6qe80cQBdBGibCDrzVVSvubTy/ntNfu4IcmvGZ9VoxndhC95TawYjHl9ybCS
FEtXo5cgmZm9ZYgTu6uY4rKMfdDMxoY/xuiH33TpHdBqnNHpbAg2PB/RxmnnNFIIHiBVpf0cLI0/
3FfYbQNghQ1nZKZCZ2PwNt5VJ4VMWUn5cxqpSxSRaQ8QVK+EOrfCO+MmAsf5LhQo1Xkt81zzhV8C
hQuIhXnlnnoj0HxEha2UjJN5Mux5GxtQpCBpoT4hm0dJ6CdxRIyn5mwwpTbCbKBDHCneQ1oPhJSz
gVk7sdE6TEL+V9Wq7mXbla2xT3CjFxg9UdYjUNdpcQO4IAgTjziXK1mDADqADx//Q1d1B3ZP6nZV
H6oY2pjtW28lfqPdblHc0VE7D0Kx6mDDObz29B3pHdL9jR4R0E61DPJEyO8EdmgWLZUnD74P+uTC
0sl/yUGmTw33l2MZZmtN9qBoW/8OVm2oaWCrelgty2ECZ9YDdQmG0g/m+nLLnTr/XwIQh2PITjw5
RG63YCfi6Km1j+YQJ28YUnu2BnEHj2d58HOy94Ndw8uKqnk4XopwP4bV/QqwJLTG0IcmAvCPrQIc
0QmHEoqeFC5BJusBnkknGIL/9F6V6q48RAXAk3hnw2mW/fDuJMkZkQbcxdsBPEtxWic2hUb/58mH
7xBF/ryB6IyVY6gmXBsrIwE1vNlACL13lpDL2eHlpmXN2XnKZrOyWdgjI4f19E1Q3Xjt1HNJTtuQ
mAODVCCc7geZ8mQVBBRxf3plrRiD8SMkkr1FrZ7o7VUBSkECE3qEUng3oYzOeQtR78XX5LYhwFzt
nuGevLKtBMxmMw53V7AwnS38zODNlsd1+midbIEb8ZpXDRXrMwdGun/wxVfOt9QFEZM/z2KFigRF
0jC6PVRsbnWTYrPy2twgA04gKOWaghK9G0lmey3q+PbhOOX92DU2C5SUmTMKyH3lH/DNN86DFB6J
XYs5B0ri8M0VpSYtc4nBo/j+rZvByRbN+lSB0CWr6Fxsx6hKk9Xd6k91wff6TbCAE+67C2tyoVQT
YZtKSz+DHmBTouWJeqkTIfEpTzLIaLkDhEUixnwACeHIL3mVNmVEpwVSO5cWQefpdQ1XKTym7PdU
IDOQBCmlEDb4JR/5SAu0/uyk045wuruWXNN+/4bkL8/iBr7mxTDatVRWIM0pq9nD6hshA9omMwf5
VzY31pdTEA5i380E+kQhVZfxIcJusL+wCSTYnD5Iz+FFWUdtiG6fhxSqHUdGd1hL1yuhKoi+s1Ig
u8t5wCXjcsP5ATO1taEmZ0RB5MxURQpE3Jxt6xEL8v/o7G8A+wx1U5dRJLenUHRFg6iNw15lGyp+
XvZweFsQjU7K8OaaH4Odz5rq0iw73CTkjzijM9llcxjHw9KdgTOrReSjTeECCdq5dgPZ7mUaF2Zv
cW8cebFK9TtNYvjcQMezr6cRzOgelv1EAgNXUTmmLvQUapPc16q0lO0SoaMg7sYm4/J0Dd/tk1SF
KuT2Oa9RIrSyMOHq+JrHk3A9mAxPlCk1hDAGwFs8KLST6VwmMtMdcnQaBckIU1mYX+1Zm8M1hQts
KJc4t7/hVSSe7uPC0NlqkJ2jF0r2Vs61EvQWm1bXhmA9ZCpB6v/Y+BgasMzKuGAqKu+CRlpMIe+Y
Tc5D8TNNXy/rCKn/omvRtL+Sgfly8DNnxHAnCaUwKrrLpEtxJBz8sHTef+ilgMtH2b0ulnetjEgE
EiTV267ZtqbHOsRqe2RP6NJqaEbtqMBzuweh7ZCxgjPG70zdtWPnN98p54dwcYKGaAfjtRBmTpGt
bh5ZepYA9LCVbjOkpCZO2zpc2mHWcx3EZcywpxBz9a4tlk/S3o1oJLIZA+oLNG6hqlX9psza/+9S
AS7lq3BAHOSgRjTz9JTI5ZvJPZVWo3CYvP4SCImZaDUbEMqT18SABjqlbQnVOT3myGn2Q968zepj
lLeRc2lXxZ9LHFLhkKP5ORmHE83CBaomh8vr4kykiiovNACFqZn/Y5ueWb1eDn+9w33zIZZ9TtmV
Ueq1Pnx+doqv6jJzmtqdOVQxelvuUYPlnZzkVxxNxY7Fgb6fIR0ewKCM4H0niW/YrtvJAjYI/nuO
LA0tyEUCjcFoG9Br7uu6gXDuV/lOS4waqZWpsQTXdOpWDicYrSZvwDNTb5v60YSDKmxkv8GjQROA
Epi9hD/ZHGDYVymXBGCXal+zk5Bw8fNJiVmujuccbLeIRm/UmsSVYmRd/TNY7sq8F5DTJW0DsM82
AVKzI69Q6kfCma1Y6amBDo7Zg0zB+bjcrqloEDHRuxYgp4vu88jD3LdtIEJ0IiiNgv1LkFEeBj0M
shZtuJtcIf+20UQbjN7vGnZArXIkDHnHSqhLhL90oL46NMq5Sy68Gb7VDD73ZCgo9ORIY74KEczM
xGJMHVlH2USjPcuMTZg7QbBcRtRWe8cWdu/dbUuYRIMd0u54lNFckdm9bBGJBYpYfMMei2+H1fPh
W8rdpzEQXOtDGArLqhcfnuuuUmv5q/g5UGVtaj2Y5GU/qTAc/fwbUenYwjpAHey7mGBypbH76OXB
vE+wMUmvX2JP3ZZdHC8Esh7qIhV4Qd99uaa2aEhYLRZytgeG0pjv6PFa292PQcfsQQOxIO11xN0O
cH/2drZltEpWovuZu7DrsxMYfLRoJCpdO1o1RxJx2ZiK//a7c9l8toIXRzVjcfsTQtvktIk0hHlj
ZWHCh+S2XtN/tgEcjcErRENnCiqq+AW3N8OiFGtbV9757eU35sDXny1Ie2x++5LasxdrujvSJL15
Apal/vOvhbdhPkk0NbzY25xosMQ6P6G81byrCAxMMEGNfwumnrl6TwkMW7kjybBB+PeJc4aO4r37
zty0q4IPQ7vqQrgbBmXa3+2DFWCqv5eVt0HnVT0Gpumg7QIyY8ssI/VbtCeV7M2suD40qWJ6SOzZ
kxbrcIK8r2Cu2y2ATeX1XdTSzvd2KgXBpwHvJhmnXgm6v+0j0imPwu6noxprqJU7ts1ygLOFoB+I
FnhcHPQOG9yY2Oo2lOTEnP45jysMRfH4L0//yBzmUjQTQOjBaO5eueSek2ZEdfkfOqK1wyhiyVqI
4S7oymR8l3u+YuY5JDYIE/+rglDMGIJG57rJZ/zeuNlfqTdAQWo6EqFvQErJEhhsihh4g1nt9eo3
WHC3f91T9NZotH36F1g2Xeohth0/60bXXdKhpc3CekPabYvDsysG4J695rNdll7RLZZFX2uIZuFY
BfV/yI3nlE5qBe7S8U0Z0qnOUCq8A+2V6XeO+z9+yFbXar/ruRv883IG043BdWZPFM9ISzUmCIt1
qsu32H0I1OAvxWmaOxCj0bdA+B54sAvD2kcJmTz7pXB5uPwJz0uI5PYclTqrkUxUtPoncMERK+bY
7kgrLhJKXZDMk2ymj92xKavWh0IiDE7k99zdJTI99lym/pbhmlRnsejDdXuwWnDLbPx5F4441eGp
UAby+xOVjOhobjWvVEWxYXXFgsA7wgFL4n2rBxK7D1Yp6Zx3MOmMmjLkKXWnp/v2PMWG1SukKnjE
K91EUxZ5+P6NKHQxBY5tzUILHn/LmODEA6MA0tCZ9RaeyZot7OjHBPQTDxIGgHZ17RRmiqtAnv5k
ec/l+dDvv+hWQPaTCGDdijtEX41VRYBflAzeV6aI/7egA4CbCUQQhr1MTmQwKXRumYzbfTVNVVuH
qAR9yNatfAuM8Z0sNog3ss8JKoRndviYk66QbFMIojHbe/vpf2KsNEgUBWFLcHCYzroZftRFDUht
+jpOnBv4beHXPlEEdmYT8ixhW38riJDbJeJfw4NHPqvgOnBylu+iK993Rpfmkz9NybD+brv8iRyo
uig6+AtpPRjFWtPe+4MVIEnthbniL0sCQhYLAJP3VAj/eME4oPSBp2xPl0sNawhlBnsYiBhQsM9z
V1KgIh5O5CJNA7cKnJOVyDIjPiqmDzeMnm9klPdF96C+cOXQ0SGPJ5RKV5PoA/VAH5ZgZUTtuAp5
rZRbr8LBIPvYGTbkFunVYikmVDubmZm5Ye4fV8XKqcTj2Z6gCx0qNtSc1LTiTa8mg/TlQ2dgheBo
Z3TSqirI9WrRXK2xQPTJRFtTkc89dxH2GQ/p6acLpF10GvHOoehApAFhJqWU2rxIkExm29OLulyG
giG3Rc8f/7y0G3vS5kCIStUXK2DVMmxDRbkrFLpAs/rJZwkgxW/3c707H/O4wbtyNzArU/kW5lT1
r8zLRj1ymE/Jiep5ubFjfV5P6UE9ZC4I7rfkp16OnMlmMgMzljd1hX+XEzWvT9NXMKkpSKCb3yXy
O2S8c9+FLUHkr7CsjxsdAmyus5DcEVmLmdC39hOy9PBAQ9uJbCQ0JoAoOzyeuoGACeQ9KyoCI77k
rhUqr1shozb9fRWWFz+IW/walokycVe5O9mrR/YteqIUtxHAiVIS+t/C08YKIBZ2MX9saCS1qZEJ
XUFmSEBWlsfwpWYUwNvyyHm6ZrI4jqOoDs12dIxrbNVxZsj0wdpyGfPVsx+0csEKXHoH+ztcRMm3
fSiFBOWapdyuLz3sHH/LMgWkF1drXkgpcCOyzoXAX0RbITu4ei1+Hp9aHJWXlRpqNTfxWHn/wfMI
ao/8fyuIzjGP/EAsxxVzwY0bjK/x063QnndbK5OpjtI9H/hXpEFXxZeUcGvdtBUgfXEHgb/d1kEt
Y4L1d3FbZzyDwe55D86/Id2I12h9txui02kdFbmwfWWUVkQ4WEC6dUpgVNLeUwhc7Kf3YRSp/0/u
LUS2kG4x0+j1Te/c1qHQ/EbBhboz41s4TWmGJyDnPL9PsnRGbF3oo/lGpbujCUuN9OdJNV+4fFUu
pY3pmVmlzzsKpVBbLhiQCyI/lkP0jk7tmXCYHtnwVBAFkeGzpG/XKL2iP5JkiPzqUT/7ZcoZoI1n
oEFtddV7xS16AhIC6UyefP+dCpjYIX/DI9CL8syUKcSQuw3rhPTOKaxOjS8roijaVx0zZlSGkQVk
9Tc+FGr8M21qREdCnpEONYFXtMn61YOMiJWso/18L9rThTNMV3pmnKJTmkgPUWBuhn8mQr56tdej
/y1vrMJEAWhxmUpptVzbkcdEPeRyVNe3kJSLOc8Q6nfYSza5kNsWH5gFWBxdsWiQ4vHlUecnFg2o
/Jo765PoEQz7MbMXgeKJ1QQDxhpfj76Q8VOEbtLdgq5H4lNcM+yJiK7YwKGolK+NRCf6yzc49KmH
UdNT1RvwAeb61MwDlpA0L7KVruEDLfzshFmXPZQweYKvkmwfBArEKxxWW+EW6CUWthFgFKGDC9To
YWRPGGU2iUl+eKSwikVBrnzvkiwBM2Y2CHPl4iZUUcQSnkEvvL3kBQeZsoJJonRA2mFda5UR79r6
nnUn8jFrDm788L0TCsLlIxtQDH4iBZrh4+XObulWdcBQtAkce1LU+tg+5xKpQWTvWRuT8f7hV63f
0MqOVWjGO4gMm254W0rbsXZM2W4LnQIk9DecYzNuGx3c/EXDG91lGwLTgC6NCmC0ZJQLjjfyhdi9
6MEQBbGd8JchRoNvkcy1RJGgw+8Y/rpbfaqofSmjmEm3DlrryduTuVFHgV1N0gBScmhAhcnihZ7z
uwfOZR0tB7sPDDHPeyUGYmn+gxLBHEiaAoJoTXj5ojYMcegtHykK8MQzhAeyIcgrJYcNb6Zvcx6P
GuA2UIyMJCGoCQPADFeWvheR4t+CSlnoURRO9h1uD1HIRNxZDchaxex3xAuvFH6QXDCXDa1CGIO4
wnk4xPWWdViwGiFMKW1+HfeG+3ErGFl2N1lB10qpL/h4sJHfvj27ruKyZGlQCo05BsScXEbBLnS+
wh3dlsjjfe+Vc25O0Wz5a0gQPyzqRgpwbSCG/S7knBtCXoysNr7ZRiLqa8Yh3M+bpPtqLyFJr1+1
UfhQX4R2/NlgMxncoz0hgiCvkvhYVf5cG3lS5i7ib1GnlZ9uBLjo5ZzmjMGwYPyhkEm+m91Psxwu
dGWeFK99CQ5pYzAVo8G7TmN38TPwrJLUtq/idBw1UCZXxAxs6LRK+EQK4g32JcsXbARhCRWdbZnW
4p02Kc/7xHkpB1isDIQxUV/CW35Ui0fka79dd/iBtA28fAvP2hXvqv3RPUV2p909JYylbUoM4QJE
+8DECDVhqK2f4dYX2+DcxLRypfpGMvOeGSs7iQmGCD9YVpwOH24cEMua7vjQRNNOXEy7tPOKQ18x
07LqnBftKyrtBHPaDeE7OH3NrK/x3/HUGqcbumW3iDLi7EK4E5avssZun3dzBpwhSq2g7/Jj/oSp
9z9XZczhUTt0yWozMMoAjPb0E77rW4kfpaMPr/PS2bZWY6nkaSW53Q7TkIHYzAsahNgUqdCSg8/2
KtTh4iGBRdU4c8JSQV6fA2NY+s+i71PZrZ652K6/UZyhLKfYGjPmvLham87u/HsKKH3Ys8bbKvLK
2x749hua/lq1Mz+BX74ao0efxAguXql458YgMfNPZBIiMoNUrPTnZdJ/rayvK3BrRo0hzp4PD8jk
Fm9FPGGb4RGN0je5GwIgEauQOKyolMShyItoD/D9TOVfydWJB9Tfc1QYURsRkvYi0vZb4PUwLb7r
yB9x/FZ+JXh2Egj7f038zzH7Fr+Ys6X22MWgA3U1PQuC+OfKUMXD8eVweQAZhxjefegpGh2+o5LN
VDYWlVmKSKWzw6jIvRpDBAvI6vUhR+Ht8EMBrjCW5Pvh8Nmmx3v4gBIvEjS/J08ixtxG/NR/t2YT
hyoXjJ8sBr7MoVF4xt0OcjgxeEzj+WrNoiqPCZXK2e6YMlfcyt3QasLhs6F4GobW9Uiiw1FF/9de
T1bZf6pWAfVP9uTIVFr7Nxd3wXEws2i0u3u812rebLgPI4w+K2s3woU7LBYNRcgXS3kAm1HMLBdw
pTZK4LA6Zmad5IW83ftSA/YnKD5bKLKqFT26Q143HFxfXgcza1WlfmYbDqIYTpcxKdAkXMlAmsqD
g6Z432Z9Jjc8/mYKMm4r9U1XUbRlnygITgEvnjMDirEinMDv9imJ+pgeOIGiaDXOg6DkTWYsMuQW
+TrAlxTDE0dYRgCtQyGanzJWYMPPjxRj6BFkiw8L+6VqxUaJ3nl5zdo+omqHI82j88e7hIbp87CE
BBrtVHYdqezmKi/U4RI4xecRxDkdgV3ZetgUsB5h3MbBBTKvn7kcLa/TL6GLEKs0sMjf4fk8qH2Z
n2dDx/Ji2nQ/5FwGhjQbe6EkNVobLbKA0vzNNBv0eIln8vvWNRTBjXlTknLINuBHvr8IH3xeC/ag
zO3eo2l7Yxm6jyw2k2y2CbzbWXeXP63rdJ4znyNA06RE+wwSwOjvWSvGBgyASiFfPqa/hcDnSoDc
Uu/EpUF3ITllz1RhIWRTzzW4miTKRSjB5IZGjgJJNwgsm1uz5A7ifkMoym5gu6igs8HuF3gh1CWF
2QM1+ciMHebIGlpE6r+9UVsYKA1OjVSyzXVEfOr+WmK0P87EMMW2Cal8grfzpOrARUhWmrsZBIIO
/lnSmOtqcAmFmdNl1OWCaKiotnAyrKS+luAX43103aobuKUUdycAb0Tc/oec6LkzlXhBL7aZzHs+
QjYDoDls4wYHsp9hMJc2FzQw57p9n4zme0l+A1Ddy87vvCytCZsQwjhuxutLu8RaawTHCVqDoNbB
zLeNbHvUBtTDHxdJPl43iiIPKpXVLJdDDrGrCAobvu83lfRsnu4itACOfmHBheOkpkc0CNq7AleD
nI5YcNgo8y7EcMR1+BR8e67Zyk5ggAxJu/aqiGTCKwKD8n/ZTEDWPYGC6tAVwlEQewG9gwB7z52B
j8V+wyzX3TuesxtNzVikGihS1hkphyrvs2AmtWtcsmOkNzGSv5D4gc9rT4KTRao4Li0jh8ZTX0Dk
+dt93dq2nV41h58Dd2b8HmMIAYaafOokF5zag9Qh1obW+pe4hQGUTU9eWWrpDAsJbcMxXFWXy4kH
q1zxbT9f6K+7sEzS4CMBQVZL+3nlasDstyE70y2JEa6VO3DzecNWURHJu8ukdXixJOt1e1HlH+x0
EawGVJ3qVFM+jhxgOqgUZLdJGvM4aLlw9/0i28X7A1mgZDguf0GT7gTiKCr8rJuHWq728eCa62Ia
EINeJdmaLaM57js2Bwsr8y9zBu4Dy6gSNSVJ+OKoNSi1Yty5A7JM6idSG/PBZT6y9wkGmtr2FRRp
7Z5nulxmQgRlVAbAZt5KI7ZsQ18OhxZMqMaIsptKvx6EChiE3q35XEnRlG2TuUvaNSXSCKNyz0GI
15jC2EpU8FHSn3oGeXHQuPNEREvysCpx4cWBolEYnl/F3gXY8d0ctGOY7jj4GtE03FdvgnDeTB7s
iLyWgAn3u13RZxbs8lVV9udHH5D++DEj8YTQx8BYzTUfgcTStBE8oIc+s5Qg/vXBH5TY4gVYJgr4
AFyfvescwCnGeZqmob8dmdBY+wPK+IQKtmfQdVKWaellKMmIXQURbV5EXNpOSJP2MIS41C2aLSIb
n6dDR8NOgj/bpjh3RNYj5/ZddmaKnDtttBh/4ZVpaGL0ZrgP+4ty2sJXgw3lMlNRineHdsC5J8mh
T+RSMcQUso7Nhk024jUlvY9xADEgS1ws9GrwFEm+SVUuugVIQ4cNCklqFALRev/hrIIhOc7sZZAH
oVKxCPrgIoUmkLQXPGeKWMIdUQAfyfR6eXPhOKQ/W7s5ibpkIlbfnHPRakucoTnIjqY7L5zhtebJ
Mb56tRccgh3slUxJbeQFAZU/2h/FlXFJ8oWiyWJtP+sCLJ+RdiNO+A9/hZQ+cWMybqe3RvAxJ8nu
mn+9jJqAOF49FEsHOXSR0JtmxLndYLTGAwGyYggiabDUdowfTNcdOKgTzA4UkSa8XDI0PQTD10qd
S96jtTiMvDVEx1b2AXlfWxkl0iX4Tzn4OKJRpqVwP+ksC/v4HR1HzOUzxsvFyabees67t/cmGt4F
Zr2I12NxZqrF5hCs69wv7DtcjOCgrmLX/MxI3qrp8T3fvBB/yoVpUBs8Kh9HBDxxc0x9y9H7wEWA
sFPs34+PZxvUqI617j2kSlHaP/6Y5/ACOIn76l8v3tK91XalOwY0qUuknYSvOyOQIjrq8SoKvznR
LaJqlcGMkv+MityJLjEdqCswiaLGed/PFOakJlLiHMZvt//MukEw02jsyjwAB842dcbM4qV3QRck
cTyGM7aPm3sXe7v+RwqroAS/jq41VxpfHnm92Zit1uxLJUzMvkLHUfWjA2UUGFJjrzmEBcHkL5NR
yyJdM/MGEp/C/3V//4wDyQDaM6xO08kwcyIfZ2ZhNPQB9K6MXSs3wYiPzOYT0yq7xVagKKWDgdVU
40DMM16Z7EJNs9h+NpQAKOwY6Zod5YeywZXinIIKodDkp/o6AlGj0tIKKwOE9zrdaLSoBXk0Tpe2
jeqaseTUjIYgfugr0DY5zx3rT8he8t6wIxQQmU+msiSricuxQKjOBEKrZVCe49a38AusliZnvtwM
V9KLqQ9gQfDSNWYngKiseRVvKLnv0lP2COH8CoGeRpPcLx8/PXGeLGMhb0sVsWWwCx/KQxGYsNLI
iyZjDlJaDl+NbtpS5yhqkQab9Ck0lZm5FdAc3Xj1YWRa4nT2iqpJg3aPh+wg/KDhCBu+S1XT4/eE
2X6/o3FxZAoCxV82P0dK1DlLP4s3W2jfbQBtxoUrfx5Ap30TrGo7PPzsu4/PqfWHGA+laVlB95pd
nJtOAHfhP/oM62NWh4+EiYn0gSXlK+a6sxs7JyPYNP5YFSJy8MHnX8O05s3RSgxCFwmspG3rlq5q
gjkypvRR1yy8uKUAjmMdD10ICvXoHCZJbtkoiyBRkNKCd4USqqb+b6/yceiM/Np1k8hIUmIvJdf/
SbSvb7pMj2DnW0bnX8anTJiiqix6YjnDG9NJcLhjCr0ydLlKr6Gm+3U02KjICenQj3IK3MtKQbQW
3+3elxBsQXcOf05vf/bcR5oTTaABfhosHEzH3WCqy9/Q5b4nBJVT2zVI4Rh77pCkrjMKdZxjKdOf
NrQhk6juHesRVvBIeI8p4e+VqhSbmYc+s9aCka0EdgWQOGkHTpDqoh2RpNhYfjc0QZjwSKK/Vidn
RYK1d5mQGQkj103cujjwGs+Hs+VADYSgT93/tkcj2jVM1p05xrt74Am6nL/mQYVmdXjLJUYDhdm9
JV8iAwVaq1ArdThjao6S0dY6yb9x5stETd6mEAgcARJU3Gnm5iiCJ1ga6j0nnjWvO4/7sSnP0neq
omy4QSeWVh2SOTyVk6QJte4MsADGk7zqZ3iLXsP2RuzwWbXSYJWeK7bldkkxvX785uQwxRrfCByv
nky5KZfuWfiYzttYA0GybrUy6+P9Hk/A5Mp8FznyfDkz+qfndhvdXdwvxosk2tFvRRxPDx4bGn1T
IS9+tQ96OCBSxfzd1ICtYjOer0Xb/gSmMhmRdw+sGYKHu8ze+wBfUQkcz5TWypZ81ENnaNVvErH8
8MCPfpszmHqbdnVi4rk5q2YYi45BFKBz7VoHPvQ8unU1/17RNndfE+O/GS0PFNDNv4IIaU9jNUFH
vxbDF4Wufm71KIeG9TPw8deKtLZ/3DsHE75IZVPG+KMl8cvfb+H6zC/LbUCbGyDBplHtJQmEd+jn
ySkYyco/xjJ++famq9yqX8psO4qtUZNmuuHS+5Nl7XqSjn2seUQx62XtJBiPoRtK1Ilq6NjU/Pd3
uvjm1VSUQjjt2+CeXNIAZkrZFj2I7hNDcecgeyKl/QrSbVyxQQPdjOUaTz0VNPFdei+9XRSC2INS
UMmfKMloW3+kQ8sy+ysiIN5YC9XFxnPEYzZE13Pni3JOoTOLioGg2aUf1cV31NjTyEYysyGXetJ2
RTf0EhL1DK9kJSz0YEFsGn/nTSeaMd5pW5PdHMe6d5zUfPtb6M288PVit1906K0nMyey3P+t7aC5
PknchRpbPpqAnwvGzTlgAGUzt0X8Js7sQAdSTPoLVMZUlbYiC9dYHSo8I9ZN0s9WkhRAgQv2GEaY
TCD7Zvh5eNd9CSVV6AkRIfGkKT7N1Ei8wQLAkrldMHm3bQETC2OWwmZxlufkOAQKAi2uRv5RSYFS
85+Y5J+jIrlgy3ScZppfivPOcWlvfSxip6F06NmTqhSwvbj5xek37+z8bcPkpMzCdOuthnRYmfuB
z7KDO8g8glt2biJrd6yHfz3THV78MeYr9rXCp0W/PVL/KNyFPlQhmb39L6VdgCS2dqJbj0vKnoJd
/p/1ZfXKiCwXGILX2r/s1FHt3vXpoFoqSTkqOBVQnvcrSL0wvZlzidCXb5Jt+j6rELRanQp6C5oF
roBmJEh831x8jbaQBOgFK3aTFlv8ES2gkh1tte8Boe816lnsT+hjfxRxnefYvzP7OxiP/BMq069P
88YOA5Ul8aJlQ9DYzDeZJUMp74Kxi6i1sjsSZOigqFKuMZl9Scqc3C2Udpko0ckGblhWXPjx5LCM
uDQ08dTLdcoI99iwuYuQeYT+k2+7nCZNoDQtLJKPC+ZYD5RJLATuZSYG3SGkZEA4ia+5VWEVXYtH
Qd8QFpVZXNEjyw7QJMJ5006L7kwLwqmNB9i/fxU3nMUorlH+ltu4Sb9xtvuL/cUbiVO3MyKU2aYT
YGyGaRzTNdjKSrFex1OEGUsTBpsxUXlss+xJzPm859KLPxQamMHgLUpuSB4A9yz4+hdXrQep82KX
vthkFeQ7tS4HYfMbeOLZ9YxtwHbDUtiBOgHYHqcmMRQlvYIxOP/aa1SGsHggO4z/qXtz+v4mk3m4
Yi2pQKYzVkQTUuz1eIAvdfVDt3tAOK3rJsRVtOeMT+IrY9OoVaRIzbpHVidgV5lORA5oh8N2eD6O
jR7ycRD2fnK7ILVz1OddsZgxb3Ph0HBdpOyFzncQ6N67Ye73vMlg7K58NbrYEyUpchCCKzvR6C+l
F8363C6fAXGvhuW/SfQU/Xj20K0awBzbKo8EoQVt+3Pu0XYxtxipVZf2Yyc8fbJcwpnHfYSPVQhq
LFLDZE+SEC86Q7ZLq7VZutAygDRTT+wOAVpL7+GVVQM3tfGUxqkos9P0CStrzzv0o0Fp0066NjIa
eO7fDn0zfo5+VlR4RXZR9bhC+ajT5v96j4oni9YpdCzJZ6kt/FMdavgq2NTLGUkxQ44RBDwebvYi
Z2ZjrGPZz7BCW6hwUBw/GHF9y2Yed+hsS6UKGCVRQLmTZzkhBOR5uq8XKJmO2Yy2f4StRvtjMbhX
/98a1XNmMzNgOx6qJM+XsMVGxx3RRD81rtR+5/cUP1b09/fAq7LacJpf6x7pCGjWj1T7ODDPkWew
1wSFB+qrCwSpcs4bCc1bkO70qSCWihchTxGu2MhzV1nW9dhpGKDFqmqBDG3zM4XaX4RlsA4oxWEJ
hTiRWwyFkmwDBXoPvqOn3UGFGStVkIDg7iFBC4AerYhWxXWB5YsU2hvXl988KTcM0Ru0x1AYuSX4
QhJhUkhHXPpylwHhWa+yedymkynL7VeW2cRKYxxQ0+etIv1r83M7/yNqPQUHT8xRJmtoqSS+jFv8
8Cobhel4r95Iz+90ksDSF640UxetuxNxSNDbabiLQ3eTF2TV3npY/WjOGGRH3+72pbkAkpAGu0zv
Ys5BllplMUIrk62F3noJVFufdny+n3hsvpjSRdt9fb8oepNraUbcZ3WxIOnva3ndHCsbWYhPiEGv
mjxoUFDrB+H2nkY96UYuc2NiUmS0udR4x4PJoLYyX2snaoWyBfS9mF5SydL+coj6/u6qlU281ozu
eAT7mc1O4zzBobxyzwyLlINjNv801rMeT7flO6XKxW/x8vJ9ZYOCpdhUXG2HLk3nJ9IZHfzdI63O
Qr42sXYpNnnDXiouwtcpJGWXREQFu/ukKV/IpJwb2vzdcLrW0MQj9/pLYsOCNqj4XvqMCc6p7qi+
OJDiZA7ZSh3gI6UStLEHlw768OiP17iqsVAsdU/z+V5JGyivDR3e8tsW7YofAnlpmrkxXRiXnulq
Y/i7CuRK7OsmVggp4bn2/BaXlwUNbNe3jx2vqhL0NdN331pS4hsoyv7Bsd6nDTwJAjArM1+E9dVX
W1EgFC2CFmkJZYaor4cBDGe+zL/7cPQSxe7fV61hW3wKHl7h9mSo/xaE+yxvDKGUCR/3ibWzLH1T
AUwZa87yNQ6s5GuUGeVgibVDelfC+QnMR9+z7O1MN1xrU5oi2hCZslC508W0SJeqRWqCN3V7XVP0
4TNhre2ljdaqGKUq1vk8EN404f3XTnThx9+vRpP3GGrtqrsgueLeymDNEHjCZZC7ZWAZk1THit4d
I858FLzSiOnTXPHhLZiWPvaOT+NJcMU9f6pgyhsJKiZW+XC/MTmYhd3OiutN1Qd+dK5SLAYlW6tn
iO6UGWGOMzrqqZ0za91X/T0VuJUxR/OQX8e+uMEz5cyNR0aw3iiLG62LejBRLiuohS04//jX1HbZ
Q61Luj4S0qpn9VchTqnpgkKYcVa4hAQ9w/P4Qiw0c3hOODpcRIeEEKJJJBJRf5se9RJhSzVOEiTI
9r5I6f99OXTBPeQqc/mq9I5XKu5MRQl4hOJcNh/CnpDN44RMcK3YTGQnM1CCUae8xTrVyGsYg13r
RjzxmG5a+xJQaSwR7MoPGDKvD1VVXs4jvCpL/jO+fiiqRDhl/uhtPHgBaQPILE6bVPpTg2rrN0Om
jsr9De6FvA7nb6O4Ud9ja5xKFHUDM/mbNyfU0MwoBFNY535PWECuTHUdkEiv/3Tpm4bKGw8H0yNM
/D2fj6wZ1voWktyr4f36cS6Bu2+sU6MKg3MBso0x52QEt9YzpNXvms8sCo2haDfQIP6JmWM2lMpo
62ejzHUyrmw9fOg1kMcI9UQ9aNzoOLXsJqQrWV5qhxnzZfy/UNwochR1G0pb9BKyOc55q8z0WiUf
p3CjFOhe9zhsm/8D/QC+T3vgBXUY8wZe0SmUi/T8vEXjlRfdI3suDy3hsuOfLrgaL9r8z1iU1FFj
wZZuRVVxS9Nu7RGP9sypxIaVLYJWR1OETDP9Fu1N2Tq/fBlRa3ywrw4N4QpSMylbIAfwqn+6g9iF
ZriGKS69Yqn2W698WGp3hZlHg7T9QzWvus9piEESLNvHfz4sJeXF3gUV3bnYpmn/LCcIf5Dl5VpR
8l8rvHX/0zBh2ZgZa/rf6gnRgq772rXasiHkupemHXFBwcvIvOQoWqNFYdA2NzqRUQXXkOegqZ/1
FR2thP2QbRytpLFYdJcBVyiJqCqJsetSXBxqfZ2aKXy2/DUaHSb+LHxvul/Y1OQpNz37TuCVm1ij
CRiM9lWr9ObfH3if5+0S4F6PLiH9dWZQnv1Xf6tsOm2zBq2DRQotOJxllJ4Xf+ExSJXUKhlGvaYq
TRisI3DMYnT5D0EBh7ZFrcKXplkRW96ebnA0Rddum3HogtJPWiRudpJLXHOEBa0oyxUkRcQBT9AI
eTMbd5nU3NTxe7blZuTTvR8wbAl/zY/JE5M2Z99A+R3hSsb+WW7h8BiwJsHLectxLmBpIa/C3rZu
HFt+eiN0SmA25zg1Oa75kCkHZ9NOkJb2Y4v8rholIgIUqeQanWSjvuqQt2f/6zrky8XNPWvDaJkU
nQC4+sHlGOM0UCwMHJ/7lHxyKzid4yymNMsYGeXEXA+XRqSSe3IL5z7SBsm+zowgL9XeUogPuXN5
WE7n3VZ6ILD/9gEXc6+upbvGsRVFtjvciakpQgYAX3pKyRoYAeppH04KRzaZI7iGJ0uvkkEw39Te
EZWkNcMTtc7p8/w7uq25w6ym+YD22AzdvHA4LT+cXLywTYx7zVNuBFDsp7BxKqNj7NBKuF4O9DUD
zWjyR6brLMv/hose0kg/andrjbCG+vgFNpt+Fbnsekn5euJXZVXs0y0gwQy3+4lSuzZMkqWYSGAC
+mZf8IAwtKja+8kuFLSIt3XRh3tee3zhRVwpoOPsPmJG9UN9WvPYVBOxEFCP7JfZfImkNpEngBoh
EBcv43DrD4itDp/V2BwLzuhBSYox3MlWn4QqnOwXUWxZ/yGNo35jdDdcVFmI5eM0lzP/K2lTFFmK
m4QVWs0QRtf/ClWZ1HRnVIT/r6CKTbFSt0EjhYZ70LG9PGDZQHfAwrKbojuBi+XkknEw9sp076ox
AEhVMUvOvKshEZaHQKwPsyJP9l38WryXMNofKx4Ciq6Od21QXmv3pmb3wiI0Ke1DsumOYydhqEn2
9R9wQZHYM0KBljMolfuQESENRzhU+KtOMVxrYa+Eepht8PJRUZHR1roD68SH+POLjzdRg0+5UfU3
Wn9MgNk+TZOwef54LRKaUa0ttG0cXsZz7iWpmWJeiqEldtSX4OeAAz8EBHe7TEmt9taDZHkjjwZL
Km9bVlDzGBlqp+gjaxunUQ25r/bo1oErn8XUFdClM4eq+FImq4EMCtkhXAm38JUUZPu/jSdu5BKC
p0fAEQIe95cr37y1/qAzj6l2KTskjpuq4+fiif6osuDFTVZOyL7YRfkIBzUyxTwW/uw5EiTNfKzR
3TedlXwvVMjfWftxyIjfkJDIk/VQRK9r5fHWn2L+T3LfPwvIHrHN2THAWvueXfgBKSp/OO36AeJv
0m5loLm3LvzbUs6feJxpCwd9Q6NLoo0QR+pdYPThR4ZPtAfqwalHrhBYau3QxhkdPhkt+k+dVcUA
GUN7i4i5tuIwdGOGxQ78ChPFD4jOlPygOm+4xL5306wcdntJFhAuHiIlOCnzlbvfZm850IcHnJIK
grXBReYdlMHUq3xVv39GS+rW/K13w7odqC577D7EzyQ2m+7CnU6OUZI5a4LYhdrIjHr0NzPgEZLc
RgMhrzYuSBzYbBJ5v+qiH4JGLpiSbkxFhGZqfh7LhXOJBudBkODIKBF4pZJ66vdA3RFD0qKQXClF
FovMy5cHJ7JWYPgChzTcCJhZmgR3zQoweAuEgUDui4BZpO+86XpW6mt42NrYFRew6j42nvR66kH/
fLMqerEyDKNX764ZY6Ug4EVhtL5K7WhmeHpuHCkADCHBHwGubushLaeO/PK+XKxGr45XcGzWghb1
Eb2QgfzY0IBBbpwiNm/c7qGDbB1xUYsiZ7Kuxxi24uSsbDrbGn4v5m6Cn7SQVZCGUVDAW+33c+4y
aQGa4S8QoJUexvTnx5nmJFBNjE5QNT3qWfvCDmHLGy/1UBXzUs0hiJwy4zJnxZFIUB8TlPNOaKrX
mZ/Pwk49QFu9RNx87r9x6CIFwN7WiKLxkOIm2VjUUv4BywVLHDKVOuakc/o0ujnLmlTwcEO1f1cL
YJI/hGFKUN7bRlOVJaVYEB22SGiua/Zw45NjQf4gir5QJeEz7TBt2qZzoflgO0w/5ObAMHZVb719
1LERhcjGZyFRTFcZpN68zMsroXu0V2Hp2mQ6GBoCTXEQV/25LPGJhOZrIKhNM/jA7tozjoG0vC8t
AdZn0PAEiefkeG/H6DHdqU/hUY1VUxBvPzkSVcKRrXSfsJLRvvXEfmLqAn1zP7aa4CRTXDLIxDJe
QbWjdiU4wJzw0POkF+6xNRlC/Nkr+GNnU9tqFI746K/p3oFo6x0bYtUgZryoycsFW/A9VCGXR3JE
sRsdqOAmOdyFHzh5Py+YH+PJLTu2gW0zpyYsje5/+pxQQbIBKrSxeoTF/dt2VtJBBsaKuDT3Zq/O
BvWoH1FdkLY2LuIVN6LED8Lo06lOWLHVLpAJr5wshNvLIS5pxfKzoLxrsFxf9PuxZLmLfmewqaS8
kDWmCvmBGudiUdkM/AfvzaY/zkXpOLlsl8xgb1yaJjpYq5zB2oIrPcRT7nGlerQ5Pgm27sPo4SIK
LThEifkSL0lfRITf8wS0ht0Ul8g8AVRMH+iQqDuwtxXAfeR/teRb4Eo8AZgDrGy4djpi+F124hhH
Ln3hULu3JIiwW2anD7tWjAljFoY62ppTbDJ9UoW+YYOaOzjC5Z9BawZiriYOssZ5CP5ksj8dGoo8
pyM4ATDQi6JWJEOiEOglG0b2RCfoSn7n4hyw34wnMtUst2J3c2R9QLXbuO9TaRgnyKv6JPRu14Z3
x86wQf4saguNhQU3iH7gB2Q8Tr9KNPcBeD7wfj7dXIJcY+L+yIiKXZs8wk9PWyVJJvkoD7Rg5v49
ZNWJBxKNMcA5NIcEPWpHaGdJ806XpopLR+e0U9cgAJK3CoVYcFf6BlypNTI4EeUxApnNvfN/J2Gv
S+3VxF1Bd9pSDn2FdeHVzdvH9SFaMCUuHl2ixF+Vpy6CLq2VuuQDfMFmHqGGAiuFtULc+F3WoW6M
ARsZpmCdjZK+lZxLubHiLFbUF+Fv4UCH6ZTXdNsTFW25gZXUxhemPNFyOSi8nUOGiVxZPylpTRUN
sWNW3qQpACQMV+CvhoMZxlX1eZvvGAzA8M8TU5Drm7JVV38TTS3cqybWN5OBrwwFCLrDwo8QAVrO
VUA9Yopnkw1z339gTvlcGKXcybEbaR5KIavGmX5yR3qNNlEgRrdzwv1BCdBrzh5lJ+3WOq2a0s0o
dUvAzje82VczHP6b3EXcoeLpdEtZEykTQl7ZOjc3QA5CJYHA1B2NNeN0FWtfi0iKiJmIzaGUbtEN
c502G6b7DEe+7UdqjOaxKK/h+hH5CypmnKZUCmqJCiWPMrHq2l24KLFjU5Zo6UuXhZH1Rn/ydbpg
9b5CQ7b8IwZJ0r5qXk8X6qHIBJb2jD6LK0vB0t8vANaT+2/hnxtqlGLH+T23GTLE7pHr3GIBAZWG
q5QYYPHAbn7WhKQaizeJwld+q9skjbfNwHAqgNoeU2SIlpe9x3QJuQUIlBy3aYGxvREe95sAitDG
nGvxYnYghdqQj8C5pNLUrCEBMITHR8T7vVZPM9GbQ9oTbb10d6dLQw0MRFdbI7sdC2TF0jvN0EJ3
wfllrQH/gJU70QWkOFO0MmhNN4CZAjCKjmxtCKTh4WJVp+DAqB+5HP6G1yEcvBU9hde8Y9ykSPRl
TFgQ2LXS8El/xgMOzGJvvFs7IZXEO2tguNO40x/NyV3UiYJHSH4JzhWLI3TESlwg/TcphTW2CcC2
ODKsTJKanqMsmwxBfug+rHm3IX3ov8uhMlkerXHqy9N16uM4GHhLbt1AdSau6AwDV/vAGOzQCVf6
7yPZHWK5GrHqLWOnAlDlQE0WV2UQzblsgeJNUlW4bZS+QVFhfy5YcJepCZXPsEzsRmN0ZGb+LBk+
CCD5EeA/HZfldMJj9YqBIkiSAErsrYXZqvAF8aU4AS/N7o6HJ3bUhykOYak9T6oSFjMb4VAtOcIm
KYwdQYXIOo1tnW4G6//9VdWuHz04uI2ifDQcAC/KQjf/N9tT/8f2rsjkx+RXsG1n0qc11IgFyxJy
r9pIJIsgvCUt3ykJ399JQ2y2VxI3NJoULxAIjfFvfifk+16xZf+VLfdbXw+WpYvXOi1U8/RODgUs
TFEDIDohhQvpslpRmsM4ywk54JW6nIF06rUS2iKXkF3EIMgbpzZOEDTeFWpeFNREMwW2gznF+eZT
HOdpIZUtk3z3c7GARb7qA9nnFswdl/hrXl7UMcOSCGCl0FkzBxaUHkmPS+MPclzOPB3W/VBGOmAo
4epToSVQfy2pvknNBVXPCmF4cgh+ZYvJRqIsl8pR0vao7fix6kzNkMUyM0zwKAmVRCWe3jbiw5FJ
lhP8n+vvO/3JyL3mHlkLS+/45X6G4zMoC6fN2NRZdjjGcpdVldwwZxzQuKhciYokianyoC1ApQ2S
S3de6L2mFLXK8jaMVH80z3ls7cfvHxN4TFvLpmDVhsAUPEdHo3QLzaoCkyGlRtje0ZmVUJMqPAUj
0Z5ris+oysQu19+ByGj7YXoIV31ukO2Gz2lTPyDj531EOmw5O6NXQR3+LjFA+WBimOoXs36ZyYL0
l4LhnCeuVGJuHzF5tXKGSTFZpAXiAEIdJUBQPflgwWVBaNdKUpipYP6NmxO17tKfJwzPmwX9CKWP
IYLXDNP8Ev73k5sEWY5///AMeaRV2jJ/hNFyR9lebR2IRmzYJVNGZ4qziz7LEUihU0tu38ANn10J
wW2TV5/bLuBqz6pDCpiDOBrxtM3VCD0SWfcxwUW9nzKazUGGX0xEAgstJsziDRKZonsc76DgHFyc
uzKVrnhxdn8Tol4A9SQMmjPsaEtrcO8oE74ZDE+gj5GHtI3ZtVed7xXMNQtxGCn22eV5vZPS0XXp
DeHvL25p2z1ydPSPG7pLrxgCOk/kF1VUgjRJSRHmH/yiMRrc0pFTVfE6LYsTCatTe3fvQKXVtYgk
xEGRNN71qn1m8zYx9fZ58ijJR3Yz0ygntNsjIBCdh+OxZ0D6Pddp2242VITMIOqlIl9Yd9lp/PgE
dOyz9YW94O1FbJzFewg385nsLGpg3YrwCOHTcjk4SWpRvvs/n03w+AKMlblq51OfvA/8HFJUGnBB
GgYg23VU2ELYI4r4IENnMhBOwg5TBpdjaV1MOUtYUAAAjs0ocNAI12IzrtT72YPohKmXMjq83cyV
N+45q2zRNqx7PkH7VeX8J8TDdHgvrz8LNdvHFpRKHR8MofbMz4lbiI7hCZS8uu0oZVtcV8CROeuA
QQYxyLcm85xAfbAC/XuBgBAuZWbijTevrnwgE/HLIKMSpt1oQ1ecHcJBuRGI3xgI0GgNM1tvE+qu
C1559kIgBydYH+BLRoecfUhpkVL7FavSCHkhryHBofPXheKrqnVI1mCKrxbSCc/rmZ9nHDobV7Fo
n5/YkhfsoRNuX24A2G8IctnzUibj+Jv4McwHPqLDfLe8824cz/Ka/9Bk8fzVACg6e4Xx7lhm7S5o
f1vmd1H3s9MlJE04ueAFmcBM0T7JgKDAlKuXY1Hyidpz4OeV9RCTRN72+w+eZp1+7rmqMlBKvznq
YqRYgCc9FOloXLipn/yC2ezaiIVRn41jCn6bDvGuMg6oeI5Ih8q7rJtg0HqvIXkPK7BaBDWY0i5H
N9UKEAwRmAHrLaaYeF+4/dbhfocyKgOwc5wlIX0ivfQcB5GwYItaurPmpVMVEooSqOSDOupFC15l
KjL8yy9JlAW6dJcWG5ZtW7DzWiRVSMSCcfaQvbmv85Upr+s52HNSKbW7WEw2eI9Bq6MeH/cQ+DSw
3McgvSikySCaNuIsooA0RoDfMDVgMmZ4EN2BL2w9OuCFgOLWbIAO0VwaBNuILL1WMyP6qKwRc39I
A3axCK6eeLqlWa1l/zAW9/Aa03iep+qYX2ENwTKCd43BctCMrsfwmjZSXFOqOVwbc331/q/HXKAA
b3ejnOLNxAGqfqlF+nYJM8t5XcucQT0hAkxNd/Aupg5vHBcZvDk3EU0zuBANNxWI+5WQ1iOPuw0U
Tu1DdbXFRQBedc3AgBxGO5kn0nV36K1c1NDgwQ+UsYx/iKPRrXtwCt0dL93dtSROvqxenga/p/DM
IbBRTzgvck7vdzuJkXYeow4phkZm8n7kdPabfy/VIWt1dunwrbzMt1xVMgF60CSjJu1wbUHGOQuL
CJlaMy56hyAyofjVyyA6W+c4r/vqJoZd0o3MGHq0cPk+6Hkika/bzeRtFJtkE55zEu0THmDZKxO5
PMlDiQ33gX/D8mWq+xvMh3oxdwMKKs+4RK6gWQwGMitVtdtJgKNAEYJchhtFtPU8IzBy0IT/0Gj8
g/HJaP4teckoClkmHyk+Q1rxfd6pVG3c4eVIZnEniB18vDtj6fsMbf+cFAC9SS3d7DZb8uj6mjJ3
/O+e7XSZL7FeHcjfw2XxM5ShulQU8gdQKvD/jyGvGzJMO6xyq3To/uKKWaPcikYceV8afsLn992R
VTFwYIoHegVzPL5zCbJDaNwsqghK7TUP3xoi2g+C1ueaU4TSgJDRCrp3XcVJ7dc23IqIaUPYQ0dF
iIJM/sc6V5bgtgfYQC4sL3l2jnHzULfqvDrVnW2dPMU1SwpKYurN8l/3VjZfutoPBgtQbLW2j4JN
4p/qdAHxXIpO/UnHUOs0s+mWN13UVUMhUYxse1tHwAKJwrMnJ3vnpD0QKdTzsFrIYnqN0iPehqsO
WWr8Y7toxWTiHfcOcYhSTv2Q4/LYhpKKXT0ngbuEiBhQgFYyuo5UbL1YP0rOIS/JQwMQNTTN7nFg
3ICkEQ3AExUCk/IUwy73+GW2sLSbNTKb5l6d/YcM0srYxD7BRz2q01tQLMfehw4Tr5pSr4/MqX2d
tiaFfYEBkRDyHjVkAqWwyU9NJVYoAP3V6i/lypRBPddI7SmNFlVsdlZpFlMO3zXcOfRAppTtTkZT
mB/LwEInAiZx80dqpV+ySoO8mp9+ESz7CXvuxDGsMeYN7Oz814vlx7sZ6kKlN6xGCcxRWtlfpejh
LRRnUn6+qjZu+CVoL7ITN0u5Ubnzqrihlvywc5vzWLPqd+oxyBMJnKWfwkVPnbJ16TZCN5dI3nYW
Pldow/v53jSFG6zEfOFZAneH0VJ/5KW63MxBHmj9XHFoWkvEG6lxAT3UjBapkuLJY4TACj3bwc88
iJyUkbdidtsXuIJtZZQU8ZnKgtx8rOqlhYwMCfS0VIRa+YMFM7LMCwe36HM4KXQ+q5hegk7XkVLx
zWamg2fDS9Sln8EMl8c9V0xAmqsPISGMaSJn/XDAxlj0j8cJ7Byq3vIMV5RA8ShAaChMUdXKueDl
d6pLnl7rKQDxLny0kSMsbYjXuD9YWF516yypq0rbr8YbklrB0w2F8myXC8k+v4WkBJ8bwOl/NRI2
0DLYwSXQKMK+ff8V6SPjVdMYL/JJoo/Xz0wFAzCp9H4rZ7LkEvxjduCiH4wUDq+Ym+4howSLvmBI
8Cyer8upQ9Y8kY8QNJvoq1EZ4IYSFAtQisK5VbJ6PQDR+0JcMBCPVxyWYglnfT2br9E9upeXW8K9
waJpNYX8G/B4FiS3VcA9+03mK4LZ++uEFnwbecPwGMFeRvqGRk5TVDcMbFCLc3spw4DsUirgs2pl
z/JGGk+x0yah7BnMU78gUF/+v1ZEGkkWhf0HYwaAukC5wnpwr/SKYLpkEJFwQSqEAZsyG+m+SVFb
/Hlxj0Wd+8uOT3NUBBYSt0WpabfRajeXdvsDduCsdBAnJNY1KByHxr3AhLjindZ8t8c2VFQHShOA
IKNUutKwkeK2WpsLZB0fHRraC8353j2Zo0mJvlYi5oxVDmsqKCTXnJqbGWMf2VSrz0Ww3Momv5jG
VOex7PMOpkJQwv2Zms/AUtc9yQVuRiYUZW4HWNXkanLE0FGupuxBugNXo1VmfIBWRnFjMiVAx4vT
5tv9rCckY7z2q5QBCDcMwiXz5Bdl/68QtsYcFLEPde+VZzq9+6HLmeNaz7dEzNyae3GxZVSibt4X
QqA7W3UqnI3x2zFZ668YHgJC8qmHD7moJSkBg/a7A3Eckc41EAsloU8+JSBg6Mb7MzkvhwmTeIvI
jwhG4yNRC8egWmJJFiVawAGgJA5zBoSXa8CvYf/iEUzMpIUDbUcuCqICbI8dc8XBijQDmlX6/JPi
liKziuZBE+G54Ybm4ccJpqDGSDUdQmg7ONnbodPKOoCkihFCChvvzI0gK1I2VWvJJHPQmK2e2J3r
E1YIHw5jAmBYmJ0UO1wJghJpyxAaDAWt9dTIUhbsDtfcByJqIEL+EIqAMoDcHThuHKSV6xrid9rD
Yuz2zn/zySDOH4XbLAGk02LoZ4X3WFv6iTLax9XYO41M6njr/eMONtIoWYx+zUvD9ncaCjw8LmYL
rotNsLHPUn1bJRkveRpPJQpYrguJA5EDBDwHvWbaxZWQ5I6/Dmr8ncsA5NMoQrOIxRATx9x2SZ7J
ejsqi6PJQtxx6VrhL0BGCLTenSaNynDyEexfVkaLP5TSR52RQDkjsF/U73txXW9EHm3QnA4kxuQq
1sgVbj81/+FUTIrElhJME+979SjYM9IFRdI4SmqRZSFhxal4vXWlla5Lv2wpR5FYWMBIkCdVAKGK
mTljmjU8nCUcaZIYwgpg+ni9Ubs8SMAUSat0n+jSXwClArWcE0zTNV4PpzHqtjtMRGAgOa23HBqj
kRN7gRFp9CjNI1U5qm4EL0lVE3XSZm//tkvge5Lp1sblSxDz7uaCIRkLYqukbeg5cYBNWM37sUbi
TIOirGjnNAINc8uPt6JWMtaAydIx4NMEHOuEA0qG4ORfrHr2IvENaI2TBQPGZGPiQBRuSWZllo20
2pK1ajqijxi02zS2rBo7o6JC5D5R/iFlpG7d4vxQLRI27lUnKrHzstDkLXB5ZfarwsXt8yJT/EQD
WNYVKaLh4ffxxPI7h69PFh84mqwnX5UziOLOglY1QdWWL81hjCntmMrkkag9p2RHsY06jhFMosOD
lE6qKCkKCRxM8XDBXBylz6D/1+5KUayF+utdX8MjSFb8fh19L15jnZn3fKCiZkR4okS1nz0EkJCp
mk6AX99YNYJgb9Q3JyvjZNV3tjst0sSRWmmtjNGq2UwhW1V8y+pJisumywoxf/CRk19bemnz351U
Hh0Vd8AI7Xj4DswAA1cvajO5VeDCGNh5YEMtuDmbCm/BTYpzymjg4cbekwwRBFA9kucY7TuwJjag
Njcr2vqH0Y2anjP5uSygJnN/VA+uMD2DRG0e99Su4RPthe5S82YmwYA2xCnPmQzYFlOWUickAQA4
KbD8UXfAzO4Rp2yTN70Gw9+R9PARuF/A4rATa6SEagkGXIhvQLG087Y275BihEpnLhSUHsfVaPFZ
so59efAv2KIEbuIn8ZArtAPQylAwUUEVko13KkTmZI4s+tTJQ30f6yx+MV7OCbx41+i+jdTYKL7M
Q8WfB22EHR27h9yH/ZDdUfzdT+/u7b5LnfcO7oHx2c2DXFK9EcMDu0EMh7LACt+qBkic4oe18dHx
lq2t2wpmbgr0nZ+6BGmxwC4WimUCTkCch4XxrA0oGZem01IinYedJO1Om2tKh1LQH4x3mEUOU5v7
lOnzDYAxpyUT9moIp1u/Cghv/oENznkSxLIwKxKReK7EbvfdzJQ9OTR6e9rhxkGFzKJBAE8B9JeH
EjlAdYs72HN1VbO/e3ZHWxZs+TCYQJ2IlVGErwZr0mSA5gV5JibvFLPFASMZ2J9P5Snglqf7ofUT
UaYZhbiAepRvckA39JvdeujQLZvTAikWmaHoKtPNm2GdxK0D42qOhx+pLsW9FOdBNJTWAnhCLIPQ
6r2u7iYUk6Ih/BysyWe+1IENNZ9kZGv2DTFhrWilej3902uM4KXzee7L7FUcVZB/R6R3U3looehy
vRSjQyfLIMgyZvCJSOsm15l+RG5GbB9RIaNtB8J5UTRz/PwLjgzOqWyxGY6+g6rIU0SLhNbZO7GL
+c/BG2o/DV6jzgus+x72CHiw5kvg3ClwvEdFRRzvApjC+DuAA6JtIFXo8nNEzuZ9T7l1oPQSGFFv
egVqBNYoweV4//+9PknQGGWwekkGV+SGjekEKpye5lXzFQgpu7gtU17NFuXHAvL+1wBbFsU7H0/S
RP/7CvuA6nHA4fpdPRkcnE59jDLwN3iwMXqUMRWBbn9L59qFNPp6rv9OLh+3Sfx/oVQ5ZEBflA54
tBIKPboFvCvnlg2z230mS4a1CUnyCOYXAK7V4JJQpboSIOWJCX7cua9hVjC4XwTqhlrVVQRvyeJs
RWYW2ZFrR3cKAGuF6xG7Yjf3XcqItMCZ5nkFT22FdyzEA5VTGjR/7Zb9mdoADAnGhwh7TFCdnamo
Yvu2Igz0ZZ5fsBAHrEhgHKIVbt2aCcFY+xJOtkuHuKGUavml9JasmoTp9QedWPkx6LFPR2ySlXyA
htMfKVvwMVVlzrJS+vixTnPN8xr8M805rbY9lLl8vLBC5G9+DpnYYIWskJTGFqpLfWr5MGHTL0dI
P9DblO9p/0eOD3ebVbycu3+R+M458GSJ2sGHKPwsgk/oWb7yIjMKKTbqiOjxEd/HVqxZ/ACWXzXt
fP0H3Q2hmoteiDucVD2s6N5pMlMCbORboLtn8wBQ4NmmAuMExEvvwrFKD8g+1uUASz1tlIoXUbgT
LDctDLmIfxARaJ4rAmY6edyP8m6P26bo+EDlZT4f0EjjwpkL1MUInQJhT+o8+3Q+g7rLGCuTxTth
WWnUoz0OQWV3lclN6ImYRneU0EH7HUp6kdRXOmPXYpJwLi1H1I1cj/nUFJJ9xSsWpGlj/gv2bu+N
0fFkp7rahllOASV7sy5lklGxu+FgoGj5LxvIqcJKKMBZldj9tpfBc6vONwmvZgzPxejlyFkyjHQL
bGvJJeRJ9JSXXFkyVwnWlhe3rTo+Gt5+qqDqnUhN6ir3DfMtJljDVVFn2XKJG+3TVqZv4svCsQDd
B+03hOK7mJlhlas6E5j+MldAeMzf2aAR8HxKdWnpYVUaeEz2ilrPY56FPoIxLOwkSTz+KbeCGSqs
yw29ZimVZna3rrssCqsvAm0/Du0W4CORxDdbAM0MmsI8+Q2crnEEVAwngnT3pwogaQ8uGw6f0r5J
zT+gVKbewdRxS32mBh5dImgDeGkoIVUYB9WriznAcXiobUraUyUy0RgQ5S96st3661oahaS/rDuX
nXtaGt+z3Sl8CM842h3MJuFphec2ndmb4W7+Z1PrhAJxUl3eg+sa+uDYxg4LbxGGn9W147rmqBmu
Ym+lYJmQbSacU59BvH5trQPLY/ahkqMh+Y9kFDK7JwjREH110WmZljuGs3GHHpEjd6YJc7Ihlv1v
KFkMccxI7dqzXCC6T+RjtlD3LC8zcdPIn33tOrs1H26cnPg/FBKQUUa5mSdan9BFZYOlmXCMYvA7
lWZUmbzOMQ+Qx/er427qxbtYqtxqJ9yZXN5IZyNSkxhNQoyumLNftCI0LkuJAxNZjopbsu3euJZV
FDGWHtQztVONG7dtpin1RUcsiFxKr8iViWFEzIGcFDsxOmiqWOmWSecRW1m0t2F2aPYUUOeXfWbv
axRHNWX2wHj2KxmCoFfBnMpz4pWKv93c2nxCdC1hKwXWovVZzXSwQ1H18MTT3Y/to8pPpsOnzA6r
+HMORKsYJzY4gQvOHNnPuDVIWGvMU4f94gquc+H1rTPgal8MYFArK/tf2p3AWHbXSyiKRPzjnLak
+725T0iUrm3FqpjvkR1LHNm62h/DpvVvP82xTlU5kcCZAXMgEVHH/LGXO5IEElCW+WRQkNOQ36nt
tES2SX7hdR79oLdTBrszidMsG3hfKGuySeys+F+HWCb2JUYy1hp5jLLuA6i0KRZ0rsOZ02npGDK2
4oSdyVfpRKxtLBmzexGJgDZHd3FgjaMteCzgmBFf//IxriAEGL4+CZKWgrauPfTUbY8B1sWJHNAl
+K0oro2PXKjVOmHGTDRyoSyJwtLpwc6OOFM0gr1p0iDSa1v8nzBW744blFj4d87hLcBKZ+HJFmvA
LDa4RPIJviwPG3r3h5r9a3Nm+pIF5FJ7tg8XTK9KFSeHsyIG+q+AA8YRkW0+s3sF6r5Vf32T2w4Y
ybwXTeZLm5T5Hrcry72FTe+UghSrVX15hU82bqliAk9L5kMoTpKRo73HYVO4h0CZjlCy+2xbjk4O
+gMFXt96+y+Vc9H+d6JO70r2OYCLxsN5aYYFmeYtpKwp9e2fncNL+p7qY32T8HiemMrAp029OzOI
jWLQllzkH7ZF1ST11AtKIheR8R/PIQGha1pWd3M78RDPhzeODhKRw6658XzlDx/bqgwSLnca+uxn
TpprE3vlZbVldsR/ckj1GGJ41cMNM6VOxOJy2amLh4ypaW9u6IR0vqJ6RRDkR1loSEqRI0rYzac7
aCy7vTaeA2Kd9sFYG8d1D6yBk57nbpmxDxKoeZEwfc4gR56yQYKWOO3DKBPx1tgdYj99qcOEijkU
iPcOIgIoMpPmAdt4BYVX4DOgL2xrdhX5hRoSBV3wwP7s3Q9xcfQXGIzMAYegJldIDLnurihNZs8U
1/OHILuNH0Bcq3GxCwvuL74GmBM95vllhywzAUJRLBHhrJ3AL/1lteCM00FdQ/997CXDl6DGXYf8
q9Ya44/RCTGq3Ws+h9tMcvOSEjByuC/Q+6/HlCK5IPOmlnufxXzA1PqZByYPolRl53lu5R4ZRjxR
PcuON88+51RDsfrMpKajMgMKr4T1dUvf44+pgtFPR/8oGavK83tlqsXNGsAgEvI5tkChZd6dAwBY
lPg5j9YSHelQ37hfxYnhIZV58yKwV3N0MC3mmE9uP676Sd7IW87/6YXVrkV17pR1PHMoUTdUw29a
F51bPgMY4+EGY/imXZTPTotfpMzRFCdK4+HiA+ACl4jJN0nGoEWRyycWv8RzDyHRTSXvd5AHImsU
exQbTyvsK6oWiD23X6yaF/EJCNg1kHoX+z5C5Y643u5xt+1mvMo0vZTUqkp6hNTF0lfbgo0EtYlh
2J2Xlqgc7MEWtnVtnZ0kED1CROU+iQc12Sj/AFjiN9UFxaGezR6HTozGMHGAlcipr/RN6mzWCGOD
ibfzrKrGYBAELOCp/D7D3QKfmYa+oXeSE6Xz092gAdIKWiQc2VvbLE6T8Xn4x0ZPSP2DAUefip1j
+vMXHunw8hAJhpFQ9hMI3lBoFAYtK5azF844Lbjyg5uUM0yXZD56gl+8hVPvLsqEclU5dEmYZmON
sp2on549uQMTlFmq82KpkCnixOEWEpuvfoLSSIxf8/7Q7Ll9fSoWmd9/wu9x/R25KE3qMCEL3SwX
q8Sg4NmXXtmyWGmHpw3FsHnR+YBTx8yRAYea88rOmg8jxQjNonO6xePgBpgnVz5DltHZblNrqVec
z0+89SsU4B3ImFE5/zjpSDJv0RyJJMZzCu3PfxKfu7Rfvani5mmUjoG7WsWpTGDVoN2nRz6FJxDk
cCdG5zO4uZa5cMFmn3Cbj9dMF3WtdvVS6JmYHNgVZEMceN+k48tuEPltRXVCUPbcJshHubnni89s
L5xA4DSxvXnSWsLAlQBuW8gLa7To3NMt+Yqf9dQn92wutJ4/kvXQP813shGCdkpEwXTmsDwxfdrQ
4j9k1yNXD/joPOA90Jg4BCwX1Q/Nk8GwrLnGF6wcS3Rfa4KbLBD5E6WAk/0DTB0qGUhZxNBtWVRC
qxo4BQEw6nnEnk/D9cRsZ6IZ6bawNSo3rmVSlc2XaabxH2ZL6gyWaLKeKT1s/EWHZsUkmDadmT5/
UQlFCR4neymhyBUX1apgNNrnRptU0uxF3O9Ro89YWCLWoIg8HVLXfSTIqHaJ3lxeJeFQDO+cNy0o
JpMCMKLw+ZlE9En+acIflrtqgw0SdvuMOovOBPppVdSWNUHwO/sheO0dd4MwMOM9P42Qyk2945Gx
iiyHktdFj3UF+tXz2HeTkdAwC4KYkawcScyveiwHg8xan439u8AQeQQws4tf6J21lUMlo2rXfIO0
ebnetBkOkYbb1RW14RhM8jobKDiK74reyFixf1UXYWmxixm7qsVVh+FMsTGkUIydzB/ETMLBaD0S
TrZMe6nPkApqKMZc4jlv5zNyfikCmzSvwEcheZMjD7QLR+6f7Sbfrv6JAIwj9DQscjewKfrb0ITV
VX/i3lkiUt2zDAETRejDzMNAGpQY9TqQLTj2SjGGYCEVF34FZkqwfzo7xVoZ4uUyK9wMTds8C+ry
nV0vEDlmXP7jWbI62KYcoKBt9wDroD0AxnhEql88FZ14jTGZG1+/NDvigyFu9GsLM8/d9FEC13VF
EhYwM9Rk7b9jK8J5ukqaD6XiYziC21NT/rph2OE8tZE/jYfEEVRb+3K08m/DKq/0KUQswKQsHz7y
QRARZV7s/vs3PUecyBUclMPZRze2TfDd5gM/rwnyGVm6X8URxiz/U47+ZVICDlAX5zpotHFa1t10
DzBIdfOFNwx6IhcI4NJzghpmtYesw6xgV2NJOMn4IZPrxHEySguv9N+8JqDsIg9iHWmAgFhzqg6R
N53OdgCc975SPvk3EWC5vMVS00T281YwRAQnXmtmq9LsYAshmTg3oOlSNit1rfbfPZHXDdgYNvoB
EnXTRRDKsSXuAAQzeksNq5RUSvCJTOgEiIKPB7bucTRBR+6D5r1sjXar5yFOJfaMAzAIhCDwny57
4uLbdCFVg2x3XIgSicm01OXEcCwjbXqm//EKJ3YPDr59Ubc/ze6Bxi+pX5xcjkcfWUE9Uvkgdf15
wl4EyzZfoJdDa3w5OEpdPpjJphB1jjf5pj3+4YGRDs4Eq3YYqQNSo5l7JTAeHPMKR3Fm5gEp7aEY
gI940ORZZz6QStnsRwBdJG00ZB1QAMNqLveFptkITpS0U3AZbur3gL5SebLA9C/gCJL2mQrDpf/x
FaV4XwLF7rb0KvPaMdAH69Rk9i26hPxHWySXtx67LfN9A9zTAWHVjn9i28tl+6pryJJjKmAo5zHH
7GqYUeKULhgbQnwp7RD6ig8BjXlHwjIRh+s4w8Zvl534Eaa8rBk4f9hs/OsC48XCTijo7G7qewke
VTePcXgUho6/PJzE9byMgAA5iam4wjeFkQ0M5OuPXSv/IHQznzKwvFIh50N3rXjvuyagPlRD2aoo
pwsrsVr0VUadzBdHSlq2H1qjOJGtSwt2cZB9LcUDk8gpz/cY9dqApCkX6Te/Mu3JOsf/NM11znEN
2+d0/oPb5Mon5DlRwb5/N5G/9FkG3GTl1hKUonDvpsVrcWozftXy8GS5hIv4QsOYFER5ZV06Ingq
bv6nyHe3s5dV1x21w4qQAr2bGaP+CG0oACabJrk1Gm259Whc2CtmRtnEL0PTK0drD4q7eS/xaqtc
QpKzUG6BhW52E54u1NAfpnqMi0vghTYwuyv5uWYKP6/CXoOoGQcoRr/mdvJqRREPPU8dbbsNovB6
qUpHc2mmDMAP6RQbMHQ9DbUNVcI3adPSeJcFh/m2qCDc/OxsV03X/XVD0syEGDjkqEOdsyKOdWEG
Xq1EGwpvIEH0wj2oXWpN8XnZG0JzW7Dy8b/2VBmtnNKMDTMMRxXLSsNgfH12KkXcawQZ/C5nUFsy
CWO/XS1RGql/1dmrnhTcHsaxgfgmy7t984+qFUAvRGCVnCA5TEfB0+hY1qhUwtCybok6N4jrhL4u
R+EKchDd0jJMIpn/OEwVuT+V8XiIgp9SEb+a0tsPbn1kghVy6Bc+eMT1QkzjlRefdIZIg8ZTX4W/
c6EtPYtG3t7j2vUioSMTyDI3/bsEtR/vI3Mm8ww83qUvNV+U2snxIIIiVMjA/qp43kE17mFKMi57
hmhTR7lBxIlzPn5WfmOxr7mizfo5JgLbQ1HS0qt7uqyG77DdNYyECFmMetM2RnNGrZV3jpWVfEa6
N7ggrrucxWAnQCkaJgEyRlMWwpYZ3VxbJzC7oqpyIQPBYUPxb3L3Kuy05dyCC1ftMTTB0xxNARRX
3StQsAwmVwqVQx8XnJClH4p8l1pv0ANy3KRN1sN87JnpPb64rSqIzp52NuQDaIA3NbQ+0RptTpyC
75lx/RZCVDljIvQ+fc8Y9tL5i8rZgX3sJ6GXTEIdv3vQZQtyDtxdkhJe57NfnTNWsWLcs/U0KiaV
nmgEuHcnLYgeNPj9vJxrGgBxiBOmIbAuleGg2T5xFdEpHzBH/cDK5YMqIh4nKIIH50IzXftiaDdJ
jMeQW3x9QPkqA7Qaa3GO0Ct7AlwTuowaJkmJNJOlcgp1F9JeB6TmCtlr23l1c0FdWzwDH3En6rQO
DxcEqiI4XTUUuQXFkT7cPRXdoyN1LfdvBRB/Rh51kPtmCn+YabwYS7PHnElFpvlCXR7rMmv6X5PK
cU6yKZWg13ecbAiHurAJWk2DThLbnfRoOm+J6zcHzC4JDFZ6KvXX40DZ75NQFlmgguZ7NnA1YoKv
sApm5Z90Xtkwk5ISYqgCWdILlDZNYpyvPkQ0igY3Y4/Y+5cJT9xAn3cJoRgcteJYRMWOZhLu7JB/
PJXsZb7BBOkBT3UpGcZOGiBB1QkGLAM0QUFCUuOFUe9QcdvtSg5UQEefLQV7ZPvAT7RLuwrvUlr0
zKH0e5+WSI0uWLjJ61QoxhYJE21s5QTzVxgGBe0/y/PfK8qZqv+szdD4qGzh8E5D6QA92L+jKn/Z
99DgEFXBo5mtYGvKzvFqQHF2im9UAiDyxeJp4aGLAJ/ILU+zxYn/zwsroU69BGp1AK62kJfek0f6
cKWvZfA/gZ56M3XxZWp08lx0gUsAqDQQ/3SV/RGDWAVsvF10buWE1L5bMIPGiOcAu9sie6gzPWMh
Xp0zPUdt4pKxoRO1fygpGHHz2G7Jg9nvjuBydmE8+wgd+ARJXkXyzI58TJDaOxwQH59fvlDBc9A3
t5lQKVPaFcdLEnRiOQye0VtqgYIFD2F8Jarlb3WvRqTbbiuANwZZMi42lezIGaJk4xPMleo9m4SQ
k6krW8Ab+yzxHcyqeyo7Kp5Ce+qhJKAfq1mItFl6ZflqXWt/7fyfq7SX3s3cgqYbA5Dalqde0PJy
E75AEBofo+ClDQO8fxDIBg6BBvzHmuaKQbKd1/qHRgyyR2PzGzER3QSr4kXwAMsKLbasKvdJLgjD
wyf8Zoj0DzrRiN0OuWhQzQPpeN+gkWZdHINavIOp2hcdkKPkmWYQPuwr4cU1ZzIA3xfYrOXNbVmB
Ni9ij/qAyQZ9gaOPi9GpLpGET67XmBc047AQrTk9vLzXBnR35Fch5Z+h9WaI+qCMVSCmpI9d9iF+
Y83gFBoHwbTfSCfuhLjMzCKQI41kWyeI3rJvfm+hrWegqoEpSqkSgsrm+PSz1s6b5I97JHDk1q/i
E3rqp13pyKrWBFpuxW3tLxwVAyIa1jgTPIfCKmo3pb79IFf2o5jolPfD5SXGO8L2gLiaYcatSAZ9
FT78m648fXO0AdL659I3zK/X81awys3Ey5aIj/xj8L+ZHW9aFrZCap/izk4CsfbSOsfWlibdd6uT
N8hXsCRgLGH80SePuTUky1jVUnZEOE/GDk/cUjHXNnm7tOzOPhMEhXV5FPnF4/LfvKfzWyLfa8us
bvB2V8hPg9vvv4NYCPZe8H26vh2GNOafl4SNV8BvN5bZHyK2q/qkaPnbxP8fBQY3DyrRLXgpFWf0
RuAQM+BqVnqsepPolFbBwedwz8Uy/2i/+KJWD3z3BP+7cMKPYOUfQgvJ1JBx8f4I1zHFiBLkVoIT
/zgy4j5j+0nGOlqp8R0sfWGl4sPIfPmGy5DFbHmvlkkQfyChsK2N6E7zp9Td/hpioWtD7nJrpP91
iVmWfkPC88OC8ffkiC5Uu66JHhr27tlnMX/l0A+puQxGvkrk/UC5qBmhflIv/EFpi4Q5pbrNQG3N
0xOYdoLJPrMu93PxWG5uWwF9YsnTWxC/wgnqwG2yHmxWvn52H9jRZCRwA4W9EP8DoLLqUL4Ok6iv
LpklcItwog0q4jlmk8NrP2ZebaHz6Z6WjDDbf1obFg3ZlTJTKrAppU/piL0yOHSzwgSFf79edJz9
K1tj6JHDXL9g4SZ9gvl4VqLjachV1RBFAxv5ilpVZaCIkOOvR5V/ThTWMHeq6xNgn8+mCFM7pF9V
Y6bKnwRDC/8BFOgFk0PG3sJAW15N2Uk/7/JOnaIZB2ZQVIHHrb9zt+txXludOmXsqWPXBy3qvDFD
2431X1ubTatTPE0HvklBdRkE6wxeGFfyyCCoWQtChQQiixztnQW2bd6XqXIbaxTw4dk+Bu5NKYbM
3XvxfzAJH6YW5YcxQEirtRr14iiGtl0KTkmWt3b6K196O8Z3LF8fC6wOs9Ou5Wi1WjWmHqX9LndA
J83yKCORdNbey0suSolKAHy7gsnKLIuLpwnQuPlvkR6EWgXdbdMWKaclRnqCwYGnW9KLJ9xx0PAc
zjaMesWv+JU/mAx+ksC+H5cVvVq5EGyip1ymFMIjTVVuAjjF3CqpHJU0F110PuyyQ0kch6MGPGgf
1BSihGgrDbek5IzbDJLOntRd90k75b6yTo+xl7MJz/VbpOBLbgr0sJeCHzdrMwzbnH4M8hb4d+IL
d8TUWaP3BygiK6OQsJHe56BnmMue+RfoiehW32FM5Uuent8Xd46inwsGviN5xSK6koredqZRDd+X
5zyIw76qsK6meQP3t0g01PgBQRIYbfX5aRKEGWXIDfQQGbX9c+kNqCkoX6ouf7DMQN9CVJjIfWqB
IKP/gqf0JwviDRczi4Vl7cXYsUu9VCBE55gukoqxsX/ttEISqhYgtqzd+czXhqkT6aWwsaXhQnE4
xTmhogXZjFe2hjXc4PcLm/9DxhmyaDtneYVHBny1NIZKmAvys4EziHq8ZzCXhn1namadf6HzLDBJ
wmagdO/ZbtVlDPuD1R10i1Sm5U3+jdS/mW0E7fTijfYh0kVrIgOAN3BPl3xDi5Xu2FVi3zjlVNEP
TlVHwQEuIZ7Xbz+GBdYuvd9BfH1u2oDuI8f09Oktl0814t94wJuv3W7iTf/DTeIUiuXuVyKZ0fMV
Jy4rRbJE+PSIjw5fONMjCTKHWGa0yI1Cu8cTcBK26HprcwH3HpHmGttuZ+34P5IibgDT1Q5uCS1J
8Bq+vNmBbtalRU6kUHhWDsLMSWKBmKi+pL3+m6llZvlA0aQ9rzqORMAZ5zQMzWJdUtv2yqNtVDRd
RB55LL4FJhZXcfaju6LmiGcxy4TAdeysxcypxLY5RnnxKbnTDbDDmOeZBwN9skf/q5GJL7xY5cUO
rt9RpJEtAYJPIDhf9QviqlOEJzIaDvSvB/IE4+NGb78LrjZNQnpRHwmF1aGBbpPQR7HnyHyebHoU
loPJBHWwhzWnpAohJiQwwY3U3oCtky/PWfX58/mDiqAfNWQ/TEWEzamINSKhiawju13XNXW+Xwx+
32QK72D4vq/x+jIsCuAhx8lkugTr3sJ9wGHbhH/8Q0+qaYU+zFcTM6P+RMAac2jxxK5Y5MX+PMLc
zic5u/IZzCIfKI1FoRS+pLFhxEXU8wKXM1XXte38a/SevZLPRA074z5SzLZntXe2ZXh5o8QD/888
LoZShqvJH1LR31gluDLjQMBDo2GWW4Pve/xSoIdI0+QCxCyOAOm/3VvJC07nUnyJBQvpKrFNZgGA
zSZO6NmoGEhiXNLNX8WfE1UoO2zehiJxNGUy87pKN1kHFp61Q65wKY8rCU6RnRPHj1u2N1H5bSpu
/stA5UZw9eqydXk05fyKUh0blBhPrO3b3SWxMWEXkdZV+9Eml6FC6EB5sQaGWnsbblzr4uBGXBMo
ocYINFwEaI4V0WPsx8950XPj91OVqDo3JS6pr9AV6xCnZR3zSOAK0TsjGEkM8kmardxLA66fjvgE
p98Chyj3kKPhopeZr52rM0kaW5SM0f0aPfW6YuRu0H0lP9ehRrM40h1uh6hFC0Nkq+bO0eHDSmwD
ukEOxyZiFkZXQEgCSZsm6r440ULSzvG4Ap/6GLC3M5ctqBSlz8xXxAfCg1y1IkiakBN9MxAcO7DE
MLfY9yPsNqISk9Ycnm4JZMABFxABUFwRjuciGBmQ4zvAoub8SPWhjjZtoz4Av7V+mt7ClvWvMDd1
pCCet6b/EV9DG+VyCj6j8jiaDn+QIEH1Mxec/spk3JUG6GrvFkpTfgnojwrExDqcFPpMVzSafeKU
dsFigQ9BADYEgoa8LVCj0d2jWuiqpuMpdY4DPeLh5smkqFNAQ5OTrnRdDRZbolV7CxLaXjsLsQOp
Bnv+DF6+DWemfLOf8MyJe8GaPCnr1kSM3H5gBnn8cnnOwOeMl+1K3IO41ts6RgDxudQjtKkH/D/A
x0Y3/Zj2zO39zeDEb/j7J+QsdgsjODNwiZ4CDrnPaJ8l1K8ClYatSpHGNPK5z9WwJqmzjQmKX0uW
EfpVOhT2inzb6e46CQqhyZSdXKImtUyfOJnuSdOZH1bIrYSY/v/mIb2mSEtgFOmiPIPQRkEchnSg
pN/46wggh0c04V/V8b673pAPBDt6GLkAuhqJC00Sam5ZAnua2HyfXGHFEOf1fEAaXsn8X2as6eKk
AePE3ZycNZ9r8nijuinQ2yy8m711lY+yC3jOOmPVhc8Ah9QMRjwzkTE5Cr/g2zak7CqG2ZR01QGM
KkvHQuk6FJ7ee5nyJ7qMX7pUzfPyM5AbwP4cRUM9AKOkp8JwUUxAdi5pmRPt5N1QAaBYOKhm0Jcd
V8cmOV0oNB6sndwAX5abEt6hw0QGuC4q2MkjGP81clcwG4nGA2KcTxnMTJfAOFxeQXKj+BvYRLvB
HHGgMqa5lSB5z300p5AUkOVOuBdP/OlEcn1ahZ0OtwuAAo6XsCHgjL0zrrKGjDBNCbNppDh9kHu6
naQMOBJRD6Bx2VKZpJEaXj2bGi80xFB2WdEGRRRLoQVSQpkIfOG9qMUcYablnVQUIBTe6hgzr2wZ
8Iq2PlUh6Wr6SBia54heVifCoBDNZCr2zBknAu7Iy5S3EBj1Y9829ZWFtErQEuo7MiE1N5QzDK2m
v4nCgLUhkS6SzjzsqJSLIbtodskxyhYNywG01ctGmjxfmDJD0xCVzlCeQg8LM7mDivt12e9M8FXs
4jgyh2ZDlqtxXJ+9wWjodNEhCQ53waSCjyNU+SvuY0F7MPUHDnQVoaoC9bUr92/CRIgqy+eVQagB
IPQvscorz5/gQkS3M9MtMuBds09UU3w/Lb9bammxmXgRD1kx7c9tpjNUgrF8buMisrLpJl7r7QNC
mcEkkOMJZFJ0q79oYC22tNPavtrAoF4hXVJxDe6cKkh2VS6i0+y25siFvAwR0q4zP5X9mm6E6TJz
w0DbpSrTvI+ZcdQTQd52EW+cCgGNMSA7ERFQu+DbvdL7iZZJOsVaAfnWwvrtVwGrOV4H3DPG4Lqw
7+D0+5XIqSDMBhOpHTxmEYeCBhAA3HJ5/9gkU/WOiJKbGDHM9DgfPPu1EqyLNMiYRp0wsMjopMkw
77ZdlzKI5xYgDCa/8h9H6Hmphwgq/D9O1qVk9rkUp7HWbihdeuNpYjgW0/x+glAHVdb6Z3gY5l0V
XvnjSPrbf8Mxm0kRpjaBAyr0E/QLiD51jzAUkfeRR4xTaZxpJmNdWnDQsVTnPb8OShS4vrBkllzO
Vcs9a7T3tllb6/jleU0aD3GgtqT5GvZkig41dRxGPxBxAvfM/xSqPhUwxeMhkYNT3qj7zHhw9qII
A01mCkv239fR2xZ668dXDx5jkVyKLjfyVvFI2O9P7UpoWQEY/kzPyM3QszdysFhlNn3n/PRvWbQy
88uZ3ybS3hysED2Y45M4h6BHAYfILq4/7msQnwkfWnUtoc0mqvrSUpBnuSM/sCCm54utEMK8/uS1
cOSNUdxnbTyfbCFvMa34SUZNu0J/hwot8qa+NSU6Vu8flsJjvxZFgGh3APlzO0OiU0QllhXs8yFY
/Yb0f1f4x4TzNh8U5vUML5L/BujTalnlmZtQmLvXg1vHmRobSI/AimwqTZbFRWege7AbOxvSSztt
BZ6+EZDhRsmv7/oVamZ0Nryp6/0I/vp3vDrTEPXxXl4vgCKBEudfDaH8pcDv3gFf/UfsLzJAK3jc
2xX9o47VqsyQy+fKgDQWBzPGLa4mopmCjzAdqUzy3tb0XF/ElbfUQimxdTv6MMTkzYwEc37TaOb5
7bkN0kMX8KIPQRRwDRtkOAhqhsitJD7t2FUR2xfmQzKjafovNvuReolJSz6yJne6aOUzVxzeXn68
fih94gfvZ6dgTvjcXGQuBJBZdek253KmT7h4SLXC4KITsJxUYV0zQIqvZeFvhvzbjqXXpqQy711d
rRqNMHM5lywhnlxUZ6U6Qh8lSpBlB+kK/KIsEZpmaofdkkzND/ys9BdLftnHOhkjlFqOSgFf8s/h
TglguZoj4EssvZ4r3ZhZl3FB8x9N7fxxr66e7SaXv9mJHHZlHRexJIXbdUlm36PWwDqoN59kVWHa
2AJPLhNEdZKhM8fwQhfVigRTZDZi5KZSvn84x8aNZ4yP3cWnYbRwqdtytcNYYnKSX/O88rkdhPLI
wtcCJmK3RW1H3ClhNOLWhWAWEyMJ8HYty7cFMthDajufyKavMG1YPdWxClErHD2JoJokVA/Q02lm
j3UhQpFnqojz5t/II0S3MZ7r61YguSX0bB6AxmdtZZn24h6gts9zbLse3QwiebGQjUUSTTGtav3n
JQEIzaasK0oxzqvOINQ4xZUNImnrVuhFxgmr3MceBt59ew6ryRqfsYs+HWtIUW1jBQQMBQIO2TG6
N77J31scjsczv6lswFdKHw2qkcEZByPkRp19k4rtNmgDS43A653FK2L2Rc0VAixxehkt4f2HMWJg
MdznJFm/vFOg4rZh/gb4mRcIbiyQBpR8AQDzNNzVsHad0LnUs2M6FtYqeDZQQfQGdQWGIDVyMa2Y
pkA1k4TMQFudnf1EiEXh7SDjgaq5YU4Z6TMZ/0+Acfq75hPl2vD6dmLeiaBJa4MaR98/KPyXWPTm
rROWKl94QYgZ5Yz0XAg3JyV2cY5DGbn26u1AgsbOdas+DTe4BuJhEW8GVRHyYBMlgNutXVS3TmcU
vyH3KBCijbWZcPLBxiH1N2yfGifWoA+I7rT6snRcbwK87gqEMnQrb4SHzh+AgYliSsjg8DVy3Ft6
N7PTh2znrcAbYOVuqHu1FApQk1o4G5wqMyPR5fC9KXMqoni/nZvQ3+YH4Pa9lwuTnii4aqcFhXmE
3x/vYNaqX1laPi+4yon2xU4WpbA1Rx3moxXhfuo9Rvq5VyFbS1g5xnuY229r2Uno5PXg9/hV6taB
dUvloUviCPJ809YsMUhW91d9SPic/ZueKlFKdLp9aNBptIAg6+cK/tnFoAww77a2ndJNRDP3MLde
dhuRPbd8gTyyK3Bsz8f1DXtWbwjbYQI8Qpm3xqcO7052J1q3UZ+r7ieLBxPZeP11Z2ZvZN55I50t
mKnQTXtG6+e+ymsw0K62CApgTBIpK0Mx0Tri6lX1VjscANMFBKXPU8t6eiyeuUbza6vTyQEY+mGn
PiBV3wgRvxt2nY5y+L1RDfjb/U43dfop9Bx/3AtGpDpPvAd26ypU8n73DUeThZPwpNhJRLUMsRmN
3QEdxSwVnsUi3WNyWiiIZGMb3tTW7qqbrbeIK7cvBpPvgmkiZ4O5eaUvu6iw/XUH9AD/uiAy6lIR
emq/uI9jRIv2BVQcCzkm+TV+2YxsxM1sJK+sjSz8HhImrPO3jXi9Pu2sekvLUaPOBkaywx2UtCzP
kBtQAsC7fopuE7M7wTW/p8g1B8QflPWE7uI60p3yOsbQsGUYRizh81+NlkcG8JlRVOrsx0XSa/NU
9aoenscVAh7YD6jYVH4ipk6FakIiS9JG+4fQs+GoW8xKsqJD5h1fM7HGAKSuGjJtOa6dPreBEXcD
LQhzfcLDu5cObkoBTVDTb34N1eQFXyQk7naL77T9vl6pZClwpIqFfdueh6fjb5XHfhBQik7T4jo9
eX+kxUZF1PSOMmOwNOuJCCUPYSd2W8Xc7BwPnhto/HX9m18pL6h+cJ33sIhxULXScO7YVKob/zw4
oWOqRmaR1SxKzQEPtwSiQLrTEZtPra7Budu+X5L6ANR3lzOcSepyYshAWEb0leWyMlo0MFseePBw
X+ou5o1BY+dU6MoGAAaD7E2HHp+MPd6r7RFXykWmquMXKBzqtWKPkhDl801Khn88zUEML6j8QrzW
fuuZajSUHUVTcxUwSTU4hWIk8C+Yb30/7+CY2PjkXh57OaHzXhdDJ7ekjiUw45iBs1wPZ3bwuhX9
CiTrgXrvZU+hmBE504W1WJM9H1VMyYGly+K/1QnkMPFelT8qFZHSCECbSZuCE2nItb4i8iyB4klC
3F9zFGowTKowykD/BW7sP5hnoKH2zCvMoCc5xUlra8RBHphJNwp6vtK+OHIN8+tQZpUuxLDj3fOA
sJugIakdO85R8jmZ5RgNubpnTRss0Xe1RVX2FBQXwKL1E3G4NU5T7/vMm4zFocO+Ra+Dn0asojyo
Oi2orOgkDVHG0EM8wtoAMm6FmUnbYNWJ7gRsf6wemIvpq1b4z6q9BmtXQXj73EExScEKreJvmj2W
Hu+VJQZGLr8EtFqM24TxOaRp9ulAX1WXJuj2WdlwFrExo91EWi3WnLI/1bf4vfl7gGlEMgLpTIER
koshMFxIArMXzvyYyrvsxo39rpRQcHEbFrZivnAqHHj2qd/g2HA365jU1109ABAmurE6NYx3ZDJw
YK+KgbpzDHH2EdazkA2X2FP1ALqcUUUjxfZ4pg5ONQoa8rgQ7H65W5XjIaVAbRZr/wnI8cOoLbwN
TAsCgt4ISazBp5roHEb6jFg4koo+x9+vrEMFBZi35+kLzJEcjpZlLhVE0v6tugR7n6BrzL4ARFmR
uHTCYN8Ehr3LSCPF36bHmADrYr5TP/0wNowvkkZOZ+gf7GtNKFvJaiq+7p/EsFu51PbC9MJPZFg4
WpvE6t6l8qrSxqeIyPl/nWbXMageycqXQN+3HzlnPXkyjHip9rKBYEQ1zwvwEihoF6ONG6zNPHJC
C3YBCS+zMDlM8R9m2YUodsBZBgsO1sOfErSxV0jkUmv1Wbz2dY1FCeG4vbvCJ1iF064IuIBueKjI
iwg97d/CyXxswGuomxRsQk/9KQnC8TYFuyFuZzlIxIg2xeZ2fRnG5d6xjKKyXq+DHK1tKXSe4qTF
++CgJqWXqZmfj9LoXS60I8AK+eSt0zNvvyR4ENcJ8JZlAWZd8K80aEMNeWiRITV822Z02A5Mk+dc
iRUdU9/X7C0Yzscl+e/6Mr6GW17hGq7c9AG38LcQgcm0KSk0Hz9lCNRGflbNXH8OdTFMfYI9Pytt
fMq5KkzHfMQg0Iw1CPC9Pzqhhcukqi0LMGL/JDsI4JhPlAQA4/errR/yk0LYxV25cRUlNMilR13l
kLeJdC/v0k/ruG4xR4H3/sjdJ5GHatDLKfDUbH87swDTKHidHDghIQ4Onzh+w9XAc0+Qk8E886rQ
YE3ZRw1hrPmfq9J/zrpXtQUI3qiyJzppb2LEeWFpA9IzKJKh+ZYAKPT9C4xXK/+fsO/C6yO91zD9
p9eVHrAKeTNy4C/lX7CyThzPKfANx+B/uDziQnW7XlxE2BUqW5qbDfhMGdbcqiLKw5qIywLjBFpY
Y9WW/ruf6aaWdDS6rFRA7w2HFzeDF0Cj2WVm6sJGrTrCgvPUTpuLvcLYJHCB4MZP3uYP/xXrzVV8
3kq6HKmuiFNrtJ8iOCCttARJzuu0+Gjc10DxUEuaTqAKkHCAIATkuQNBp2Wy3vesKiH4g7y4aNeX
bfaLcU7jVD7Ai6etgg+MppxlUKNR3zkAJkJZGKxPvvxCsT50aNSRnkbl7T7G132uRh5IO7QD91k3
9L1UbfIMA89+O6umVX4w5w7t+LUwlFpArjPORmXqeiDchKcbqb2WdNkWQ5U4r2OAD3QJkjvxXkIz
bg2HtEMGiyNd/UQ5hXe3VRI5asCitJULrl6RdMdCcpWZjlh74zDOigzN2ZDQ9looE/S+jKQ+aKYZ
giCmpTn7hf9JmKgy+bhutn7jxMJdq3QZ6MuHljoiEJ3c8y37SrF94JP/xQt9b6R7F5RL51XcbuCR
p3C04jXbGknEOHrVjzTOp1m+3o5WSh76Hj05NBM1D1Rc1JocDfuhOJw9e7JtyyfNoyAUSmdh3kXk
yhgc30mQXRBdL6M49AfgBzLJjRrRpNNiaoqZQJiL4zw5sxLzVtTuohwwdt/1rmko1I5/sIhIGNdK
gXqv/+e99KtrkshBZjNTQ1kzlOqzxYyKLsGDRcw7Ty+ErNjG5aEeFtq/X+IXinvYMwILZrY7ZJiD
a101pR8SVXn+MA7gV7qh8rPkG51PWrjS90UrdSbPSl5SedKOlqqz76xjizPsTvWNFEHJ44IIv3rG
xDGvQ31GhdF6wI2Cm15iqAcznJvNF6APSqk/xEogRFMvuqanI0NqRTSZWclDS5W6v6fQeArqxGKP
djGRk1o7rzi17CwqdKxG/BT28xbQalGouPtYsQXxMAkt+Xqkif8NxGfjRxgos3l5ml/7f9AZLb4Z
ZVrp9S9JPgP1oNwaAp9xEWjJgbOKYwwZ664CWZNI6kDgqYNwpyNUKCZDQm+lUGVt2nKBVFaLGYyU
icTi0l4jKZlzkJwsnSpJSi7gkEveRZzKTgMmrGRybiuh/s0Ov81jR/O9Wz6duaHmlSvurICC7wDa
fd/zKpSwiLslPVfIHjPB0z9GQuz29RF/gx6mFnM4XddswrYShFdCS3AxowaiBUcwS52tmyqcZ4pK
eBSIplBeU9E6EqFHbCRJV0OQk2QlTkIynG14RHeYYrAFyLjoatYDIhIXKW4WLI1BuCUkDNQZmtWN
FLwq4JNpvbDQabSgILMD75h2QtSGPE/r2sQ8dzXThGNd5a//UbiXGxO7KRcCtfj4SwqKGzWB6oCE
pnZM7fuKMSnZ0ULMRT5tkMYhCNEri9CUHCAChjv6DRRi88mXqcGEFt0aJI5qz9LiUoYTWNIowutO
IXi/QrDteOhzow3hsRubVMyQc/XtANScb13beXiy1DgQNFGldtVNXSJ0OZZgyKg5HT2/S8RJ8pVh
bKVqWkIUrCW0mr6OzDXTieGBxwYhJMiHAswIvmvpBVjOjKSvDyHyyO2xrPN2gdfNnYMDY7v54yxR
nRNkXwpb7zqdBZnVs0zL19VbnDZawOT+uSLq8H8SSyrhT+QY6r1ntRRRu7VbO397lJhEW8kXKXPG
bXypAMVNgancAd3J55z87p3e9gFooPN+XqnFLufLIRcxoQSSUFdCi+L7Lz0cPrHWi/8ovBMAU11r
DsHfrI4IsNd3WlpBrWJl9ccBi0eH98MLTtGPLLCCQi49wBB/qlPAu+FUL1rXQWOwkbhJqd5zWbTS
Pbs3Ty6V4b1UZIeXhXHaJj6fNsGMUMSUIuWluju7kOGuX/qliD8bjZy1/oW+rKsptL8pyvIw6pKi
+cCLkBXggSen7nJNsdkP3IsdMn2XSrm94h2TeK8piVg+j2RPu6DYaaL8yhO6+V218A0CjuHIj7Do
qmGiuQIveZLCF/yNKfDHGVoiuRqusmkLccMvOySr54MfObr0IE7HtzT67YomUgS6LwMnKE5dS0Rt
55On0X2lRDatkt24pSrbqk/ZqZz9Y7ynGtCiq4hObWxDsvg7YdG5PlW43PY+tMHc85eaYYe43uWI
3dcNqLqTPOQaM475StdzEMnsVzaDGpjti2jC7hNVDT6/ldXI4qolZSYKH2/JZ8SV1ibjuJHu5Vkk
zut1JlJLWtrdaz2MAy1TYDaSgYYBEkIfN+gJO87JjccpJzA2HYPH7eH9xicciwvBoWYJy62f+B/x
KVwPX8Ocnuc5DlwasfQtmmxIXmF6CN9c98qPPG5NIQ9yy5sVzx6i4gm1YhYO6pYniuEJ9aD0+Q0d
V36UEcfAH35spruO6GehJcVw0J5qKq94rGMkxfXVzipoHx06Rr4qH88Z9+9WYWi9p8sqFlizYN0z
6y8ngWG8whz66HmGq7pRNLlvkiYKSKzR8aUR+4CAfX9CG7SLfcD3Mt0gsI0KgbrbsmPs5b5sB6BU
Tgw/5vBLqkZrUVND4bDrSEwDtwarO7RFYLj3icuLF2Q3BKkdpvrRm+ZRLUaWupmAjZu4olglYMsV
JxIJH2mRrwf/e2UA8/e56n1VpyxNvfeqf3ORoyl6PpQTtoEjomZUY0H1YF9EsMdHh6GxSF2Awvt/
48WZN7fBx9iCzzP4qTI/pGYycmaf7bfcAlHy2TENkunjxAxYRr/UKlNisWnInjlz3M1Du/hFavNz
6qzKsWepjd/t/buclk1Zej17cpxtGpwq8AZRh6ZlIVbY2AH3rrXxS+9CELFSHjOmzBhUMorn9v0Y
FX726hIoVZ2RpDSJ4aXAuyawFyKxyoQKZmL0aMdhBJRNYUWKiJewSigl/qLgDnKoV2NMtj1HvdX+
HaFFraw0aZrrpGnWmTaS6z3bCW+QRu4b4t2E78HjNrUK+DLBIoA5QoqN/rRAnIRXisIAUThv/Inn
GCLSOHPKMBARyp15sTQWjd+Dm47WxNXxd6SzSqPV1IFwW/NPmLvWNmZQY1yYUa/qprV/+CvLYtSV
tPS05GIfBIVllH1VobfTUOVrfkhKLqzxd5teaxBtr131Apw6HqbwP2D2PWEOB6GKxpP/p9c5Odi1
CZ8JqBKY17CfG2Sri+VQ4uT9nclVCLnRG3ozhuXIkKNTaHP29LH4viU7bkj8n96CUYyWtNsJdSno
CXnWJ4oqXkUsov76kTQot1NmbZmsOT5cvXLFKuKSznNq8WMyDtoP5jGtn9mzvb3RLU+K9w93QCXS
/XOdoiVtGptQrwRouzCnCf3pt0+rVpWDscVwWr5vROXMZ6c3iRumMNIcU276XfCo8yuvvH4VRVi7
lxjExqduBAGZKKKHXRxs4ZWIszluETPoFU1f0sdLMQdpFkj4iXnuBiyvsG2yDOIE1+iOXWIwlJBw
ZB7xkyCHRpwtWvBINi/BUV7lxYMXpna8eJXMsG6+MCp3OPrDLqhAdfPQHr/IVlPWaUipI91nO9FL
spjY6bbGc5V0EJ+zlZjqz0C479kiGBUh9sFLd5+6HqYE5UuFMbqXBJCgqkjeBHoRFqUExTO6tA8p
bZ1pKBtj/A2Dd6eEE8xenj3VGWw2H7p/Ux1KY+MYbH5AH5cfgwGwFG0edWxRw3qV4/fmRDy1C2j6
a/q6kGxHe7ABhKg7rFTbuTAQQx9lpukSpa8uiGzNQRHWAT+VJkueNw4JmblFVBYx05yYtSJSDZLw
rI+sjS4Py+JqNcAac7w/Kz6eabbWIcVJPICkoSgs6j2nRdbai2b8GDzz2sF9vudBBODmo2G7vlAv
R9hO7jzaWSvbEV6sYmVhieUfjdSZradKSTdV91gPwu/S10xcxJPq2SMjw5ZVcqoCYgih8pG+R6um
e54OheHmkOhX4qMoQtBVP42bUN0eBdHtlzIuZgTu28McFUt1PRru2WaO9m8RkjPQVd+Iy1bcjkko
ImXTFy+7neTi4Kh7uFZ8UNZceFes/dJkvA4VNpEfK5MCVbrligSQkTx+WnztsJvvkIo9r+sFmGxO
OlDY7kJo2DIVW/DFA/4ipHujKRT88s1vIm8ZAW2ElefQlrFAnlihN/OEifzubLXZ1PGCCLMNkInl
fu9u2rfU9ZhHBVnAHsZmJ4zWdTJ5gCRLaONBYixTii9+y40AeKZ2hD+nPy9yEu3KauzRRaf3G/IG
e2ztZypE0KfHDXW257caXHjmBZSf0KfhDCnwCIXYOVfp1xJ9epYl0FYTHgYBqRLhMEIoZGpLLCC8
7YMZrvTeDmpRBMwXwPWj2IKWO/+7G5g6pZCDvlqS9xnHpTgrQf+49d/CX6TJsCD6Pr2bEPsmbi15
xxK2cAIg/dPucxsmsy0gldaeL3uIB2c2pUj8wLTt+TQieqnCay+T8oTw79sngDIpfneWFyU53RCw
+ZsoVenxsnZyZRLqRi7Beyp3ArUjY22sF0Q5jYrBvJmDOa1w60+QVHBq8lh6nULH7PRPbN5+FP06
CIsanXHr9bri5WWb5qzJNC0u8qFiMUbx7hlYn1DYoUN28XjWGj8gA5lrBM7KqRXGZgrmBLDiYtq4
Tyzor03OYJC9vnMS8QZHgV1k+oyYYjxqWaunkJknb9zG/GrxIowSuuY6qlRcVkWzgrXHAwWbCWDJ
ubgLBI79UiP68+mL8Oa0CpWjb7XJxYdbg/M0CLuewPRfF1a63imgHir7sFzIj2TXPrVfvhe3uHZg
jaWJ7zBNIyV1oaRMli/QEoGdFbUdn80y56AcWntIvbAdgb1YvRL6qp8LOS7VGcLXYLBC/YGSvKDO
iYCmdI53aguTZjZ6/UuwlAkUjIjTGzjWQ/FV72SqQUdWvfGsed4OWmaaWwN8Z1axbjKgsN+oVQJY
yGUMNF4oMY+51DMasYJAIZTz82ygVOgGJEiuQC8pvvp8fUScs/eQc1t4AvHFWTvMVJsWK+m5VScx
IuRZ/hNfByiDKj/q0EoihpOBCqeoKVe3fTcZhk3rGL9PYtneavbebon3KBvKf3owtiFFb2/okywl
LH4icxVZv2JWS5qyyRRhZUjYu8Rm0gKyp8ZWN+th058GojKH3yvhfkr4hCAyMnSbPQ2zHb89Orpg
fMidbB2lkkBvZ8yBOBLZ66XTpNRG51lAEGnF8kkRjjXU5sXIq6vPLXn3C4TmFUSJZCLX/y/URD+x
mLNU8ASZc3omvS2R/ynZiFAzU+Zl9wE4miOmZIemjyveDnz7CfHntWiAaB8iJX+v51GkNyMf+mZk
SaFR00spJDyjDR8d90Xk4FWcGzCmBmebeXaY+Zj43zPWDAYIeslq21NLKPe0voLqK17c+k8+HpNK
ikOfc8mRDmSOp6ZpI3IzIlUGGZQWq736XmRFrJ2voeOu4ko+kxwwID7rqcoNpBba0qSi1kQYTgkA
J18BOJKecnbn9xeYhIm4C/jsViQQP9OIpMh7wz2+h0DHvZRxfJiWTF58KJgNotcT2FcoWBLEilW0
lw5wU1wNe0+aSoO2XBGUo73e8sosMcdRSDHWuYVGl1A1gqf2eUTmwC8FKtRlJ7OcIJwlHn7qgrjH
0FO919rQ+15skgA7q6PXvYxpZLPe6y+b5bAiRato6z4w0O70836qbiqSaIAP7lwawzoFIX1JmXJf
WhsChJN37CyC/ArdX5/7QZeE2GBUjHUJJ5sBckJ3ZVa+GhyepN8C42wU/KFOOdGzYdsnljn+5sBM
mGIGRJiGFp8dcAwJ5xVA4Fco7VQpanT/bSulGbakSfhv6z8420wll9bp5QhiYLHHhA9A/Qq0G1rX
MFe2g+51WFqkS2Rf9QTZn/b53W3cqxizL/8QhASZb3VVbKz6f6NSPsmLjUQedTevaMv+Aov5rLjf
ww/eW78ZSFN/m7w7W/hwYYitlMyeNHVPEIYLFhbo/1edwaTckU/bvjBKKl6XX2dniRsGKsCE40Jp
7BI5Z2dMmpvrThBVs1r2I5oB9cMBACNfCMJwgXG/LXG71GABmKCGRmVyHKIXqFCt2IDULEQ15ZAx
ryARTBPM9yISfc64TzN5e0k0DfyeHxJgSHdzCc2qVf0lZyNRmycmCi4l7PckxX+BMOrFyvqzE9FL
ml88ApMot0oOin4Q3aF5e9BZqGuAGG6B6o3eH8X4G1zgBx+tqusMM5b6hsfD4jRbXs1wba6mH3sD
jIPe8PLcD9ScBvAR5iXnZSMXgQG44yZBgMclvT/1SKYUlMxEoKKaCvf8bpvrjArdPVHcbP7+y9B+
I4yBALreHq5R13R6jeNjvniGgXzQrCP1FP/6C9M7zug1ZqYNcfpd5Gl+qY07vp8ln1hWmPIw9ar+
cb0JY/G3nqow0XDzwLHyDJ1OGA+IqgsD1xJxRPGY4Sv7zTZYMJzxMomvl33hAuVF7L7AfMxnUeIw
bvsZFZc629Kbtk6gzKmFCHTL0FhbV9q/+4qh1qM5a1mT9rJpYb0va2s+M8eBxLYS03xZBUOo+MiS
xZnKjrLYYgcldTyJWs+7ttrceB21lezeuClK9MtiKRkfIrTrDOl8SmKpj5hVZiT8m1FiNygZ7LHJ
qix/ufNEosEgVxNQMwPm2JwbSbgK8hLcl6G7ngf5D0rLCeqJkmY9IUtjmYyeoAp4XAvM2LQXzm58
8+F6AZ4m2gXgAE/wJwWl+iEVODI6POmn/03LSNkNlEGesqiPrtvWf7EQvNb4Yqvm7fLWSEoBOaLY
ilk4foU6oGXlRVqV0ymD92nHSwczrqMGxgKN3laW5P68VSRCRy8dwh8AJB28muOlPVvA2cG9CYFq
b2IhEOx2/BnQAIchtl2yRW3zTC5ce8KRumHiyoHRVJFlhEzahLHsZULr9SHzC7GwZQ6Bn832iMEv
UV09s8M9jHg3P8ONvtmpzeWPdO/eXSOs4V8lvff5NVRphVOCYXWdPT53K1hKiqJSWeO3aHPM3pUf
VxTzP1hEydVkJWiHMJGoslpvv2xBIrGOOZB0IVthu0DSkEWpPosoioAbAQTYubpa/Woc2FEBr8w9
x1tlbwTbsnT0L90Vm3TaDOP8XSkyh33NfCTnVVvs86emgOwCaPmCZ+eD+jrzM49R5DKnPBzYX1r5
EuUdv0tuVe+Q3+dO/gWAPEZ2hLMIEHnLmML+r88BnBt8Q1Jewn3dPWg1JNbcXyU2h6iO6H9cUWCs
AtFzg1USPKhBhKf4Wey5uukJiJgZrpzOnSwdtTHEv5HzhRw3XE2pDf+XkUW17SkoQ8oLobqSdWEo
8cKkTv6FV+E74tpAjpEslOJFlnP1eH+hY31/f9Dnv/MTy2Xjk8Qc/XMKRZ0pohETCxWXJ93kpZOu
STvPANaIYt5CU1R6jNLGHdHUkDM2tHmnrupYfK4Y964T++U4D9oIHmZVMiz6xDPgP7FBAIkgU3wL
IE7hOuIn6wYcxf9OtGZ7ALZJrQr43mgqGJ0Wdddk24Mi0x9ooQOQFI94alvHKo7DwPYUIg2p+gnr
/iGYkkRm31hR/GpdGuCEbx6HqpLWuuk/DULXpYcmoxbn3PPKWbySPsDi1swoXUJwq9ohEa0oWTeb
fOR29LSWwvlsZKWqMvc2z5bsUlwwsS84AgtAo5XpN7/kqMIQS6yTrzGadztD6Oxg/+zvNJadlrJO
8quKSjAqT7eifsSVr5qaGZZQa8F7tN05+/Z65EFcVkG9lpMOb5YyQnhC66oSg9Y/DIosf8Oy0cJy
6k/m/XiJHDxtusZMO5mzIxBVf/66oXQysLXi+g4ltShAi++zN5gkHSfXn0819mQhrMJA/1d0vYCN
Q6zmztfTbSCjjKn226yCgd/Q2kc1oONQpeIq2o15npg/7UuCG/mvctH7gSFHQWsuJ0XfWxgAiHNv
31aIF4bCgbhJcR13c3kmoQW9qf86E377EyYaS/eyjlbKp0gm43yvp/M0dmQ32xW33aTcdIvUiz7f
GzrP3QScR+hvNMrD5lYTGLJCeMMW1wVdt1Z+KrGzjnU1VFYAC6Wij7Td6jfBojEu6i3pF2j6CxwI
CstO5jZ2KvbEXrib/hT/VM+QuT4aMg909N0KXGuY8NwQSwiuerEGL7FZQNnNRX7RT+GZCg6p0+Vf
7Iqrf/073Vc6nJSCGOp0W23ggqf2z3nVwmCgLT8V8C6yquVDhAEtgHbYjRxsTimxZ+EQpFcr5M1o
MI8TeqVOAI1r+kwvcQk6dBslCEG6negFxCkJtWwZ6vra8nxDvb5XE2nysQ8PfffUfKnty/r0jafM
Za6rF5qsKo5miL1VBMS6uHJ2MQa5T9pKdJ9tICTFOuoFihCbqR6PXtKWORteuG8CyoL6h8rlpz1y
slDaneYPyEsXm3ag99o3k/s30dZ+1EORVDAtCBS3aSm0RyzBC2ZwyVnHKpcNfxLv+6c78Auea5hB
PmbtMBZb9wsP5PFUOP7dpGqbVUpDJaZsVWrUro1FaZMOQ9jiuRN0nMU+/YP+zlTCIzQA5FvrHpxB
CBaebllYNoEjeAYInXEGimr8qgfHRj4NP3t4dzqT3jO+e8ZTEj4CkNFpRqVvTS3YVkcyH0NF9qtB
efvEnVEKUHWPEDNhqdCr4LLOcDnq9A2aFE2Wy4YzPWSqN/rll/6cVIfNzw8S6x8t6S7uzBmenOcF
hUgn6kr1B4SrTKwMac6U4OE3NEGyj+wZPeLilpXY+BzjixNbk9tiVlaw/ZJnHSWFT4tkOlKQJomc
53s80tjetSdoBX1WrbHvxqrBkiBFDUjVua1Vsq2N4YzRW3P59eroUgiQTHjmMvvFTGOFGEuJZDDN
H6AO7TU9d0LeKNhWhKDxzO8B3c1mvhORXf6qeddi0QzSL08xVu+IL77Tj/FRsNXhgW51yDocP6NA
JprCUgMPDJZHSQuNhMK3g7pbH5KpMTX9HfajOOUCAacpyuUg8HZHErbw0L+mZillbjaQuxUUm5OX
XKsSHs+XqbNkLutUjN93SW4/fy3L285AulBobKlNnuan83RYEan/vijfDuDRY5bAstOA4K0D0UVr
ji5WTcKss4a/ci2oUO27n+HOzoAsIfKMLBeP6bSm/1kBIrEjqWHFF9sJ0InXGXAv1vQ+dIn3k7+E
yXKbyEo8Mlodahua3QEIbiQ+d9OWPnvLCq3NUk8z9wCxwgatFh0dXhLpIKpsf+E15csNRFzJlN2p
UKgZYB/MfiQrLpJ7pfpzhf+0peMapWrks9Hg6qswN9arNiBpL+2eAnvvbHbPthEFg7YQ3nqxSCKG
P4sz9OoauMtKQ95ffe7IlPZ2/QaUcoEL5c+Of/u1bAlBNE07UaqGfMsoRqt0XMLoY8ly38/3oeut
8OdsTMhjrr0OWB806ytvrTuSHCOdNb9rx/e66wZK6ODrrFjE6y7gtgvCTHyPTZfPcFytaRGJXDxz
7akfCJ2wFFglMrxCylRqgVfHwQO8hQgJnYwnbXbvvNM56fq4GdofQb6jyjGLSLQn+fcrfdqsKKut
PmAeZFiNaZ95u+Du29Oz8+TJ8w5FisR2ND9/SXgIskjpajT8jDlltIa4HpJs99PvDQ4AHEcutDKN
xcuBjFTu8mPMTqDrfQR6Rb/T4/uydGimpu4laMgSmhGuzw6alEBrXOx7nDfG5pZcr7K7GCoueYkU
TqgPJiTkeS+VjSMTf0t/9oWr9llJDRULySym4tipBRqA0Oy5nGVmO3h7+SS3UZ5qSnekbA3G9dq+
cEDFJ6e0b6nn0X81TBJKwpVHs3vgrcAzVYupf9kJF8+H9X/TPnftjqeRvmM9yvYXNzKzWgcLwIcv
E8b7b7lanGgrTJTll94xxrLyS50s7+tGUbXM2VKs0bRWduqrVEAkDNaR9jkf9Y15nZRso4RGdNEW
Oq/t0J9ds6e0eKUuYI46/SaLWw/0RzafnEhCvTH1o9VNrqmevlDnzjlaTT7XePLWlDrB6xv7L+gY
/cGmHgiFeMvx4xEqWfv5g1QMvG3o5i/fzWphER+377F0bd5TcbD8oA3debH8dDg5D8EZtiDdribo
MqIM+w1a8SM55QQkUoZvVHksf3BR7AQoW/rJgHLcN6kPy5fQb4Rz1v+WMm9mhi2guqTPv+8IBY9P
2T2zBk3QisH+PM/YavxoEjlIIykV7C8qJf3ETOjUMj4ymp2DtbmVT25r31LXFuH6BMTTFeUdZjzk
mtjQjUJxHYIv+GqPJpLcYxE02IHzVlv0CvuBBPNFVrboMg8tIyPCCAw9Ug7v30oVm7QmczTbQHPZ
NnXZ4JIQeJZwPGGeiJbWYnAEI23nlTlRINgNOohPrFC1xatuywyKX729DthKy1avs84g6rIsbtY0
8PFsCxjXil/4f9kKz0TOX21tPH33KD9cyzyIu/kRfwgdzNESzQuU3iBIfoXRk3oK6zPGxE6+Yexe
Kz8o7lNXZ11taXKA0gBIQQkP4o6NbsyGGZgbtKKEXzQjoSqmQHbtlKTyp1Hgt1DyX0kBvdh26ZV1
qbQ7+v5GzUxgwet5DqZnXQ1LfPpSphM9PuejYPS+nWR5yoR/56wZj+szMxBOzm9K872a8HXE1Ohv
qbmOAYGeivizeTnvomVJJ3V8uEMDtHAMtaCCSTPIGcltnxWERW8CVLdGaam+FyPi10FPdEZj1tSC
yjKrbWxOeYufehbvK3iH9VcujUD/n629HwQjsxBx5+Z8bcqkjaahOUlFfUmIwT8jmpHtNqdnHqyR
eRWwcwai9d/ghwAezt4Dyf5m+i/4KX6x2HlqySQsMPP7rbKLgJaYX3J3ym3vfKwtyXehOGKL94Bk
7y6k/iRTUFBKtR63ZbmEez99ikMoclPuJk1CH7mhhjTzRuOJUjwwKBIVc/9dhkD2MaahFohPEUC1
Pq2N86RDMKtx6pXpl723PY3vUe7i8jzmIY7pEU5MlI7IZlbXASqBCinpriJFIjkXUST3bt0dSEg4
J0829ApxM2ucFMMM9PKQ9/bPnU2+jD0BiaMDOqXZx8qff5MY9lPOqMuaaQhPQuanKPDRNmsIF3Jj
xSNxruYcEj6lVnsnMp4oowaUAOyNtZcbJ0Cexgyimuluw8o5mmLFkccyFZoW1hOSDhRs8xV1AkMa
qc9/UWGuSKYnTO7QV3gvI5X7oqQ/PxiCTLp0oU22R9qlOHnOXJun1zp8ozm14bcjUKdxU8wPXiX6
EXZpftrL9463spHJ3lpd2flO+wZBYq7m8IBRWrpVbm1Jexey+q+KsdLpPDz/xeOEBeZK1s1mhOZt
g9MWti5GBvepy+oRconJh0xYPHk5Wrb0S9K/eOSc6PUPISXGyUuzXnNkGlWqGtF0mzChnDIpjxw2
JBdhn9l1EBFSA6nBgaDHJetiGw2k9V+d8B826fY1970wMT0Hv10T9iP81RT2opDKFPygTxDbV49W
UEANYAPZiIvz7m8hu9oKnroefTc2ld2W4KdccLO7i4vJs5BmJLswOr3BrsHpMVginlOwcoKSd6hZ
OFLpYPzzi9tPnY+9UZgXq14fGJf8NmtPsGzYMnENk0Fsa3aV1tntSTC/oANf5lq9BMespns8lzBA
3EX+zjhKt22JB/UBrghBugjJKTaePuvj/ngtq+jobkB0GHzmxBsjR5ytx8cdBl5bH82DCDn8WwYf
BDU3jyB+iJRiGhMq57t+SkNLB9VRTUPRw3vprlbH1WwWe5v12RuthknZsi1k7ykFw8qxyv6QPRc6
yriGyU73aC104TpJLwImhhnDNhnHF2Vz+4VYDJiX8f9y+HuoorJ2QySh4Qn1ueu/QZ7NgXNbKhvM
ef8MReffVf0R6Yk3vW5/srVbQ6vq23mQEoChpXrXn9E0hG7nIW0bKk02/o42LgBHclBmuqg8mwPd
IakU43G4M4yJW/RCVWRaLqejIqm9cR874x1PHdT2I9lMBeL3VCXTPSWctCuVpMbZpEsoPTcDd2it
xGAOgFGtnUV3Cie0KTe+MHeFsS+RWC1beJ5rQ4qJJ7iPZNAUZfHivd1znUhjo1EIvzja4gHg5cUJ
4yr6QR+6zh2S7CnCgdR5yE/YcdMYGJR46uJTYr3DDn27U7pze2qMCa+j4wCo7+fkN6JQSvQ8npND
njiTkPbdmPL48ISUYUec7VD/XLm0D3L9CIc/CSicZXiweLGjeSDDRCex7Oo9ArleLjfJq96lHN6R
6ODumu898X2nKaKZi67GtUz0xZwbHj7p4ec+fiJIBNyrT1q7aFVV/dg0FAjM6ZOFUqJQeNklNbJn
ZYJs/9Kz4CheHcUc5vRqVyOTWgE6r3QXxvH9pKt5kpNPutnp5HlEr1Y3WAtyDsHYcPqOg1s0l2tY
joulRNtT9BIcmHzMQdSJvbcBfuhAaH3cyN8ckGBE2Fz6rFWN+/dejmbgk3+shOWg94xJjiUpRUcS
/BbLH2wfpz7jBjCRl7okYt8rY2X1bt5hvWrp5zl9AtEIarV+SXGRlzCzK4VuA/xgR35O14gx9uAz
M15jvMkCqW34pd16fdnaCFYDGfEycJNhbEc8CXcoiGmbG2uB9eNJfTqcgmYTq6m2KZhbKZpwPKjf
ScFmY332R9exezFTuZQNs7ANQ4veaMULtJKltH4QSlnJ4bY77jHOyrRkivXJ7b1OOZcKuJLUcIcI
TEc0lnFBGJlAtNpcsrAK3WHbdrYmMcD7l280o7UanbJwxEIW8zZ4585z0cR3JQvw0QWK2WC7kjhi
JuL3ZSw2Hp1oCRVH58Xbu7psvrdUMXyLGk4ouhn24aMflhuMv+mFRxIS5OGlulx9hEwZzqBU0zxV
KbDlSng1pGYIuYZClS1la6iwH/5kaoLc4n6FfShPAFEgDGxaAFVRwt7un5xCwyuFjK+JgiDGyG2w
f/rpRtzbm+Isxs5V965Kr6FOY0ii5cgOWOBbiTUm1Ucg8RmKBurYko3m7Q3YOIFvN94b+If5N6T/
GTfdTlnGZJTXfdDm1Yf5oiUkJCgGy3x/+Ag5dEI1L4vOBnAk0AI9Cf+UjUfIVJXeJepSkT41bpkR
dmqlgnRzJ6OwYTzEDL96lwtxpuLb7voKY36Ik7HfunDspGkrWYdlNT5QiHwrB8RcD4OrBf/YSxtR
TIU4WLXwXlJhUiXAhc51Mdalf6aOMd4mSbKqNvMC5n+qZhKhzCBQPnVsWyADAuHg6bb2SHOulrhb
i7bdEwS8S30/S+vOTmsNweLNyLclzVA497/feVG/KmbCp4ggb/F6KOcRpusIN7XMiNyFyWd4jDY7
DsTaYSuV8i6K4Zt3ZeqBsHFWrlZC39SHp+lnb+3XBvZXHbdooplFLuwitaWpc8qOCPzFrm/iKfya
BrZZXMd/3OKPwdHNNtppogxVA2aOK7MLvfpxHdiAq44MFXsNeFI9EK/2tlJjfSURw71zIoqkOXFV
dMWihUQbKk1jizX0TOsTwyGygZH1ub3AJxbMLfheXFe3V5ZwYScIRxvuCTXcpUgytuPjWM10K101
L4QurQmEC1V7kJvQYxhPaFKBx5AWFoLiOilY26N2jWH4IVWNDFh2veY3bpLQvQk93nCytlOrEPm7
Bmr3fmyT4U4H+58yAgk/vq5LLMYilBONqKIeDxaXtsc55D3qFFLLUtCjCV1ihNTjKss3dNUSHMAs
od+ml8z1to0vXOsCg/oaNVgYVanMWcnMpt6YCjgKDCGsslJ7hvRXriaDqbnfKW8Crl1IpRq4ADtd
cXG5+oB/QovTrmKv7FNN0tuJU4G0638it+AzoS9SWnYSzahbt+TTh2mnGZRANFw2WJ388W4xHC2f
jb8Hg6hR5LjS4F/fD2yNyAFIYnyDYSx8ArGo6O2FHl9zI6Zz+j8Gip9mIhu0vmFThkq98Gkb7LTw
jXOFNYIX/8HonFj0uEeRvWYv7DxHWKRMAw5r91wcq9oJkA/10d8TtdDUQXiREZIzteebOuBWCd+U
RgQ4PeSI4amS9LILMIj/4MByHib3RwGc1EQbWG10Ha/a9wwa67wXerDrisiJC/s0b5ltcR/EvOs5
VNTJvrpgEKzJ1tGn+eShtu3GiDlZZHCUdw+1BmxMcuLZfqYr003GEu94fNJr3Q70N26zyAXkeCqI
Rty9YUXYbv4cQemrXEON+7yPmkpONr3sT82hd1dYxOYkkX4CkAV7C6ZuirmxufuDlJLszLrUfdVa
T2GCexkx/r/SoXGm+UT8FP+XC8F5FdV4FN+cLijAK6+aBF181bojB0KpyWWPdOGnKlFAf53SYGmC
jIh9Q9A5Y9nZlXecaotnRoYd2i+l8nxHv5o9Xln7359WQz09psryhgecqacTO+76h7AyFYTg4vKx
NUzJ53eLJxz9uUfugdRBFEovb1e4WlpEmXvOz4BQiO3P0dEKeDUaVHGRnbsTYOCtd5h2BPYIp44Y
vXTpo1GnpPjoS5J/jkPFmswgqfdGBxuPvOTOA41c+00uRfnacLS34ZMs1U1DKFcE7aGZ836bf3Fc
xjHFHrJh2H4KB1Y/tlQAgzAMfBrQ128JTvX2wjnRR1DzGiTqlaIKC1+mRhaDhACKW8OW8cY+a1pV
zJ0+l6lxcfudm9vkgAFnj6N2p5ZVndsHyd2IDBgeOJKQyYY0k0z7euAc5QbyMPDrYWahiP+pdwA5
rfS4CGfrYOHCHRXVeBn3OwczlHnjqATusWBRvD6nQG7MZNqvj7ciT69OAVZGo168umc07HDR/fbn
ZfEE7uIWecXQf7d7qEENX+tnPyhkU1tyEzjchAor7vTyLBp4YCzQiILompqDmcvi85mclVATDBUd
50gNwd75hpbwO4b4Ukv1mpLItETfF9MEav6ZKjyPPiN/q+cDZBUTWDkjc1ImOWTRi9ThVLZyzd2a
3poB9wAB1pmPuboAn6Q70miiah4jd99UcKI+qGMaVLwdz89M41UktyhfVjIWU9LeY6HDafo+QxC/
6SKmCrodroSii8nEwOJv9L/QDjmz9R8n3mTkSHC829KwEgc5ouxBbm2eVrHx1+sLH4DfVFR2AHkh
A2xNomX6EGUtmsQ8npjdtNxiasFzBFpqcc2s2ddBe/cyoDVSGA4pdd8WocyEotByKYwPcXplGHBS
nYccRBqc1BMulR7ebYHXTLc3G9fyAp/womS+BBQ8/Bmwngp/h0QSb4s3eDnRHimO9Dvziz3ceTGE
frV0dzPr/9D2DH7Iy08Z+AEPrcL5XFMJBvWPR+9Hv9rssnZxs3ZYraoLIs9N0v4ke8mZTtB7ADqO
vLaemjUS+ApPRIfVl1YpqJa6X/td+gA3mwXNub0jA+1yIz9ZNM3wiquGSXAnBVYcNNGlkNN7i8pr
0lXi9ipr9NDlPAo7sLCj7asBMejSMbhy1mT16cHlLzWB/snIwXCCso1cCwZA4AX1KLCbIuQSGL9P
ONsIG4X8ZlgUq/TxLx5k6+0KsdKAqKjUnqURPFIK9yGovE+USDtwcEmGmXs3ZsUzOS7FLgmRsajj
lyltRjR0ImFboJNCfvcfmeHRYCHwpFgYYF4HcMoF2Wih9DDpNa2cUWajzasCNa4zGXitEYCSIiPh
pWaUddG3t6dYwIVySgge2LuHxk3YR6k111bN+b8KVF0rCYsC6NqxYm6r8kWYe/aEiNExDORY8nX6
eP92dQuU6R0QkHTAms73I5ZLDnDNAvq1oKBmVreHP2OezYmDjGSah3W9PYHSweWu5i5g/84EJZbA
hJgyeY+X1ED4ibKZxaGcIYSYf8yoGvsPwjR/a85n9N8hGvjjSEXuaOKMPTjwVdmJ2KNKHRPXaPKb
AWnJmKsmc572BJa10jvZmsF0vHAQRX5akoShUkai9SCCJCQGZQTlkw6I5Ay35oFt0C0lrPZ1Hjrv
l9Kfm9C2wPb1iITTqVMvP7QguWIu/cSskr+rR0EnA2bNH38/6PHsE0umu+mGusecMh8Pq5GUodof
BsIzBHHknKra5r7+DmLfw1Dg1t0rmx6cOCiJ/0XKN5YSyXWM+TW5YmFmkm03CBvUKkgdnwFneMhB
T/9V0iJJwuW0SdWtS9o9a70o3qzpnaHTOdrFwHDhTgiHt/HG1JX+QqOeak+PjWLaGuNAvV5ZehWR
1gMkHJzUmDUrepYAMHvuJijoiGihgvflTozjFK5adJ7s65TzT1Ac5UKn38aboXBzqLRPl5/O6dgX
q3qRJxMUp9SPNJ0zQcKZTNTDgSzsZIXl0DwD8f5UT1e2vzQgvCPrpCB1L6uodUje5fJI8ruEpcHA
+aw/IT0hEzETYaQfkosJlbwuLzj+J3/Zyh346huTR2Xg7x/SHuyFq3cZ6yFkE2cvzaTeHgozGC2t
R2288pkxkIVhEV/ZB5G08ZF4mL8jV+Kv/I7tye33rGk0KI/kborTkEoOyR0Qhe6PXNEiJ0MF6qfg
RpsOap/HROoS1Qh8WXPV4l25NmD3yr5XLl4JWIDFS+w+ZSr0VYG8I+c9VQ3C+ta7iJflU4sS/PHM
Pccgl7JL9e2rQU5/09fufdsO5c2+fGB3ZX9nP30aZ6Xbln/CC2d9vQBE+Nbj2DQGX4vUOh9+MZMk
tmHMqotorZ5nYfq8F0VtCwx0WylDVsGv8yzG85U6iBM+aET+jkbiYdwCDIl4+JGq4ToqPOONAEUY
3XmQntMg3j8Z/7VUrdCAacyjuKhRQsK4NHj4Tqu2EwxDpVPAA0vfQtzl+r9rQiTNX42lpAZrJhnO
laXOFQEX1NESNdSmQEjpeZTobZYxCNGOLFShAE+Zab4j2M398X7evjnOUzVgs9dN58EBuZlnH5WO
aosea5nbUVAzHa92YICAsl3PxqhkBAJPqoHtPZjz09NEeZTOu7YgiLpNQAQVeUbobFOVcYIx6a9T
HMyuYmTLuvdRXg7thtKvDH43Ror9XFuiM/gUqlLoa3hl78AAUil7bgdy8PDCeUDdNGb9BG2E5QDH
RFlGVjF1OOpX5A37GIpf35KEigFP9IEMBoR7iwbdVErLXXaxFflxrj1QuMaiHsKyua82VJdh1XLc
p1qcqTo9X/errFfo38SE06VxkA8c2CqOKEjxSIl/RvROa44R6mOiSWbi5xdt6DAETKpXVeYbfyez
auhZCTm07cxKgmGgtHbC9UZPHQQUR+d/a7HCVwsDhU8/yVU1uoxyZ9r5JTdKp3YHK76o7gOOR8GX
5NtFNQJtdJJxfZ7wWfj0nv/zgEix4XedXhFH1ga9LdGS1h92xGxRAsG7ag0dYxr2OFQKz1f84dq/
+CaVsy7U9sl4QBaUAcGIXFN72FTa6IQR7AWy7KY9Kzn/bWRie/X+LOMyBESlhxjukMvRPcZvsNsd
Z3wuCvJPYTOkUEuIMSy2exuUOTA2DEZelZZgQH7jYki/uuSxxh3u7/IKbFQ1gQE7QL/roDW48zSF
mLOe1u4bkd8ky9xO0m5a1+LIHqv2yiT/OxcgFIhgJJlhGow1nrSsOd1UBi4pSwx4+U1D7ZjY/u29
iUZRNATlTJyoVscOiv70oZyshNTf8CoJCOgB8EIDQZUt//jrlRzmo9OY1mwfdRr6gTLlIUSnypMs
ETVSi9QLAmphsYhb2vVK5iszMlUeIeVnfVZEKz8Ip/FalcowZqh6JvzhDSnrOoeFB7uIRd4R8VN2
V/amFUUPEedu763AAq5iWNpJ4Dm9eD8pSaI+oEBGcgvGwJwUk6ifB/kuFy7bFXHTUPJvP2uBxjNy
66G206sxABxTXLvENWudxq8Rw3idsxyLIiC4znLiWvTdFWIFUbj52mf3b3+pvbMimSXB7I0H3oc+
D49WbCVhJMmpaM7TKZbp0aFsNSD8v911eU/ODENa6LxwX7OnOCYiGGfgUp0ZrG4n8S3jPRrNbF2f
FhhiyftFWkm9xRcK3baRgs6WS88p6wAdVlFXDsOpmMQMzBVY8m84iRLwZItXCusxBIQE6OHapIBE
6W7q4YgsxuZUY7ZbFFMbiyVCJ4P18tLuBz0robCxJadgtPZ4yyl+OiU3KeXEJ7VkKxwfkl8U/WWr
pCp9ldKnES/1PqODYB48IxaTocHEwwLTqm57/X9XBdwTTwg61hhc50Ij8LLApFzJzeE3wKJYUUt5
2UHwISpZaIAyWuhgDrdmshmYs2qXsq3zQxZlo0BMuV6pCELT1HxD5e1xfdRym6Et+qZrFaZCy35d
FAOnnp4+heAOcXRVGiMgmyTyGBZV2tiqf4JRF0s8mP03X/rRkVUOygq9uaSO1CZzXXVkkxnGBTPM
SxeoryuNJeK5OMnNMuFCMBSXnX1as5o5jgVKm1KCg1i1FY5W451lU3OfRzYlyIXf0JrEvBiTKuLq
obqt/mOvlEV+E/PDygicms1LA/n1q8E8opJbOV+8L+/iRSvYt4Rk/S1mbvoWWQCYVVq7F5bZi4cv
USx7en76osAHmjjdEuPsPwvhUX5d2r5ea5Xo7x0YunVA0kYfQdnJI7MH3/HBTrLR/7dSvtVnEEgz
nmbWEsJEyew+edo7JBkwRppKGvkKMZ3iHP4Hg2zi7E3yvPhhxmI+Dn8egQ+i08MsyOahPtNGavd3
QN31HiZdh7SAfn1Tld1FhcCpq4SY2Wm1xZhtphCopkDaHixhSX/mW90lQ8fzCR0pY/cRrJ5w7e4X
FWfNJuheSe4cCppAsxvcndWdLZxC0N7qgXq2uWJv9ti3MzObKYJ62itsPwQ/vGFnwGyw42hgDUrn
lRLELabMNHv9CUMdwJmwj3TDt7Yv80Ik1D8N4Zijn9/cxNpOlORTf8N+c7GR6ib9HHLyYagDWdxP
v0H/5pC5Yj82p2FTwIOY+Yz0xP+sF094CDB+wizLxh8RlhBBbq2bSpqxRSVwEmR1DZGbY+7mkHGz
UEOgVw229y9R7mq4XBmb4jelSZSqQwus0asapVSl6vagTmiELQ/envC2rYX6Gyl4ay7aMGogEjOW
jDAh39G52GHjUWaHJzM5/bjMyIdTAUlcWy1RC7JbrxLUCEwlqdW+9juhOmJKweA5JDX3uzjSa7Rx
udkquT9DJRVulanbYWs/UBFMQrNCgFmSzW2SupxHwepLU9qVAmB6H2tfLfBqGwwbXu1Qq6RPRMc8
D1oPZE8HdHCMXizz7iIN772tAtocQehqM7WeCR+ay3F+skiIx88jj4DQmhWHmCPkvrj9+kntda0l
P61hZOtrMegBOC7bKZQ+zpYlnSpEwjxhqZkbYPo+BXviJPnhL+yhSt88nZk1KeGGO7h55PxF/3b7
sua5fu7skhNJvFTreNxL0K2Hay0sEqrQtI6Gv9YwntB1nEWIxqswHdLEQuuvOQ+NdE5Dk5/4qt4E
qDIwIZdZMDls2PquKdT3/wSTtqk3yJzRiqjyZ/w3plz7QtfJGvqR/wIveIKAjr6vzV4T2vQRmuKJ
egYOkkbFXtweIyjqiWA1tjiVgJP3D4tMqMp5nQY+dB6sh1ZQMFOvbvHTctNNVGW6cSiwQG7O5wIs
AnPurgSIPnoqJEYTejCwQy5UqVgAOLMWzkQwZr5KCD2JO3VaJNmS43ZHCG7hbCWTegDupofl6OTG
KoqcWqD+CkXnZofNTzgJOMYO6r9Fnk/1W3Zk00YF9oDmnSRyzp4qapTEyJc1Vw0AVkkvfGbFiQWM
pKoQTqKZ7a0U1FtvLV/sT5zNbgjc2w+xUCMIEvMWXHFhpLN4uIYfWt90STwYQZACWHYx/nqhhljL
/OoOLeFvnQ3nMsGZ3wp3zqzmseD+vK6HgfPcz+PxhsSc/rliE4ihNa97M/jg9F0zKKa4cM28XU0v
1qW0XYX2KQ3MO2U2nf0gT8FcTRBmd+bT9eDy7gNlU6UFrkecnjIgaao1Lr88DdAAGBmfwv5KWJ+D
q+WOHKfxGyuKwLJQ1rrwjGVYjHYRsIcOKC3jo0+U3wuQlncUjzaTzrEO6R1/u2MCKukpDEB3ZcDO
NYew792EADdNiTj2pflj/Pq942wJ2ZDtQDEBflYdVApaBpe4xnOX2f2u4Aut0NtqyNMrJAm2FEsg
BCpViDb7YknZhCJbseYBDNrLSTEt5svsrYQjsuuo9VOuJ1AVR4iO3xPgkfQtE1Dm4wcr3xf0vq3q
Ate5ZRMhmIGmGvNXcg5R4GFtySJRF6u3wK94Q7wPlBDrjwXpnADeXlD20Ra66pjnQXm+NCRFkZ+U
xW+iM+SRUHb6OhDWqwGFoHn2zfNyzfdaMl4yK/5r+C8xC+PfqRiKLLYRsQUTGI5k9GE7fK0FSR7s
it8MOXZOqEJ2WkDA9TznQQbHU5cryapQE6mBR2VJxZowtICXDebFeIqjdVcx9dzSz8UXaZiZO6bH
e6z9xotDyRAH+Nocs2q8oefojYj8ypHKgzThz7sU3c6ir+yUg70+N54QhRyuCAQaWonK5pWiT5fM
9JwzhIQm6E6EHz9ZpnqcUzSXKqikiW98i3Ntky7bZeDoFDPLZBnjuPozTU1K7I3aFmjCJEcUVS3u
IfB+rJtqf9psMCoenFWxaSnC3Raj9Z4Z825gVAFQu2tppNEcevQctif4lPCZHnAdmBbmGHR6SGtQ
vph+b5cNfF5CyEfOksWE4swNe6pRCtM5h2Q7kw8FtO7LlXVzcDUucVczGgxdI4dmWFPjTvu5Afpn
Db2eXth9YaSgp9L7VajL8J8JL8UlUNl5spoT6/ARrNfOWWf6AdTiPUGQW9399X5Br4uwl7K58/pl
rdvyp0YD/OfcjMx8qKLwOYhooW9cSQtOCTvovPTtjUgYPggvJNF9WB9uztOt6rJk/rXK9aObtssR
v9EHQMyn6FWnTd9xiK7wp6jaLNFADZtI7iFjLgxufRHigFebY8X+tVWgZNMdp9Ms8JV9XMQmu8Re
CER18tCC3104dGDWVsCXwwhkBh1Pumv8Y2Y2R3h6oLC4PI1OZrhp8/QEk+f5iY8zVYz7eg7b9OD0
oA0JJlBbZZX1hZVRr5e+QxbjhDQPEeTGVOPixBpwVvuxVCzt61LalpBKITVDxUzn3Olvny8phydr
c1dqQLj0n3ST9XZv/Ks1yoOPCyFhce+X+KFbYlKpxCid3x3w+HQ7iseUgP2IOQ3/vpwB1mkHxHwg
wG+ppy9oROfJaJayEXpI5CzfiuKG8YPCcLtLBNJns75ej9vyZyKOkkC+Pm47ey1ARfB8z6J9nyoV
tT5V9431pBnGzBL5EuLkX7hr/AJdfKRl2DzIDGGRnQuIplHt5i/R5Quptl561PH0fr4Yx/FO+RbL
lNVNJ5f0ybf2RDXn6XmslkJ/Mdb9JI81pwEHSuuzfHAa338MAQtcuzYkKpSEWEepQPMyGYQr6536
nGIdWT+NNZikde2Z52VfPwRnumGOi2R062ZUjtnNT1QnKlWyGQg6ME/WMNkes/WIx7y2lEvS+mQA
v82vLQ/ucjVUGJ8K+qeIkS3uZ7l9wigjOAkbKqiKyzW4edGLxMDvyjCUZ6OSVOcJYD3w3yCaHClr
OPqy7FXC5a+TyeZJ1PMX4UVhff+VCoi7jZVvtE5RsFrbQy6ftcXD9hO+SVN/SksD60p3Qb3+qo1M
1H9Yr9MmJ0tzFiSr/XRCHN4OHa3OayudqDTnY2Om5ftlE7IpbTLbUQnQW51Av0AcfWyp87BOWFYq
kfZ1LBqpvqIzEyDHDdk9a/PsSkrIsYMkDeC2WdhwvZmQ2/rj64Z/DPFRLQ/8grOZyqX2enoih9Nb
zK5HifwNzjzrZnGYO77D97LnYUkG8F6HOQUu3t/wFUf7s+eCcukw+dofxxaRdtScvUoPx5s860tC
F2KQAFzbyIN7LMazeNQgYJqcnm7kNBcKm9tGjV1agoDJbTJ3LddcjTK/15HP+KXZY+QmRX0qWMU/
4ucbJpJ75EBwl7LTYe3OWqU/8XI34lfmxVMOjwBvjv0NIEO4R5dXrIsk6p/3NCwf6rFBlq6bGBM7
xyW6iTigAKNr6uuCaO7mCr9JBAJzercEMzNK1wiW4ptSohcpcaBZV52Pf/7E3w17B2F28rNzFggi
sTKvABRVudICv/C9CdtvdOTTMx/x6FA9YKpgR0rgi/BiOxDA+/XuSxuhy6/Mg09NzqnuuHKdDD5P
pRm0dm7+QXJg0xGqy2aluApFSh/Tvncp5cP2P7CmZnF4x/c2QAS7qIhZHIPtnZYKkhkGXPFyhN7H
5IQygyDL1BmOXryMXMO8GD6OHOzyK0y2pxCKuFQnVMxPXi/jSBo3itLg18DfPJRCph+g+krq76ax
j8PFUnf+UqVXJ7BzJ7vTxbJTwx7TH4sgJmvFr+CPHtMiflm6opRq+c2tUDg3vFuaPJogbIp0VTrK
5fbMikhmn2WLrR/VuNRBXH3v8juKFSpr4MGMH2SsYdg01IJntM21XFOokO6crVLFml5EV6ipG19l
NL+ON2up67rRRWgi++AdbteFFoZhgk4klJ5Pa4ALKplRAlVpUTAiPp4QNr6yhRTSrsR3VrYmrnnP
PPBY6lYieGOHDfVZ2xN2fSMHXs3LslV95orsLl1NaX32rB02sF66H9tCNVx3SQGVh456siVGecdd
VjRjrz5OYEYbFOyI76MVzleCQWF9niErHFQrAf/7ipsVgUkNWt25CfI2b1q+tPELihnwkIxY0Dgv
dtEsIUb17aGKLfHzWaTwZ/isOx3ACroevJyzcgLztOLioAImMdJPtnmUt1Wl0uxrrVBsxE2t9lps
SyNzCT7mc/98EOYNZjNsOqqtP/zzesaNrqFr8lip/1mXcfmnygAFh6V1y+9eOronNk+jITkZyFXR
NzecK4TUxuzicpyQcwYalntBaxGz8ps6ZDXgvcBVQAOeXSYQDvyZOfL1NF/otGjfCWOSfS/2j4qw
7U89YkMCx9/Qp8EAY1nlX8qc20aaK2w1yB8Ma5FY6A0tXHm+4a7f+lfKw0K+YFm86izGlue96O3z
JyP5P6ZcLK4a+ks3eqIFFou/re012k+uGcnOSzN+YuD1oq9co8mFVrbHgRlvhyxxFKfClT3LQfZM
uDwXrjVeR8vSmBKsMg+GiMelRkKA91oZ7lz+URyJufEzEEz3qsAV89nyjKmYikNoSXPZyNkwr0aH
8ByBbeJtlx2wjUA8/pZUzBXgKDoNxWSxcb2EW8/1I6hgKiueTKPTXbCszuKx2yWF1d+5L4fjaEvj
RP3eju333tWfTvac/bPVcbBNJmM0jeSjfpkrZSaJLxZjutoYSNvRM6xKvWQpaezLrA44+SzUKAqa
lDNahpEReznEwSevZACKhwwVqcg1XxZZsYkUpsKnr/yHEg/xOn+nuwkxkzOSR0BTUliAR29UyC1L
W2+07Bb0O+NyP9dOQ1c6DMY7QCeP4SSLNx28+UlRwneuQNvro6it28gTzrbKNHuEd0nqWG54pvfI
WP5pDEKTLQ93feAPf/claCuGE8zIjyVpTOSsjqLetAb+11LVXV43gngBmmII/SUK+zc+JaUfqaOM
rVDmrSHzd+jFubaDLxPuupvLlgzCEOD/NfylPIAnrVYe1o3kIGfKfxYBiMh1AhExpGcD8Z5DGdMb
gRCN08FeDz71RjJSYfo2DMJ27Vh2XyYH0OTkKcJt+8NYgiUlOH9bZlxGwqRVEMlvG65xquazY7JO
RGcMLs3YPhd3w5nh1MpCbHYZyQSbNTyuBbPDr2/tCD4Y4L+hyXUFQOna8aNDEX5sKcy8bEYgKu4U
2B0RDoXIflJSpybvZ/b4xcrx/9xZElDDSD8SWbdSq6mMz8iyBu1obxeoqjG75W7hoyEJeGdnzFA7
o5dzYACcveQjui9G8RbekFhqwD3ZFCE/Av8bqfebsEweVWx/PoHulKqi+y3lESH8QuKUdQ/E5qD5
nR7+lcl3bXQDDfNRHIuWVTzyxbSwgi0bjYL8SCn/1WyxyRsfi8rV6YwGqEahAREPHckKFHnywPUN
gjdNuFc/MOYNJ0iI9n97+hZPSAukaEkY5Y4JkhF4l5OWOIFFhxUgqcz4Kd2+mzYFwTrSKGwqZrLw
rDlXO2ECUUIOV6o3BJ0njIMarYZAUj+PCu9/UE53JAuMoLvflpwAFTI8FVAvNwSMZRBZRP7YlULD
KjJcmBJxpCmvC5e/TZKbcb2sLFK6vySZIThDmCyjq011wL3qbhIM8tV3KBWNcvy6wAKnKI3TRC5l
7r1eLFM9+bcDyBJ4AAzpBXL39ukJErs+1YYb1+6FcHKIEtmeEM4GT/PWIR9lEsvhariu0U2scPOZ
7/gr09IMq7IGYeAvDekPNh+6gKt3pCvi9zrM53xZmmeRBv3/D6kyQ1onkQzIXiliyuj7rVUMZtdW
HM0HVvqUzy5fwipr0e+g5S8wM4Opu+9fmRF/XG/GlhvfUQGmRqR53UTJ2cPCgX/RH/TI265zT89C
h9Fq2mrcrxYeukjHKm45Ld+UarsxD3aQc2ejZaxIcwCkVNpyKCdapGV3UlL0X7ppqBPjqTL2rGbp
1laoqw0D1TAKHgHDgABeEfphl+D4+aRUueKmIhXW+qCFCq3aLGOI1pFeccWN91dkqj7vfgVZ5Gxg
69YRWDbQrsRdiffrVordIka6Wx4xiRHnwFYRiD//jLbRP5xz8cOW36oN8yFzodbf73vbdZhEChhU
0JHhSYMrCbwzqUMXBHpz6aIAhieIoDOSrGsv0EmGN1zIOQuKNP5eQ6L8EuiAGcwsMt4LbDDMfdxV
GC2FMPwCpUMxedCGPERt/A6SRMTkLulWloRQHY2YPl6UgOFIp0kH5ftUpqlbUMBYuGdXU5u6T2mI
r82oTe9HLZe0ld2rOzLI2tDg7BSVNp0IGUr3g83iPclaI3RuX0/4oJJSomAUf4lt1lhhkWUrK69V
oKcx5ebgJBSW8MDR1Gi5WMjnB3SW4JeQSC96Yxnept0d5nRv3EadVG9QlKyNj6GjxNtc928guRex
AGJDKZVOP4toLJSF8AKnnuvUN8fXoJ/L4+cMHF5RWrGPpVTK5KY8/CtlIDRD5ke5l1XcnC/rMcFe
J4hnbj+bbCzrkDLABKOgLpd6Mk8PwUZrLqXoZnESNXxhKyYCeOw/qS4+0QoOuw4ePxqxUizhLM3u
SgKx8LmDll6eLCMNu/agNxvhnHnRTvZIRyUCEwPp3y3QjKybaX+UB1bJqULmLbDPO3h125iY1zf3
cJFw+Ful31m2GWETzx/I4QMyiGw9Tjvx/z2tFWr9DAjxqqQGkZYQUczIgW1Pmh6pD35EcyNIq+HO
dZls4rngiOXBBnENYhB9/xsv8ot8+YUfgBnLyk5JtOyYxlm3tPdw35OeivzdtioNC7pfKhFlPTf6
KdtivyOy3wGKovXr7WLLa/SJoUMepqVbmeoDuSPnNGP8/RVZfQjWbueV+Yr5X4MlWYpaqKlINNn8
8LYfzZk/d7j1V+zyskIyGmCaQIQgP1QIUVxGtlP0+z6SJElU12g8mmyfymfE/DwXHU6FACcFHYJr
CHdTEEqisoatwXfkOPhXhBRzIerSNZe3JSd0B61hknmRgEuduXl0pryc1pH3+D26EAHODBnaIr5x
QHyuMoJCGC+bf/mOSVdAtHW5uK/lKdmQEFrK6L09vS6ymoKwID5QFldpUjgH3NK9URvnk9mTANJB
Zi+Y2cScN3u9Cxs4PTHwqtMElI4yVWdER36KH1/eG6ue+Az/1HxrCjDnBgceIhGByDPZdFrEh8X8
kN0lAeCJacu2IQwNs5tk9ZGGw+NbDiUX3B5rXemU/GmDPMT5o3wnNulgyabDEGMkw6BQRmhrvw2g
II3rHptW80p4/zEyZXZ9+0vIzAhPhdgL7LfZdPDym3ryAR3X33V6GJ6S9FFEmFivuIgo+UIldAbj
YISeJKGcvchRTuNcegNKUlD38jJyG3VZ89W6mmH3FalpcPV02hAPv7Ol8CyuqKKs/upgZ2jx0X+J
z0ozUUVa7hf9cHeyVzhCgSl0jSmQ1Gj72SkAIBQwRPGOHW5cDb25arfHrkX4td33SYoxzlSznbua
TWL6DESq5v2kGwJi+8MlLIhBvnOCOD/J0boBAEc8z+mamtMeoibk8lRK8V3uwHhM8+YqUXZcGows
ZhGsmtr8BFZ2sopQ6CCYQsEB2UAxKwdUmycAlVcD80PGz9kj8AGMOM2G6m4/tAVsK4K/zmm8VLZY
YOKhi2rZfOOA3QMHznGsjroz0MEkBvn2ynfIV1rziQJ/X+VorTNE5q+3I0i31b2SoEPS8hK9HSCn
Qjc4HRXBdkRpZIZyBBuc2zKX9e9TCzlyjrRN9d4oLGr+XmW2OTY1hd3XPigC68nymGsRn1p0jAiQ
89Bf8dATkvpKekKhOrvq3plqf78VXis8zLdJJIzcfP7+4GxdPnqqaEp6FwXRZxhyKio6KqoeWq/7
2fYio+j4i0GpENN6SEtfIPzx+RSJuWCpJJrzanldF2FPwzScJW+qMQTtku6b0D7xri1cAhsLILzt
RE6SJXXY6Myt8BAtjvFaPJdj76k5HcDI0VkBGxMpevUD5BcI6/ddmAuHGK/VPtN0BB43Rvwjgds2
rzbTf8vo/31avo51bOMyCFsobO+i0D488hJNTucbCsLqVImeJ81iDBx7lS3yD9I8EsrGgN/32LmZ
u8CG0ruav3Id7cChdaT2EWMCosU+5L6XmXb+R1J2PuMz5/I6tJOA9+W9LwhffKwfMivoG/upvV9w
LOjIVmgKKMqVy8ujYIYHPpJlN9OQSdUhH0VaW+q+rG/YRnQfGC3p5J8tYjAG40G/LnPRY1LE6A/f
2TctDWo1prp34CUloXjKisesAZRGkTXNSokxjpNtKjlLn0XvfABNMzyzRDyvhlIaMW4h2dDj/IdY
9DrR5+pxv4Zj+xW/jF/8lACxx+lL8z4vtVZiA1EqO0L8ftOFJFDanzu4UTdD0ClOQJ+Q76Y54B8R
S1lTxGMX4zj6S07ynuMe8NL5xFIB8PG3nZTbAyKajwEbapr8BOfgvfPzSB2XxIc589nTyBfoRGR9
oqPjTeRviATII+7UwjdJtT4AylTiGZlnGggftpp2ZCtcnxCu0S88eYmO9K39eONENdNvZmOLZL9B
T6vyXZ4jh6t8P3YncNmWfHKeJDq1OV3qU9xaJRRI8hPtvizttnuZVSXW2Tat/NQNUrViUuv8yApK
9a61UCJirNqa7pKYyRmyG3QCphZcxaxq4tsvhxWSfryaQQSd90e3Cd15R/30rUYg2KOBu6Fcyz2g
+SgJ565g51nVq99E3Q2B65ULPVMLqlaYCHxr+nPhtlvRgjgpLxnlUcKejLH5RIGDhkjLNo1L10Th
cHoI8JVmEEiboi5+ojMUe3ikD5/jwroxg4LQX+WPZXctPIvpHFI7/5pE5jRP9kXcC/sYseI8DNya
Y3rOqC/86u/Ar4w8xYP/lSfsB21DPbA8dG/fe1tSXl6ERoQYA8Q5dWA33rFI1VPibn9/pZA8k8xQ
TnJieiixxLVK7g/PzU87ondjqysZDLeYx04tgKWWazrulITLF7lHVU+rsA/g7S7DhWCXdfAWL3tk
6a1FTHzRUwXbbwIN9IUF2Gb8uc0wgMNJzWshKLn2AjwJEqm1+XfdP2nwWuMopnqx4AK9xXFasbpH
CmFwMxBM7GrTFAjt5b0IvwxFSs0NxNZxISHCNthd+ck+yJE3gGirmSS8GqxZYEPR4195sieAt+g5
MweOHNSye+Zeds0etwNo0wHKwwATlvvq/wNQr4c9X2iOlugh60Og2j69dag4V03nvh450hIIgyV8
1ViQQQ/5FrQENLwKYw9LovJsp6v9bJc5ZEzwcrmM6gl9gsabLK7pHB76VJN6GXWrCUj3rEs9BvpI
A9d3Lf5HDimmQl1eHjKNu9oodONahIQR+tdtUixj12laXPPHknKkJruzxkb3qX95gsaBULg3Reuj
PKNJpwJNxWHOrA1msTXINxGVkyJnvdEAQkOxQ0KLq7U8IWSXMhvEnz/gpzv0dApgA08gBM51dX10
vKXq7cGLPLGc5SzqMoTypSrbaye8y9HjbkAHhnrO6ahYMajSmq4DozBQbjZdy21NmydOguMFbeqw
t5J9pyLNgbG0pDI7njAHi3qHYQqfqN1FcXxgy9dch5veksvh7Oj1a7ooyVfKPSZyEUi9gSkTk3H+
uS0qFrgdzzeuby4NcEqpeJlP15GK8EniuLYuMw5v0qY44UJwreY9+EJSDnRmEjo0xooNqLg/I+n/
xn1JZlzbXvnHzuP+5KH3VBCDNO6fUOnMCk5+MT3uTodiH7THFRV3F7/LBK9xFvsffusEAbiIbl3C
Jk5gWjVeE2xEytkzdatL1aDCl5lptJkfSRut5p13VXXNRANKGtJaajY3Giw/aPBIVv/U6k0+si4c
VP9+IDxHnds4yXp20SwPR3ZoEf77NVqGTUCBdTAorIxY2j2D/mYzv/MTBlRdP9tFGfmDxh8B/CIe
tGTc/8Mk4sABDv7H8gjZ5aNhKJxEIOCyk6D8SYty0iyU+aTWy21yP/LVQpC7uCkNOAB58SL8exWA
1LMkolWH/MsSgS5M6MSpRNvUoHs61JPBFa7y3gtynsFFBVN/Cw1yXQYAOsOU4fFus0W3xdrCnuJP
Di70aNWULbmARfu1JMz3HUhU2hCA9O+a6s/6nlCPDOC2v2wiuBzhDcMcCwZefx2FDYENA5Dwle5t
RN6qaE59lGtHffEsd6J30hXbRlAS5caHW2Tw3scurFnURaj43d04Ljc4jLf3alsfzZ3heJzBI6dY
DB9Ze2L3BvzDAPkDfGs8viTdfXHsujzLbO3tWcds1IWTX6/P97vhbMLD+akofnfeHsj80l4CVcQ2
qnQR89LTLYWhAL1ujEHLwNUn+1kQt2JiYK1uvuQCOt3zbslx5blqyU1w5i6kG/s/XQ2GOohDYx04
rl50xIOu7h9kzVinM59Fc6kc1Fk6zUQSPhItJrQuok49rJnOaF5YW2FLcgeUCzF+HY8HnIInzywq
eJ5nIxHbQcTHjebpmDAjl43rN1d2lWEnMYeUuyujdfDhUeCXuvT64TaGNmgiqFlDtrkYJvVrs+TC
qswxLXO5tKYUAuSghyRVs3oyj82zawEmxAuoKHCPuUh8VFrFWqbRlFc675qouRk3rt1uG3OwCFAO
cUBB5PxTREFOPb58TCV+HSJV6vxhr47tsrN52oVQrOUgd28crxm9ww5XA1OyOqK0zhZ04PYLcY86
XqrspWbcU4mqqaH/aepDS7NNf+pc+8iEMqNyYaccbnvdB+BOJdk6HUDT0FMayymzk0Uj2907wm/H
ueGbBBcRdg+OaaBOHpwGpamm+fp1GxyBYSEVQyWzOu7s8jWGlTxtLojEdk3Uw1A/NIUf4En9AnJQ
906a0bE4/tdt25NqkRHJUuWpLMRHwXIP6i64+2UdJBwLr93aoNqVr5EdupnYERMFmLioAP3asJF1
CbP3yYZSVD0eR0Lq2wsl0ArG2/SfeFDyTGxLhD2oeEZcXPxFkgPtueBGp3in+aIB/FZD3Hk7ugXU
Y4wkjB9qC+d0cVdD5TkjqJmvGUyUTWiCWU80abpQqKT0FwwL9qohCG7+rqaxQd62RXGDbyaGN21x
5lCbrNZW9/05co0SwYwQDvaNwEl0t4mXe8MGqeAc6Gc9FHgSnlwe80m0FMfTDsX+iIlEx0uenQeL
bwVTAVfYmJua/LgRKxwD+HnIVL2+uvA7O4Do5gtDRyeJfOn9kMIGsa1HZpF21PoQHdklTYIErBQ8
zGlpHlbD+YIi1da5kYALNCoDhQ7bA+hT9LW0qp35sTXhORYgQKobXHJgXKlq2zPjZKYrzLEftG5x
jXFqyR29vFiFhazDou5fQ6yoVwEYweUUGCAmHFaGCNJi3YLnQdPVJQ83/VTPS90Sw1XrZTyOuLYD
krZkAx4acNSHfOr6g9o2rNXZEWxHM+QFMLVXanjcQ3V9rUZSYWdufIzbETStioFH9JV1W7s+hafh
xA45ICxwx5snrRRGSx7QXyZhNLkz34JuXRpIm0wLCPLr5zx6caZeiHD2J5ySC6frQStOqtFKpnTA
4Kq08vQJks7dVHE41nNt01o7q0zL0sSfnwHJBl/hSSkUy22UKEq5RuH9XkvfUwuZgW46Gvjemqwc
XMQdDLZzif2lDL3S4dwdrQKYY3rqJm7mpfQerqs+fg3Ryxt6QHpm1MuG5UMU+7YAVoLTEucorxIH
kkdbaHEvkdITaxI6yvvBOLkep6DT3e/gLerdPDJDohBTNY87306W3MeaSeiv5Sd971RZkRNI3X8K
tvwCdswmXD12fQS3bMy85VVXHuH7bV7Q7nAhUbNeNBV/8rRWH49SKJtF8hez6kyFHrfP5CT+0Hyy
ZhkyFLIBalp9Mq/1TD0oTZvfMy69rCCLWXxflvDV0/r9FlzAXxcZZECTtPOlMuNJrBQAFrRZeni9
c643LwjJbRJZuWCn5GkDAuDq24HitkUVuNJD5taQOy1m8KgyhT7VAJmoE7rRwpRC5nZfCxwYecAl
CoFyYxi1brOYVtSJjDCrgCmUEaaWUKI8kupluFEss84lvi4yaf9tjBBoA6lcPqN0tGTkoCChgTtc
L4UVGlLxSMnvecjdAofvPtDDEUqZQoNak6NCVafsQblVZpVn77wxFNhG3kcP9yfMoUYtlsZFH1DZ
vwSbbox0mdFHpJFj+65aon6/RgrO5F+hb62n/aT+q9vqf/S+obkqDOXp/n4qxl/H/rnNq23Mzooc
yVAaf9Mv0ThONjcZ8RBAdBBdyD8f8fbu9rPU45qMHDpZ7PZ244L/u3YWDK11C6aKY1HQIem1hC8A
x5pPOAM8Ir81OdSLbfpPcXcXupTeksiC+ccVt6q5zN8C5HigXx2GKfRJNU5jq3hQ8EBEsQscGM/j
Lm3DeBYK47ePhs/bT5TWp5sF6qglhHki5PuGLdXL+ftnZD+zIAFDoQ2As4e0QecJubTgNTyw2kbK
W8TQDwDv8+f0jXFcDBrDiCILz5cPYya/qwR2uwUV7Q9ReaDdmOiXLJICs8pmiyjV3/4H9dcivRct
rjLRWRVlfh2098MiaFUO0ceky90eHRIrp5GTHPBeUe/xuByG+DTJmO9XUtvUMgwzkEr0pTRpUBrf
JqawtjTajVrv4pr/ogeKWFOavsmG/u5RgGt/g097YWfzbDuQh60StEh/rtWAjtxiEfzzTC3k0mT0
BCzcE2kbYqOFd6y1kJ58oqgFcLxYuS4fwZxVBqfoxPiGWXMSYEljEJf/Mv8ZfyS28vwk0Hn1vdFr
XZaDqtJN6LeEQw/CjvKfQD57ISdXl4AiMvTAQdYH4IFPCQzIXqminSgGl5j3pw4oSggWk+f2zuuh
4R7EAKKtnHFwY1m3mtC77JvwHVoOK9rm1Vn/iRqd7QnENQbSUffzfxCpkDpAhP0De9xE6faggNw7
NTc6rfHdRLTmopd+Ybqp7ZTxirJiWENGDav4VL8GkPIsxvNFu8l1tTQV0f+CeGS9/2rQ8J0KfvAQ
LQ5i70ojsIMsdsmQ3AWNlHWAWFiLrjmTFkGArDivoeS5h9qcwoDUMv/e53NPzQwCJaWwKfeuV5lT
3opYQ6drFh2FvDY6wFzD3sHOeF/n/gLTfnHnP3mxJEAUb8aBAIHTkrgHHYX4/5AbSovEbyPFbWOS
d8YlbvZ+mfcj4UA7cGpUzCsP4xfJgaderyh0O0i7ASMNZ23/pBcI4rJBqvL6YtjKKkmLvKd1Am8E
iI3YI1z4l257zs4bXu6qZp2CvmUvih5XFmC+uwyBgoZ9CRU3tWhOeWdYCOAFy1KBJXiXP8+bw4Ca
CpCSjUdaZCdOBJ2qWaKfkDh85D1agL/N5K3DSn2wNnw0ATTPZCV+N5+FBFqD4+0h4Sx30ZAjzxZn
ije4xaspowM9cwgIW8MtYWvWmipDyXErXYp0KYMT1M1o2Q/aXnpcxvhTU99Pf6hd6Q72JCqVboEL
0XrLuHJnJ+H2A2wAJhzkJB8Mp7gfBE1IoJFodEKpZibavFkHWgfBHERVQBrD5fbKEzPbGUs/GHcU
cdvMdYG9J1Tf7WN7fSVPhnA9kIned6LQB10yS4bVUcOmfMkbjWPOQbl3A4AqIFy2alUDTcqBp+hj
F/iZ1+ZGGwx1do8WheFN50ZsGZ/MR3ReP4Lmvg/MU+jW7NzDK592lFy5HFcL8/ITOHJA9X016WOm
79jQ2Q8QjhDPJ+Cx8kdtR3g2z13/M05BrSoCd7+crDUl1HuN3LkEqxxyH54RqXvYPJVkGQj26H18
0Yfzk64H1bOiyom1VMT/pnJE3qIQPL51cfZj9ltALki428Fdwk8F6coVpCrcjcvwkh7Q0HtSdHVD
p70Ed8eaCA1Hxxp2Tb4QuNOsfWWic191kIVrQTnh7crjOpCtUIB2pGgckBGXlNkP5xcKBFhdgpPS
9lw6ljs6/ITo+P1+8SinmrTumyonAYtfTNt31m2EpTX0s1fPcr8WxEFj7Oh9fMD6WNuMPcisCkK0
bG97iejcby7mGU4V08jdxwigztLGXjKlebf0+EIZODpLnACi8fhwVCuiuks0qS1rfQry/9FNW9VJ
sXkfidA3CakDoXYgjHCI9PoSTJczrM1hvfZATyg2+c+XUkz1xAldxQec3JIXKW2jMm2RwxdVYQqg
yRvwTCTZ33YTg9BL3N2jmLSAXoqvtBnIH9d53h3IcRHjHMRAMtl7M33eIHXtGNMktCJkqKeZjXAW
jrY8qGMm2YlXonni+eclP2H+q4gGKXilOioWJdp/VvhBWoucmPj0Qofx+dlhY6TX+WKTzDjjDf8t
mi8hMTIvGthIE1vbTZGJvQP8xoIC1s3hfDK7dMznGH+Gu9wKTBi+ZWOrs//9buGrtuUWZDwJ8I2V
OW+zuO3+opyZSfjni0ZmL6IAJrxM2scYXljxhJl7xSd7iSzcRS4ERV4jz4Jc+Y0q1qecF9h73Fnx
pD1GrwuE9EN/sZmiY4ER40xnQH0jPfmt3ZPIpGnxlTWhMBF/mTSAPMCL6/6Yg18uKJbaMVJDPOKW
qxRMAMrclRWipKOFkV/1aOZLafMj5KdYApJgdKJBrpcwLmzLLzCKpjAIW/9+wIlk1OoczU2lwWA9
pKZauI/2euSv+O6gtxmzHu7h1eh8ZOcNmlGm4rkTzEho2NnLwfYt/7vwLxrO2B+LoM3mDrWvYzyL
W0UmFaZ9ep/KsPRV0J1gk/d/jX4xTQt99pg/tfe739BsFeL4CAed88Xb00NgLD0gjy32JwH7k1ki
fiLCKrNx4OdnF2ClTR25XA3DuBNYTJuRplIrICmFnmfA86Lwx5hbgtufteq1dAyKHdRVLFLKra9G
ySb28b5HrC8UfnYTPzFRybxVsUkzIl1cU4yTV4t8cdKmZn/rYnf2ByMmZq8S+0FXziHvUj1do700
6jKaIOTnujA13gbrqLTDOOFzV1jobFrz/Di6EU4+TcmouDH3icOx3fXrOzLWDXY3RIDq2QUuQPBm
ZzRAaiLuqxAeLNGnqs5QiJrhvaOysZ58ONKXxtnetz2PnC+rfgEsmjVQ8i7zkmGgRewV/7T0B6VH
cPqDS5jH7bDG737INS12NRQVNp0kNLj5ah0GQlMyFKYhtlYJQBehy5hWQtwM91p3q3ixEqDKZl4S
bd1rQxT9dg1wC/KawG0K+okMoSBTE30HyiWFFV3DiH544FYQIe0yhJlUb8+RnL1K9GKncH7n2TvR
z3YXHxVya7leQO0/A3RvJf6LWjshCmPzdAdR4vQp5EZjQxOAiEyvqxIpfc2LIvyOhdx9UHLy50cI
0hkT9KFD+JQDZHuVwwouBo9GBOpkVERuCJusiikSyAULEiSjncY9IPqBxVVzT7MjfngHNRY3K7P5
gbl6QhCwvhZ7tBa0rO9wUYu1wGq86cWBDA966l063cDuxFSYDl470yhOuuKOL581n0Ezo0+XL17g
3ek5H432E1emAtTTbAnaF0ZaS5H4yoMtKnGYz5Sy5svpnbW+djHg/rEagnJI7OgluLSeC0SJrEVg
WV5POtGxI+rcO4ydxTKfCOwDbZfbW+6qyX2FHkx+t0LIZW0zGwzGu0dHsHqv5bpSgSNuHe0x6GeV
rqTGQEg1z5Ne4RM56OsKiXOje/hn8a06GYl3NBdpIiSJMx5OkS3wAwu9wdZRX2scWtDIOdeYs/4t
Tfx00RNh/yLYwucgIFGaubWVVFAqoivxtK4lZdAY2pm90/+nk/8wDj1ampvf3PITiA7C2i0pvPJh
NfNxUki0LVzwozmDQ/BUH8VG4zT6sIcvOmf75PBX1achRgQlHQUKJ6nW6Wqq2zlg24CYDssztqih
kfAOtJ6DpK9hxP3avEplYXKGpW9E6ZgCkRbQUsIyE783t0N4foPLH5CMCFjts+Bf/ZdX23kDm7VA
iAtXPRrna4rjSlPmXnn10fnQnge9NBN9jI5tWo7DIpQGj/eyGtwuGZJ04bPaqlFIwoAllLabd7jR
DiiInrC0zdOMxSHEypr1KPJ4cWI1PeCRDDqHW1+mqSaU7L3oSryHSC60vOUqp8NbktVkWl6qfM8M
h6tlTFGh4hBBJCUOLxo2jBG9OeX7weNfX8mKjfN4pm+wa3endJEBp8Q++uR8g5M/BuTYAyyirkRL
wTMVKTydE5He7pzI9hdgSCxbxncdOyLa7XGQ83qljoIh3RilZDWzzE2QjU46ZawNp9OK/caD/i+h
+fa7dSdSeOCCkIrOZLaunloJmUGaGwuH9cIglMqZIZ0ga62/JGyTrclH7cxuLaG4AYYHjnWmldL3
MxjcQw7PMeF8HD0ObyAd89TKJG4I8KMOBYeISE1yEsxbd/lmSnrXQxbexV19hI+11b0iaj+D4DEH
skVrXKQii3Htes6Bmeoy+hWbfAMtpNxt8KEYFzW9dRXpOys3ZWCR94SYmBgVRmocX3M5mF5AikFW
bd9qxZEJlmR47r3rw4rWQHiSMpOcNIqAgBuALok/684VFpMxFU4ggi1mTX0rxby1UEX4lQv+kDf5
XLd2fnh6R/d32Jp/bLQJuZdYMzp+sqRdhQh/raCEr6081A8WlfA1c/qwvP+grJm9iTCtUGDH7HE4
etQ6L5UocRHCL736EcX2YDd7+bYNt0wDhd0aMbK59yq6igOZCWCEi0t+6Z2Qn2j9foIPX9fM4lXw
DwN2u+46wkPzj5YzNJz2CUBK29skeZ6LR0C7/bwMxwkv3PwSsAFNW7+rNbDjk6fgImt8Cnw6avpK
hRojIbm/qO2gZD+MhEmS4SnoVoAG3/zXeAgp3q+VlrtemgjM+Ss5ISzyS63npwyBdRM190M7+fJC
wV3ivpn5/qHB85pvTxWRc+DW0QI+YeQdL08TdGukz/0k6VfdbLmib+Fisr5wOersjc6A92jbAW+I
lWA07YYhy7PqQKxPvdLm0p5N69Qnf5ySyTgyNxs5hFuDcnLgsXx/Pr7muMIGTXJA3uRZvC1LGoTn
SjjqRiRfE+Fr17nhBPVpppLKS/2kw62edsOrrfAvUM1+XUordqJZb7gvlVpRiIfg9E2cuqWgIXHO
BdDp7QxTBhNGsne9QcrZJbEd0vVj7I0m2EyF1KqKumF7fwzlDqBJ/zmUlo62y1luip/CK0cUQ7o7
sdDH86gTSn1y+quAHwPutznmY4QIcOITFXCcpSt5PJCSuZ54C5NJBZO/aAStYVeT4uoY0jDBDBOY
4iwNIiqZ3YAkzrFzLBFTHpRDFdRJloS8MJZjAjQU1NEqxr5vIlnr3Cm6Lh5xXXve7eJKZpYKuu7q
4zmajZGSJeMj8KfsJXmeGW+9dJIQTlUyCI0JHvDZNDqp5VC6QZZTEKyWnIsd9dSwscPaEti7mu9o
dKDiImCAJ0O9gEgBmoAaSHOn/fyvzT9+AW5RVXhC1SCjkrgxWM+VCZ1kxjZbZWGMfPSUFP6xO+kc
LZlK9RioUNrXTHBwTOFtjxP5TgKP3KOC3fA7IU6kkRBA7CyEbPmP+25d4tFo3GSWNgKNWTfzQ0Oq
rTdY/+p5MLsPAPgcsqu3v9lBZvSkT9Ny5xuEee4wVXSTK/TUUb84qW2KDSeNmQFzG0Z2jQy0LoFy
bbI8Vn2k0ys55deT2eg9yxmKi/6QLnOeAsjeS8HhFN3K0ZuplNcrTEcLbAQz4SYCqkvyFASbgqu+
acCxiZCw1uErCYLFNumDjCftz4VoWsjsuwuB3MTqTFS38RZpcpfBpTUUyMedKBtGRpPWncGotKCE
dsnEPd5cc8clVO2ZamtdRszVcrCoYAb6dsvDTpKapbJwLLHAObffNdwHoUgFZ+cY+vjnRYOOQ4fL
SxuCcO5JhD6PpaR1hilUPOTQEpkMHqC02GH5mPsZUjmB8FkgM7j6aIiUmzqz7KesKQwgoHeCk+BB
8NdaARTs4ZFwncaSdJLAEszPHDa8NAXcdsxJ2A3YayKfkXzsuS66OVg/7uChMU/91CLeA+hX0jU8
slYSXQ1f1fn1d4Z3eBWjhNY9jKFo65iJQL3xzF8OtsXQ6tWfeztOW4kH/onuo1vGhfAGE6JntBW1
mYfukoT9knrINkF+9p/TeX8sRTRbuzzE+IvywEOzPK11Np6Ec4f64hijKPPNZrTaE+lS/6rhHENP
qv54mll4C52xddXM66nCy1M7a6bCnZzufQMMt97YPEihDgIHpr9BjCqIQGXapn7GQY9shF0ahKNu
kfheBgUAbiVYFjDERAC0a/pAX2HXuShOjjfhnU50F3TJ16TVmmxgEMHLpJjUBvEHWlic55ygtgvb
SVHar7ldbj/loFoFbXnU2jIAyPoLLkoTtDuLZwJ/6W+LwJHrF06lOCCNKY8bqZa5eUHL1l5+BVWt
pDXQ7sim35QCylcbPfujb7lekbXE2z7bUGsYl9Rx1tTQjCFxPe7A3pepY5C2VKAzkwvpqUum0gO4
WeA+ko+eXgNNNW5CmkiTNS5wNNswz5f5N1JFqDsg3gZvvoD/4vtb6ICWgRlFVFqaLsKkEme9JX/8
QOH+MSny4XfQJ3pwkriHC3Yt7X3ExmXUye7P5i/T/g3eS8sgpp7IDjJ1L79lE1oEHXCQGqHvZZNj
14QThTg/fib26BnRs8b0nlU8fSzO7H+/Feka6eMXtTVu+tRaU0y5OvUaKfhJaUv1F+nhl2df4rfk
9srddREzRrLoYVxMRdMZZN44b+SpFcdvOHZeuIR9IoSlSk1bqk8wSw5Nm+I2Ynxum+fLpSp3jRnF
N48IjV/0NLyVFUg/4b/2oJwPEb8yg3HJtyLqc8D16e0OkH6g8pgmr71+MFUDwZEjlfhT7dq0Vdqq
MhPVJdH8UP8Jn/fGx37OQiPUedPc5LLQvxLIoktWBBfE1t2vmDC7mj9pV/y1Vd1ntiT0qxRuffJd
+dtR48GPmRSJqLGlt9m5cS4VHbbYnaWiXnr11EAiBlyPwCEcQjw+WZkNBnO1V+vHnsyCMYRfvc1U
EcK6hoL+oMsuKPJzRNNGo47ZFS2HAdpAdo1rHYcJ1p2lMrHxcqAXA4fOhkcNBUE/X7RP7ygmNqyR
eIkLKyiywM6U7TMJdLvXV7ygG+ebKcpCEWF+0xOL/g3B3YO0z4FDR0pfPxHH3qmYZnmdTdcEu+Y0
lW9pUAB58JNyEoqmAjxMmBh5WvFBjY0Vp58yyMSC7t42MRZNNKwkgNl/YOeGUegWL/fiQIXtpMkl
Dvl0OpjdW4GfwbZkkydTh4EDtZDZSNAPac915tfSfdbZiJ2bK2WJ7POKBhA8cbCX5yEUimLqsWCt
6lGJZ9KnUGQFd1vtVwv5zrU47t4eVMzhJmcR7w8DoMvLkjXurZGQ82HTnp4laXdkFo/V+s9us7l/
Mj7JC846sRMuY5IQrwIoGeiC1y2AZ/ZBZs5eRoVvh0RKm3uaKXtUzSx1cb+vKK3D+5awEy5Hvyt1
iXxeuZi4sswO7NNqlnNVaio8sE9T1SwmCQprIcAvgTMhIQ0ktDdXCKsh3766yaaI2ZwV936e25lO
ejr7yfNEmNzA6YpnpuF5+f4Wkhc4lUsHiU6jvyqT6MstPDm8/UsF8c7AcdF5ien3UEvn8b9Fee5u
iNlJ+/sXUP690jaLX9z0opM26EfNv4GZOc4oTnSLgbaZEXuchNn8sRCPc2EqrULgGub+pts1du0h
Dz0Z6gF1YyMXvwZ3NJkdO8DhV/kpC1i8WF/J8GRJ4uaFt5b8We8O692KbFn5bpxN4+2BhXavDW9E
kpnHwlSMmcpP6rC5CI5OzuOOTtN/EMXQj55BKLwrG7DCNclUM77los11GGUqdWb3jdMQk5GoC9rH
nG4RGMIarSawiv3aJtuepo39XgW55TaDJxy1IG5NzOImwWjjJDBAghRTc7V6X4Rfh/0jqPBtg9hk
pI+8z8T202x2H3Cq0EybBqMD6+yrOMGfUKcb2O1xn54M8NwoKShOaxyFTr2mhLEno3oCexnyOYM7
lvCXFi2Jyjue2lmT0L9EqQfmKMWa+pYNcUyFSnjxK14ThzTpcS0GaZWVRZp24QL1mfwtk7JWITrE
aDVlGHFUiYYKsnis/lC27RXKS2H69YWe1IGfIQtdllFo1fRK10+bEmwkkRtM/sgYE4GZoVKSU+n9
BLQ5un1v/cJ+QGZa8wFjUyqiLZ8XxmCgzKNTAQjFy+B7dLMoq4bsMYAZQuqrc7r4eplU51j9TxIO
reWkUKcl3Psq1BMl8yuPts4G05T/uFtVODzTm+cgzNyvbuaARyTTpxjhPaeC+AbTHnJsIuJq7IBQ
PETVL3x4z+OtuXJ2qN67nOMjHNo1UheBRsEgLhX8QgnCiBezX8fvL719xqgMWLvEnQjo9+FbsKKn
W8pVlt0euG0qbjU9f5FH1jBej1G1tSv2Ht6R7v7a0MHJx8Z52/rJrxgO3S0vR+gG1Sq7kiqVnJSi
iPPxio0Y1AklaSWyrxXAxzmujha1Zg/9sRTWYxyy5cGIUcL9fAoyDatS4vagJ6J+QArorB3jOo8H
XXwZEayybgfGmV9RzSjL3aLTYvtG6y2WsL+MOxkMSCq/8DAQC16Tv+iM7cS5Uf4yQz4CgzMG/5la
EA6YVaOR4s6XiVvHKNYgCnw5URP7N5c28sUk3SIIcCx+nRrKNps8FTe1Ug7tnw7RBhI4NC/H77fz
JcOePs/npZSONLnSYPfMIAtiwI+nI+AoiHTf9wctWRY5YugrPY8+0rcYssK4ihlUgEtpj2V26pb7
lAKvJ6NpO4QOgJYG7+4r7jXFlCUv8dnFOyly3SYQS843mtwe5WJGzeM9+Ru9STujxN0/ZP92ccpe
4Cr53sJ6iJJAxZJuJfV4xZjFHULFqk8ZrgX6iDIJxmT/d50YBVHejq3KGvO9IG1oG9cYT2HsWP8J
KIVsA2EebsZHXeznUVWd71yToYwRkncqY+YG4vrRvLtTLiPnFKftvVSPImE6lzzvMraW5M2xSXp0
FZRVRYeD3lP8S/uEYEuB168hRFxKr276kXyv6hJotM5ofk5oI2aty5Dia+RAND9NTYXLR/w1nHIn
ex3LlXtkCblMOH3JDpLi9M3lKonSLFKbayo5+Pxqpx+Awx0IrqgiTOHf6I5qsYbV0UQ8A8KRybRn
+6e5kuZbtD1SjFV3MjvAhcNeTEbTHazuotwx/gCcuEqZuFcRp2OfjOPpRh3WllvSvoUPzioleYUx
V8ERZIw4i5Fj7NF7dQ1zpQtXdokn5II7EZTr5lrYA81nW6EWG4wdPtcTRLc0DiQi/jr2u1F0QKT7
nsuGV4eU0ALglaYCPH0SxdZn/AkncT4wJQ5QyAcczaFnwQxuBDpI2cGYvyNp1d9qM+7xEj620HOl
hTMRQeYYvSd7H5nMejujax2SeUyeTD66MtB9F8+My2wF0D0MhKQ6WpniGSXySDFEPD9Dm384zjNG
taBIXHSNEydtFLAI0g0Wk/6dhzQkT0Tx2tIIHBiqWM/JzO0klfkeeenfMw26j74t6pin18vdqg58
J4X0lkWzz9NwDs+K/G2XsMY4ayd6uT9jv5k9Kht0svCYSkV+B1SnL4lfv2ivsI7AGSMnnQMPLOp6
n6JnHPA/6AA8YOdZOMN0f02fiyrQH/C+6Y3H+4JZgzwVq0KTrYwzPUsntwBOEyyDWmhy+pXF05BF
sVc7YsPaXj/MVZkg4offzQrS6VCpIUNcToBlWZFlZF4oV05t8puTg14kP644LeY1Zw3hYxElu/5D
IV2By3PqxL5ij2AdIijtwepMQmkIMovci4C7RQYv3f4fegKjkcs2TxzuOiMBm7IznGSsrLZk26yn
8mJYnfseMZlsasKy107vgNE0h9dtGJryGlZRtlUAc/c6nLXmHf452As778KovY/3E8BQXUrtyZW3
xx+taaRPQ8UVjKtSfUGPZ+CLTYZuDW0N/o8k2WwF0CvQU0jGITFMZR3ub6St8l3PfDfOUK6hqNca
d8LB8tqR1w+iwFxxRs4NWqSa8Iqx78iD1W16p4e6mXiTx5d0l+8yMzyynLDJS72IEJtRAOSdJO4p
0q4IhCO7+y/WcIqMIdAGB8+fAehs32/mB1TGYlibQqLqGmpLjMm2MmfgxIetX8j42JRPn65I/asF
WTYtGAQ+4nQUQRR6eCuTMzUYOtbWNixRvKWJneTs/M/6Rsim1XTlebmFw45GiGS3ecRvXmEIwazM
AeXkaj9nz27CU8XjeexFP6UeRXnXpj24yjQpCGDYarE+6guGSWCZzPH/AGys0+DzTbfKuTQ5kfqo
/eZP8/E7Jyrgl9Ea/8sSPvi8YCdSMVDdmIgwKvMMKJLGQLBbCEz8qjtq3Imf9Tx84D8ovjCAUUd+
UA/y14AV49RODFXYLfmwMVB4fSAaosHBgHN8z2OI8UNihtblaguakLD+H/RWeOdma60GmJU54ZK0
nrCJO+9ZD/MpcJ4PZMPk9eCch5k60xYjXylVHNYFwYg2N5PUJtXjSx7q09NrWA7u9QPjvn5eim9s
+XgOWYKEuj/11SaG87PYe0RUBy6LTBTusmcqAqHGdRXN+pDvY6gd3fHDeNZdN5ZYiUY+TQRueGpm
365Z1/dq3TBQ3yYKPCpw5mGCBtTtWhF+Q0qur9Sd5V3s48YSFqVMpoey4X1ghKOJbgfk53UEPuOL
/p6ed9dhJNQdGAWSucvLnIB6WAaEa0akjpGCRMKUXI7JBCymjXKkRY5HRU6JMNf3m507N8ig4KHb
JFbCn/e7jEKLe1dxtltvtZzhNpH0K5/iU9rSdpNbPHkicCiAfizvND5xkItE+ypHFpjKDoz7BYKK
uYDf6i2WQA46PfvngPWcn/5CTheSETULWbZLa9+dtB+dT6r8mEtEVRX/OizxX85MO6v06nTk7KVB
H7pswVoxY+Z3WyjmpqhnYiZuf8bA8GHdTNaUAiK4B7MeFZBnt9oU8lBErPBzr8VsnSNbLVbO22vP
JZQALMDUuEle1VGRuVTOVjunpO6kOOKmCIYnSmqnIwUtvJgyIn82+SM/dGqcveS22YfaTY21Ag0M
ZfgbUu3W1vK1g/mbroveQZlYpe91SULknOV8Jj8/vEuF1rpa3p89shfoQV+CXO78MTs5KPKD/oOr
fuogvvYoFr5/n1Og4dPJl6XJM1ytsp26agRH3uku5MhO60GJvcT8hut+NP+9jzvez3zDbTUVQBA2
vGRH5lMxbwhJRk6kKXWPcK6u51JFV0nvjYOwz8aBmBf135gWFbDbGo08Lw051GJ3wqGjRCn0RcgS
+0A8ZN6awrthM05twnqjc+QBuqv7moHnZkQSbl2fM95MdYBPDLPHUVbhtcOrIoCMfPWkqpE9Sgld
bPfMdvetSR3s+U/+2cZFJW0xFAqu76CXihEzfE1b0t12iosJs59uyvt1z+6WzKUCOw05nDmk5LHq
6ZoZnH3n/jq/izAVXnkuD5R16t3VVMzJJAaDfzG66hlprqfQHc0FkzIE1rybAA4yLVCqzl9QVeZT
QQ6IDsW9aoKWnRYAvcnmuh9xtM8GOg2aejZ4nVXOZlNTQEcchcAhQEK5qfU0W/acfb8nLivMpEMs
SiJx+c9dzthLHEI5+3ijx1DpScxTM/EtW8KzCrd3VXU9TEcU+cnb3r/8xZC3hsuKiYmbW0/il8T6
rUzB1LkfSvjhU10bLGL7+tHjjZmtpjkZ9+njriTnOSVJWBAEFWnciScvRXOxCIfUGU2iFMekdBPE
7KJJjMukfoLJAIuXVpcagCFpzNCNYIkx+QepNNbIjChXcQbGv3MfUvFuEkxHhYA8yPyDASjbEzPi
D7wcZD8uLuvXvpmRqADTNLpevB9uaiW2i2GLHEQ28GbBIsnuMs9bwonsU5rWaE9yZidCgxed/juQ
bHhEn9YXPEFuj65aERIha+T2Ic/ZRSdHuxmDLLPf75W78/syB+JQGEKxebnAvR3kGk+Mg+HG4inu
cnwmCWeMxbRU0a+40YeB8jYVQ/QjvuOAyKClFUk+QeVPWmW028s8ZF402QYcvO54jSbxXeSIRw+v
44jtnYpy1VCUs0ssY+83r1vptebVdtlA4iZNZ9VIsHEwZ267uHYURdmVAvnMV0CpSf/QQ+MLoHFe
NpFShgelL/umGu4/nvbqAkM1mLcrfgfgAnALxgf7raXlkZInnZqcfDC4fPAnCM3BeVRyS5YYI1Q4
WnOg8pZoQ9GTq7HvCimPlTjVP6ZhTP09m1n1Ok/vOSrxW/t5lfG/7CQ+o83/QT+61Cgl0lSpzU+u
zYnjwC3YG6R2oaPDjPVggE80BGFi0JUP9asVtE1+fmv+k942b3jB5gorc3zn/fq+gbLuB5yOu6ya
00eOHH2DcdIma6d7agyUespI3yr8JnfjM8nYvTRLxkL3EI+11FP5A37lO0h78Fgo+Y7b3PAvOcmm
ApGesuOZFjWFgtY4Ti50KuqLdBJxwI+/p81nO0YuVIgVSV6OHGyBVsauzWWtWptT7HANfi7darmu
It3iCzgEcJ3cGq6HG8QUZ+UqOxPIhvllY2mviHQkeH1kQCzs5qqvWsObnLrnHTamIRecCajGBXvl
uMHdHvjlTnBCiHZK/19G2+glabLg+vxYptq9Jn10g82hXB0eYGmQ82cLZ68l/cp5BHr6lnpdkhhj
xUQTfzmGkpF5tRgOnPbVfST5Jm7Irc+M0PeAiRH5jU2jlYbmKDVR7NJ13jhy7yHxx4TsTJK9lL4e
GvPn5Q5C/9m6kIMFOz+89A+WjyB2UJfqZbbK6X/daDYeFdJbSHkVyvrY9S2Tr+5sOPJ+3Y0YsaEX
LS17WShitQGaJDN3yCLCmPtfPPz03dx2MsKW7p0jvIFMkWTopsrHhhuKovF+uj8DS2Ms6ixGxwjs
lrJGUIhTtwni+abCnZ+muYXgs/WV27J/ONlvgXIeXMOuWX6w9J3Y+oDy9QaCgFGSJ7PxnM8q4IIW
j24SgZSOAnvqWzAkkJ4QAjt40KmaipkYUB4pVVUDu7+uwHmtulQD4+SuVyaaCufUE+L5tozbwPkK
ABH4xQf299R4mNA8VV0I0JQ1PK0PkenUzYoMpdMpY/adoRnaghbBuA0U6VB06MKm6zr9VCy0T44C
5yr0XIwySF05ltxjI5HitMExRJChrCKIirYliO8HWTthtu/BNYkeadAKGr3O3lZcPPxob9H7dX1Q
BFk/KFrRgvQQQ/9ZN0Wc/5Jfd7S5FrN6t/IfC3sImPUaC0Sb3adN2JSxjORJQlCPnlMPcbRreyed
EZLvMv2CFg1luwSww1YMlIE/9jDb9Iv5lU7vM6/zYgWEWCtihQbC3FeduPbaJi/17ksUQE1bGFVe
U+Bsn7nKcCEY5D8SRYJmXAOXqCuCdd804JnpSemxe7OWDC+qIxsl62WujJfz5TIIDonwnmrKSAn5
9Qttrs3vHKBDOBAJodGm0Mfqa/eIajzudYXLpbFr9OTYA6lSkZVjzxjBy1Eme5XdK9AmLM1scAVE
Q/JRgjJ9iGV7FOKNNf8gQ7bOnu37O5sgwFhQzkJV+TZR3Y4NS2dGYlbVorE0fRIiareg3CoRgUG3
NYUyDvOn5plaO08pgDfLss7uxBsIPzOlj2IHNvrzYJUrTsEBgQqwW3YsyGtDztRIk1NSlF/dvs5b
Za+rDMR87687G+9BY1Ae0M4ZsWsveS+DFPX6r/DnRCpkvEwd+wCv0bXg1hNgfiTirN8+1fOsRMlu
kV9OsaMajAYUtb5Gv689d81La/B2gl9XJgG7e+U6y0nrdLAp+M8CnOfMGu23a2BWLKnnyEtPL+Mg
et7Ya6uJM4uLWqztaSBMULRpKkBqlpofI5uVToP5iB0EU8gcltw/93Kgg1IuOwOKLjEnZMssIAN6
UR1lvwiPjq3rg0A7YfgAbaPpgmbtXIPBZurvMubYyfaOGdSnz587jXMI37SJDzeozP7dYmFnLxn6
AN6/DdqG3JMD3EP/+azg4HY2zdmR1K46Wlg4U/j33p5S1Z+cNQuoWeo/OYm/dyd4Io5D7PVfS+o7
hRdshg8ze2hzqAi7pWU+5DcESQ6ITpAcclKrRgNgyzpVZISg3f4RLErIqR/bPQyF+MSpnOWVK/XC
+QRmw+2kInIUqOBW2v6xZ76qrEeVJ7rZDJLwNc45EZjRJSEt28+Y9/96ZCIp1OhikUsU6S8rhdeM
jj7sjfGrA1HE6pNzcpEKE7X/MBMUnZT/wJVRsMTcsR9/7cjojWyrbgnZJSNHBnaL9wUYYQZnb+su
yincIA3JK95MNc78ic4U+wpVD36+eLwc+fWOOrW8DzZsnkzRdsGyHopx/oLljS/UJY/tFmUd8pUK
nhjjQ3UH4Gm2HlWsW+UNUZ9lBwQlh1+HtQwM505ZBreRmK8QWvfh9izRJl/XY61u7yITWRom+kKe
jaBZSHBUIu27MkWd3Xk7M9b9D9hyKUH5U4c3yyoHVyM+9m+gwIlm70pZo8AsTEPGq6BhKJrUejmw
axEiv72HLO97IQmajk+InBAo4OZoavVJEx1KZMrx/o0wJdWJf3HAm2QCuLps+RQYnidTn6UEq3Sa
rOcR6wT/yRRIn7VVf3qTuvY9YeyHc6kzReQ8P23dS3XoitAvZIh+K4/SEXupBj4bgbFjxoiGq63M
oYmxNVrSK9qtUslDJ1VNN0cbtMfUmp/od85I5+lwYO4564s5+nO6isGzJJ31VQwfJ9Gz5b3839RO
9pzLiROGFGNva5msBgkcT5s2BfAmHJWp0aabXj4Jgj2+SUZVq2RASNVVA2ZmOZaCgD/xUlcEPJm/
wtqgSvK4v0H1eNbdgfnJ9AiOPCrhX5E/E9WVN0JuGRM+jPkr+sQzcLMokJDHDXQRdCne/VgUOwKJ
tHrCnVANBxk/wOn5lUF7V985yBM1FVsimUrVk4/V1heuoECtkxHK0w1r8iFJVzrUD4nu8rFLClhV
jszEEGF23meAVLZlyp4uOogMpNA3oVLrFcKaHulLDrg61rENhkiATjf1VYugl+ulV/TCv06mI50b
C+2hZONg2bWXdpU2iUlq1lnQA5E1FwuVMgqVTSJ2M7P6v+khqC03AfsUru8KnZX5ubvnaIBY34L+
8DqeCtW3Batx2RhWUUIR/ykrXWhAQL49DzP3k1Gtt6F08sc/tBFPxGq0V673E7q7kWaML6dVj+JV
KFjThHHSF3EAnF8j/hDdjuQmxrAiMW56C3uD2iNQ/gtY9J7Dt64mosMD+BMbRL0G2YBfypAFJhpA
9IUnHnGG6SqqtLdJxQd9mr5IDf3D0H9NO5qfviQBk5y7EdI4qm99ay50mLn5GtQv6w54Py+jMz0m
y+UgaekTryxKME4jIPPEAdJtGEM2yMAzGm8W5ilCoiZkD6j+WPuw0AzV8eMJIo34fS5r/ysPKH1D
OCMBiqVLCywfK3TlaI58DOCg1C/RMHjcv9ddVDW5Wa7IWCVj3TgWncq5F+U8GZPOnEibQWaQOHJq
NQLmhSFtG0cVxq030+U3pS26dR7Wyz3OEsTogd73u28KjmWx8R1JOeljky8eihMHUOakMxkYZGvD
5Sra1o/Ya+d89+eyZCZaaI27r+enCnRtLP1xiV9n46lRbU5nUaiVjMHZ8Kojwn3G1jbmR3m5Ml5I
swbdXYRtVHF3wK+GUgzweorDyx6SLz4VOcYhoFu1OXHugYfYwcJJnvNTDRuduvsfTqkpkoIjGSXn
A11IwSQubRIA3vUJJLe0pmQHs1+NbuMRg/yVmS+HY9xZ1OSx8fQPMJZsXiMVe4iy+L527xCPYdC9
w8tWxq000oPi/ydtSuqz+HqIM9w2DgFIw+Ij8LQ5nndv5aOlLTMAnmB8JHIlq8Kk54SGQ8KLmr/W
J0j5X5kPydX2CrU05DEcatuqC5PsZcXiHGsnHpXIFpI9VT0HG4TOkvTS3h2LpikH803G74SyvLve
Vp0V4V8SRFzPfU+CzaLl93aLKHtCp4R0mBF1l5Xmz7dqBtXyDh1V4vEP8LcZm6y3/z10OmKeNl5Z
zVacqrX30EC8M7Hel3oDHHW3dJ0hY0NtwsdicFGYK3eIdkeM9MTDghdjiHtVnmfIoy6QvPT9sYNx
uqjNQ67h1a0Tg1HrYRyoLoj5oTRj4WVtyGlgpEuu8mQI3RpVlz+I0rEL0OZsaa9fnkgLS6ZFAP1/
tgPn7ISByDnjW1n85dGG0SXOblwsA4oAvFSnDCLvkap94FKZ4lTrRZC8fjNObQHm04sFVlefBQx0
x3NGE8jem09HZgs9/K+jCVJVkgc+MENDVn0TnZKcvtfBKo4gMJWV1+QkvlV2Jadw+Opsp5IEyNKT
NZmWBJ4NoOPyv0sY2wyl/ug+LxujVHmJpM6hX2D26gyVqwpgN+Ex8EYf8gfYveLsgv0ZQjOk9Ud+
Mip93RUaf7k2Kmk/SRdL9xCUj/ugGshUy+iJJHuUfw71BqbO/55CEOpLH68kQdQn/BcjdN4QwApr
Cj83TtAnQZU1bduAEF/uql/9ju+M+obYzHoX+P5Koe+hf49KyqrXczaXPHaJlgcDb71YrQE6vm2a
19fARchbPAGGVYtpNAppBSsY/NavBFmg7l4ldvLfcZ0dIzyJVK5oCQEW6ALugLHDbGFHf1XdeF8g
5R4WNgK2pi7OA6tX5WZmw+20Vab11VYrF67r/fYwPGPn5ooYtVxUHePScsJiVOhUzSzHkGcCLuY3
JXMOy81RTQt/KIV4ep0rJbwJ7z1gkxEIIYsTncqorErW4eymPTvJXg1+7RsLi1ouLaw3UJqG7jk/
gLLwGoTH2ej3eyXiffUHw2U+nm7fbY2afY7BL+UROXBlUPqlatA44JMly5pn7OGzt9CO38aT8z5L
4JarV3momK7cGLb5x6rAzJ3RDR9li1TjnotncunmPvKEXElB9yOoBPOxAWHMNkbqK+h5Gn9wAypZ
T3IX+t/PtKwesJKyM1ZMzyX7Lzcby/2rYLdOV+hGz+ASCnw4kC44L82v0nzi1/f1NO/sxYcH3p0m
SqUpvbk7fShwlbL1GbtQ2IhyvZBmWiyipmHftJiOrhtRyJr2zuiA8qlqjTKaqO52Pjek7xd9kjhB
Wevd8u9lOYcePDOcRQI8tlOHVLJ4tajoXQaig7gaBPgRqL+B1THBQLE/kgL6HgWO3uHCob19mM1d
KIPo3m2gaGSM5Pkd/r2qSF+eWLLWDJDau0+8Bobqvou3RilY98+n0f/ueDm0I/uh2peX3X2Gb4L1
AnY21fgKGW3pZHRwXAKwgfbJhLdA/6dls4LDZ8Z7wuErh8lT09BmCfXRR7/MRBxDIF30CARK6p8r
xc4xYarUaO2p/pwk7vssKAkSDNcrVKhNUOX45/qCtKABMtFoxbEGojSvNUu3OFtz3HT2pje24JY5
BkvQuGuk8Xbu+zK7rvxNLmm2oKUHM1MqG1KrMrXXNxydDX2JcK8uQtG7qLcRLfxxiQLvlHK+f5NI
mC6blW2ny9xi+AGPWMi7SPNHBMIoKI5IlRkoBmI+vfdAMOw/90tAsa2Glo4LOchsABi6h6LHDEe/
V0BPo7mcvp+s2gtCH9MVOxrGm8Qxio5iXTn+vg5E2nnQcZli4ZYp7ZLfaaaBlc9Qyleu4xv0Sh0i
nf3q8R69Aoap1GNDgZ+AvUAMhc7TkmQ0M60TJmQs59HACvq5wuO9ZQdB46wUbeUhz9ui2LaB4n2C
u4OekouAGCr7wYoHEeSTbFAG2j5rHefFakYaUBOF/jCJw2iWt54sryLNBUpFwFn6UAs9EFOHtDXy
R6vH2fKhGls4ooCPzRnNxUCO6xwdg4iUsOQNErvWP3ThkffXYpObWa8XABfG8Wayx5zPt+dd/3HF
IAAyKWEJkSYlt3hr3JIkXBj61K5HoJUoYArlio64SQwGZIT7m9kEGOkohrznjVGhap588Yzr+ASl
+PGTlIifLzwbNIf5mC+JyXJtJua6wqB2W9yRsOgwOtaHtIiixc/fILr01Cx7aL97MPjWEr/XNYFA
kXiCl2DJwTQgZw/FCcdI200eQJRxsdZu/l50qK+rYcD2xCWLTIkL8xRJKPCdAgQrRH4hmvJ9LVrS
mdtKyBMQsycOyU+mf9KcjrlmQmwlnrneMKTV+OX9Ca0FojNBEJYk8q25UBrOy7Zl+gyl/yrqHEER
gSN4JV6fz4YzcNM7U+s8Pp20xAiw7JYu4ZX1/ypSDty4W6y/be/ubTH6JFR5UKXH89u8ReI3mrBG
RJssOpLAmBqDxThi7rID1zS2SI5pL5hofGfIUzpJ/TJFLHfj4jNj2eXxRkZ3LvoZq7WboU7FTzaQ
RUNi/i6Ay77BCMQ96S4swS5FuDDLah33wyGEGOKlQlIeyRX+UTqrAWV6ZyVhUg2CVtKwZkPpXKTc
VdEuZ09kkt4uTzDNqViHNzCAh+H/vCWXAQQ1UCFZjYIS6kLlJoVcRqH93CbsEB0YZ/EGvhU+tI3X
SED05EtXpL5No8AnrAYh5uLLkPy5LRzGLseMNS29OKw4xqbhVdsuJofAiK65Ajwj+u53RLPxLgG0
RmiNPTuA2JWCiOThC/Imh4RGMDaYTON4mstmtrdhHRJUmTWkE6wTpQrr1GA+7ih40FlictOxZf6l
iPfSxEXWYJ8YND9ZpBRPNU+aVGgijsrafaTNBagvrzEyCxLO2vKt99hZ0tNo1rqjBb0/U5AuWCtg
v5ycLBECptGhGDeYgFy1IZzkQseIG87fok7oSH0THsU7CDp7vcebICrn9CKpz6yOSVAawyd3vsBz
NELjj914p8G/BQEgod1DyuSL7sBMFh13WVP+3zIwRI2dwc3FE2wYQnWP4Jz+5dlttnLt06+ecFYg
PDyprh1Pc9ICm7jGTES5yHCzi16+6A4TpGwnP9QyiQ2JiJJyJcAJpvhVjSgDIIK8efFTw7XJlc1G
5OI720P4TR+yxLWBC3lGyzRLH4RvjzlHGAfseDn08F5U5kCo2SI6yx7HIyiatjeEc9MqRY/wEyak
13/mLZL2UhR36Amr9OYj7RS8jNb+z463S88xygz8ZGg1kbfnS0Y5uUgRECxJ6ayGx+TwpasWw1Ks
w4RvDIksEy8fjyvO6+cOLmkHpZfGxlzvqLFbqY0NAILTW1NnRjCc+Qd71jmQ2vo0OiAlfzb+Po19
dSkpz7ybYnrXnrTmfzu35c77xdk2zJ7xLEtPOq2FH4laInvtkQ+mrGj1MsIZ1XUZwLEUeNKFcjoC
hry5YgHQJRStjdcMiShz45ovz67NKnhKkiGc1ysJUQ1oD/sEQq9Rz64LBSF0mHeZO2BL/sac6blb
MvsH/F20bwelfcH7TqtI06ELU0zWWgmWvhetUHwlBk6Ep6qi4ODJqlqzbLG42loWjQPVkEZ2x5uJ
s5h0C3a3+JSD1vxGd8CU4KE1ncqxx2yQ36JLEsTenQo1yDRW0oz8rqFMKTGDUeISfDUkqYI+CDyh
RFzos62ph1t50jjCTzfKGRyH67RZbqzjc7MSvqJaOcC0kNGsS2QduCalBaPHJg7NVwVHeHJ/Tj5a
nEVtGUnFdF/UhDuvYsEVnm/GNnQPZWtp9AFklFm7yL9xG2s0mYFzCdUUKG/ootXWevB/DXwHmPiA
BJEXv/iCf0Fz4Bv2rU4YjM+UB2ftD1bQPAsYX/4CWsluS0LgWa80eo1bLhWoObvYI/tFQgh7pAQ0
JkUit9IMiTu/8O3ErPTMpJmRoXC5jzyDV9P/cnhYVOe63O3Nrz+FH0FW5EoiVhvojzwn6cc8wJFn
dsz1EEpl+OpoFox4aXg7wOm5S0Rokw+GwV4Nl8toowEqt+Irlq4NFlfy3Zu6x9NfKqSHzxxUlRS1
39TRNLhMKu1X+C8UBxB8TjlBOYSpqPyiuFlxFZ6Sxog5rfEU15UFZGsLgo/Ax7ET8FswTmMP5xUA
T8UAvpGOoeM+kcO/a93ukpdloiHrRTMPN2nYDcGhcXKJ1soanezPqdP1BS2smlBq5U2EmA8czgZN
/9JW8H0/Xx8vPBFeLBScJ94G6OqsvGFaZd2VNCXWWfI1xhEfQ4pMcNh8OkgZDwbYLFccSUS0d2nn
ZXK6ry00kkqTr1izlJ/Vw3xg8UoBESWFXbUuK60i3/fop0sPYwr9wuiHGHK5PcKgyeG7Sl7dfjzj
b9o+McZ/dj1r7Gi3TtHHjvqv3Ls38vkWmnkVAQ2hbwEJ5WrajNOelt4OFI2hD3XZMemO/J7HTvW2
AFnaScExxDMUQKuz/kSD7aVDOl+YZM+vKzJjziof9WUKcBHV6k60a5xi/upIGoZRz9ybZEwWAp30
/WO/EgtOtRQ76vRChjgjkX5HNgdL+ZAKpw1TAh8BNzkQWHTYIAGfUuUI40th0zoTMi3jMAuSUWTV
+TvGEYU+EnSif6AJyxbOapG4jvt62BuX2HI1euwDR0nurZH47F1S0IpC14W4bXmDQ4Ox8grf3nPC
L28mrJFAYCMiAx12sEYPSg3Byt7jghpIxCQXR652VjlIUerLqg0C7Ww12LdeAdF0UuUshzciTmbi
oBvfkb1M7ADMBmdgWYW0RGtxoqXFm1ExaoiXunKoj5mxsyzB4q07ngZQfV8Lsk1bbqhl4ue/2dtx
TLQmT3/LgJlLFsJ1Wo+GZ5LvGWNXvcxj60X8R6MHswGNUUqjVbjLSYyMq6L/CaeRS5tA+p9Lraw7
AeaxNi0gsvZNj6pgaMSf7EUzf1Mxup9J/zUxsSrELMd8todksrVTHIdS1NPwJfnnlbJyA9TF7Rhs
mItWyNlT7YdcqYYu5JHR+Zu69BV8lp5BUyyO1E9Wk27aRMfoU7nYPGGOJ7PRcQuje84DLmR62eQT
T1vyn4gXb0tttynz6IWNZy5+morU3z1Yblbuvi0ErDxYUjPCSw2UdLz+nZoDhb3sXHC9VTWA9OQN
vVbn6I5jwpPdBfLPbJdTE3Ddbop/LcAu4U5IbrTfiomDaOSTq/1/4e7c5ndEYUPLvl8B0CpkMjkz
YD0VsBTa3Py1+MD7Tn87XulW/DuKa8SJ3fQ9RKqKVFWkq6HPI40FNjt1bl9kHU0NA1vgWn4/4VVH
UpjtVDgg/wgV4P3e9CMDpIJE94mAtiwZUbUgfuqhza5IUf0bViW3KLurN2q7yeakyjBfEUO1lVDz
oWoaiQvm1walV9SwXQGFm/NccIw/nd8ukXAtO5WTZWD+lToa8IW8BhUpSnvcxvEnHy6vKSWJWDUQ
a7ytG3bOguMPbp+SGY1PFK5Xbk9wyYabWPsqn8sMS8+35ZCgPsH0nXdkyo3jEWSGbk92pPHfFso6
ZW6GQ5ox0RczqOdIecj6iRfTzHISz8iV0soc8LugkHQT75yoeVSydfC5jrk/2TDJRpqvuvY9UnCj
PED1QEVxi4DmmQ9HMSiWU3Da96BCjmYkXvcWc/F2/AzF4gErhHr4X6YEUsDdgNge3oZwm7D+fFvL
klxgsNQP37HK1QL+R9ag2DNNLGd3vQ49gIsnOt+oQf0gPkIZjPzUj8ypAq6d+/do/KM5xfInYyZh
yu67dcDi8KLnD9U3+IIpOXRyayu6e0nqqMiDEDhDgIds35rEYB3ypr2J1DcPuWWDnIYAyI8rMHxr
LndRxsKptRqbXZExDgUNN48sve69W/GtZchigQUqS+RRDbNreayJAFFqm7Ha0VWclVyFjof54CEn
03xDcOia3Hp5rde4+NVidDoT55TJ5Qrb2T+NdT+2lDGTt9ONdniwlXEtA0f87ppnd9iR65yR7YlO
rNEoi7UADfb/4l6ZFc3j+a41RuHQS+S0O+JXNIvxU/vtFTTVaHi9owU0eBaSWcjEgdrytJJg9ZEn
m9LlwdYvhvHtYivmlDM2xBh15vXhLfppfOFfdSI3NyT7jIknrW+za+XsDX6vz/SIwHI7ACIu+yGo
Uy5RGWGEeTBnjBebUBGbEp5uDI1p1Vd4ZHTXzK3dyrHzZh0TnNM636bE1m2t96DJIS+l8rDRVhKe
7FJOB3GZ7OGgY2ZzcYZl/yqkwx4Y4DbAF3veBnRYyji5BYTVPvpqqVPem+SEpGQ7FDMwleskGWjE
XFasPnspBEPES9c88ObidhFw0idigh2N/jlbohAWu494y+WEmjto0cZwvnIJkTs4ZmKES7VcZFke
gVSo0pYsKY+8T0T/UUNgeoAEsfihU+ziqyOqKv+Qq7EKauAO/DbDCJk8J17OMQ+piJMfCCL0Mhvl
chSbj326ODejNHMtaY30FzPIR51DNu58y6g1wo/leRvFom7ceFdG1ZCCqMe3+IokBLO0GeQmB5ey
eMeih14yPJuz8sGJnDwhFrapTOy5B4R8KeK2kjjXj+SJhzj9ECz2O/8IGvgLFksNW74Huv/PL9D5
r/TTVn2vfQ76YWmyn5R1uAEJqOHcvsLpUasg+EsVoSM/Fv/QWknrl1+DIfEoIA2siCVKOLdHQJdh
Hdw2dcmT6Dw0A5TrsOOIot8yaNMxGtojGig1Q8DqwKi6SG8BrUK9EbYmCeIrm8Kjj8piDjope/VZ
P/drtxVIUmZ1OA9C351FX8DFdLD9Lq65IefdV20VKFlKqDSotfvhtY2CH/s+QRWq20OW/ffQN3jT
5dwdD5uDMsRmV2bJIcDPFthipO7nXrED0AVqEd6FQNePpu8t8AlJYO+8rQ6hw5vkUFgz5KhihRIH
fRoq460z70J+g7DqCvERiJYScnjAa3LP2ccRJS+qND4KRJN3iimbrs9W4d9TC8auPCnkWSatbn5a
jqEGS7nIh0ZXs35MxPfdzG+EXhyXocvRenp3MQvHSWI7ncNds/QyfYytRA15ZJR+Ok1gRbo/mxgA
qGiQHFpzlhaNhhCwv1rS3zelfcCy8PAAQAcTtkqh4AvkqwEFvtcR5GPiq6B6Mw8vzIl8juDrVJKw
VkaNjj6Y0LgfzJmiLOgeIovj7HfcK0c1dCrUZRaI/PuyGlUrWBeLUYqBdcgjQjoHL2XvchTPFP7R
89nzAkKTdiuw5NOZ+CHNJFZWdYZ/gB5IjRZmPnBNlMgR+Sgc9ycXaObXV4EEommxJSc9IvdmX1J1
zn9bmjSBTr6RulD9NDnOBF5jOzbKHkLfYZnTUb9XdaIrNr7rNJWzTeL2v5QNlH6fLdtQiqsmCKU4
8mtvELjPPVrqfa8ljUmGt3wqnkjPUV8zo4iEI54kZnXBUiFiZXQJ0iS7DNJBpj5tnDdL8YCCN4uu
V9F/lpdVeDzpoywdwUBj4/Q07AnaLHL2VoNOWN311C4eoQNMwmRVYLsKwt5YnsDrQ/4UKs9G/QDd
iWuexS14Pcx3h2Ad70nLuB6ZsGGRh5Ta/8tBW+zO5Ik33C/iD6bQvD4msivSIsts0G9mLPgnwRY5
5rcl8DA+PLWD8cmZKvJmckNc76hGNY/DtQDPmAeyqLJdggJ9MfntHOsYimTHBfnr/nMTjTjJwLGZ
Eg4sqRCtX5fELsZMYSz91wcNR1Qcx1nirzGO3NXw+hWZ/KY4Gq7sNEVRh11vaO5ivT5gQxQgvV53
CTOUtljzwPj+FM0EcPGEsyfEHeL2u7gDFYOxwN9CikvyE13q+nAIAWKsFUZzpbWb2wcT0GZp6Wph
bWSBx5Sfhx1lOysvIi7kPVp2Ne66icALEKmCz+kGdDuzVxSLl2EjU2cRuvkEPs4j5fiR7/7b8F3Y
Tq6hPMDlzBNeCV96SmzCYzb147ZuqSELxgn4rlTMv8F5oagJHu9a6lXen3b3OBZw/5xAxcowMiAM
jU1rR//EfPDze+HJe88Xidm7rFb3/N29fefQgHWieM/Vug8glBJQXgvz0Se0Pq2sOEkGhp3eLO3f
E7BhRN9KL8eHWf6DEg/OhF0Se7fYArKe3HJ7P5H0FXLr864wdeqN9mJOrsHvDL0E/2hfP/Om7wQj
LjnOXGtueLExzpDJNU8gNqiXDLwV43jQp5IN9VPj4IIrMYUmj/PIi/GQM7OP85XnyqegrFbqqwgS
7VV9+imd7wO6n58wPejak5fUiYZlhDG3KFNVyWCLkEYAh5aXMgk4bjydRfP+c88SAWum+hJDAObz
YxpU+vvtSNml/oAXnkXqvDvCaPizzjLLJ9Zh3+eZ+hJZ5c9Mhmoum9yW5PI4BOX3W3r3EC0fkYwi
HgL9ZGRjr+uni3sIIiq4RmFRRIOMfnGMsD6SQhLV4qqw2Y65Arh6busBr1ZZGJhOSR0krAzWWpn8
dgzFGuSDq9HJ5MyFnQ3iIhyEc3ySws3OLYPMTG24s+46aOCTBKaJ6uEdRWn4ryJiufrfjffQ+57a
mz3acmZOdNYZILn4EFAVukBRn5Fi1toAYdQ5hXA404GAVg9GXsisppcvWInPqd6HaZQLyA59oEQf
QKKvwmOwRuKKdbWS+jNgPVb68OfH0otZhz4odglNQ7+1NxurK0NYg16RGx+x16iM6prJLO+OyplH
s1xgOUi4AYB4e5WvoB4l59Qyoy1Jhk2y+KEulWlpI+QFMfJTV2pRYu9sSIvazRT8yAN29KntACo/
FuYaNIzIKmQQfnnJwyFP5htgPtld4OpKtX79z2NktzQNGCCDxweWo+rSWxF2H/daIZy+9oR4vGLN
WAtmSopzCO4ux3uMucMdktKldtBHKkNaTyMnqmXNCIEGD2XkHemJUYlMJiXyeZHpMa3VnkLNfdbe
KSYXuBpgeE7/ebmqndBeCCINULIR7VtMuPlblY4OKR/Z5W9MSp5eWVARMKsivmG7KoPGu7+WQXBN
JiTZ4QGtk2kJ/vU84UjhuhbsR4GEmAgosCx3CtrbOdJKV5AER2UbeN2KDbrQnIRzLnZbkKTwEfC/
xc6f8mvTeRzgkN1WWIuElF+Jrq6pi9QgPzA9G750CVvMfQObmnHoIcUZzlN9gFWiXX40FiD+i3L9
9YGs/wVgPY5xtzBDwuiH9rjpbSp2kr0sW/yIs/2OZ6gyc62NfM6y5invor+SWrFhzfx/RW7GhaZr
dRBltvIyWkaTqUQOMiJqpeCstqOeIJaf8gb9iTEOND3CNDz/d3lzccbHe8BoCYtd0aPupeXn7W7r
1WSXZwJ5wdPYHHUTzDc31huogElvHCyD4JF8jS5LsXR0sw0P3P0tNFPuIKtDc9106s4dtTkc9anF
0B+Ygsrck632DMnkdW2Q7xF+IBPZGFV5f9E/CevC34m+DFmAfmteXl6alttDRWFZ5FaloBSwPcso
iQ0JMYWTyDIWkCxobjVxdfS4jf6V/47HVRuKJkC5S0fgy+yQlbxMVgWsoYXgUs3RNLzp/8aTNAbm
bNEpafo62bRpz/O7meKxnfI5q8YmGKKgLOn6LAcgDV9TIpP9L08kmnr1CY/fINz31z5MaMm1dFVt
w2dJ46RAApAchZN+9G3sIep/qOHW7eCIu1eG0Wh/z2lWb/rP+WoxSFOdt/ZMPlYX3LGMGJ39bP4E
lAiqnbX/YKYCREGcbOpxrEzMDWzVs1Cx1VkqB0aHk/RyGd4rykxXWFPV0c1ZOaBMh0OeGv8KuzXC
bc5Gjof5pZtpc0ziFYXLKQLwV0nZlww60cs2yy87LINCQOVYWm2ZsY71/hE1yTDaKCBMsZH9fVse
3ze5BVqQ9ICCxMzYndzgWDsHCmczJ0FdhFFV5QVkG8jG5RO9VAkipKt1SAtBV96plLRhpt0nv7tS
a9xf56nbIoQhOlccrhY4UQJwSXUhbqYYExpaM6schsxlowCwmVFv0KOTRMdLpHs+3FsOZoYePna3
267ytM0j7Wp1nkPl/JoStuuPUIa1qP/DOier8G6YJDyel5S7cpKb8Tx6lgrtju1gvnC8l26Wsz1x
GoF9mpDT/9WsaX6T07XI+Is2toyEQpfBnGw+xUK2NhMwdffLXle/xJJykscuJ48oNEThqRtPGMZ2
3LuuS+v6zi/jROX09fFQxsHFq309RRpS5faIZEiehcBeK3ezB17+j3/hv4M1qK4auel6sG/aLYSE
1QNUlbAfmMUKI5HFHrlWxA7TEw2/8nUpZmXeFPcrxY7sCZLss/xGrMVVyFwpXj2umL3yNhgok7Kp
s3OtmqP24HT35K9UWa4Q7ZsHAB0f2/CDRCqPSJSFOmldaSDY4AEv6ihy1bqe/m96UfNOg/Phgf+O
NpzoruooRajUfPN03opqtPo6nhjItW5uP9VZLxI1m2gfFgj8YFNiT1cJoxj0H+nUCij6+/yCdurr
tid6MmnpBiv3F9/8Sjeh1Yu/GtNlIZUaXJ8vvs2SqJtiW6HlvKhKXOi+f3t2wkIxFT5BT1hIbnBZ
TNHkH/KZYi86L4Ot6YUzyrHzTUEkZ/D8LM8+Dtw1DXagcabZfK+vdBWZUeZXvaF8oIKfJvD0vQ/k
g0yZDbNqyxcoLFZiktHx9OkQoD8Nz/calK1Lw1W0p7+YTskdyqQmXFHKGicRXZDXKXi9PODGjxzF
Qq9RFrOaAufOqddYNIMDLL45nAsdJmPQnxK5WclO7wZW6R9rmmLjPUW6gOuQUitfJ7mrMLiAvgJo
KxMSpWDmt+x5Ei7axUVmZ7VZhTcvDRqFG7mr2iUe3x4QL98cyYNlezSYE9nzm1MQBy/wtpBNZZHZ
2dHHpRWCFvrQNBY6DBqDwy6yTQ/EctPRUeLrBYEdoQXMOPat4xlNIAoxl6ACfbDpoiyyMxLzDyFQ
yXsCzRZ20jUv+Z/vTZIm0baH3DGe1JbZvtj7+IPQJeN6yY4CWsG6TVZH7ooWQAA0ru6O1tIvpnuP
qGVSKrdFvNOg/t9BtlysT7la01ta41giBv5PLCEnmQtNK0gqSqdoMpQ/ijag7pme42g68RF83Yqo
DxmsZIW46wqlOgL0dhU8GiDoHHkDtUYCB1xVd+1vBsVePU+kbfWK9iWVESAisHcUb8TSdYO2Nvj+
79jGenSe0NvNt30ymmm6fuWzAM0hem+vrWB7M7Tou9fKaxMySCst07rdE+U9EN88T04J6YZFDwM+
6JFeCdDE7O80OMokHYrv5z1q6HyU7HzIczm+kQNNWDgXc2hAIVVAFZNJuLwWXvPoXd8RPrmRYhIQ
PTPdWzS5CyZ+RezBglZ4r95ih4p11RXbF3AON1boBGM0rnUnw8xXo5A/I+NV4/RVJpnlLCXhtKCu
mqWSTyFumfaBUNSKOnjB5VXnwzgOItOwX7Y5Ni1wbtrN8upW3kpaZlhY+nSe/T7iBilPMWB3U+E/
bwp9e9O1d5vCLJtPmMHJZfKG/snxDjqRsHPawt2N2VSHXN9ZOAkSsS/XvlJjDhLvu0RIJ2seSV2a
FNzouTaItXiOMLerFV9o8LDmS4sOrzoNmQcT7NlG+xGotsDPgzYY5aYhybSjMn9unxYCy4HBf445
T38k8hgxgj49uk8wTKL9WYxVwPaOob8ACjn4HuBkWUyV4EJSCEa6lht2zYOzHkt4Fbn6l7LfFdPI
pQw5CEOQu9+n5jYiW7+eBn8D6AnapptZ0eER67h/I2jfq5O7/GNF4ufNolk7yJYq/mczJhBwgOLa
NEHRbEe9DfDgGLoP8hKRtXuxzIuyr/w/134SzEOtb7g1lI4esooR8kSk+6SkeUIUAZp/c68ujYcD
pPuvei8UWgyMv22aBCGr//ZyEeLUMiT5k12K6EyFaEmbpVAKasljbfm/vuDU2ua1kJ0D5Uo81Bm4
q+80YpLsf4YwT18X2oQ1QxA3uzvt5rdPunSaYsB/e4DFBPGha6MoFfD5wZ3rkg2CLv1viXqbGuPC
9RdSbcRp8X5LnCEYGfHgHFWdEXrPqs+/dqrPpRISpdajh+dlhv34ckkD5BCLlpe935AEhs8IPqcb
fRmXOinV71gxNKYGghJR7DtmQHhqfjMI5jyf3XXGGqvb7mXrfsEgPkWZjuZcH/oYZxqZl9XYnRyY
UTiqZWeAEtbkP4IexLCDgadMcVWz6QcO/VEBjDtsmlocGe0zdg5YtElT7AoaDsr7FNillrOcGCQG
207Fut9I3F3qvKw76bJVj8bMCm6LFRjpX+PALDKTo9eZ3tW42GXGwIBq2ZcfCWju/HvDbNss9iY0
69e2Tl3IFb+VzpWCalKgrzI9o6ilhea7fiJ7F8+ptF+OGE7faP2GC4UAKuETVx5VZ07xlQ3ghqgE
+aXkY6HmaudX+gJZi/tGSxU5oXQhoHrdN2+3tel3R/andizs8OzdI5DOJynvkZxlzx9gSXygArCC
44Jx37wBDXrKomYTTLPRN28aMo1E2INy++LQc6ify/dZgFcPMJHaxKsZUVq2D2MVUoT+5a/ub029
a2c09cr2uq3XVQWTOa7oFnCLNmJRYWVlQ/mHuNp8jcb+NLMQwdsAmtx1hr5qgmPzH7A+ngbAPS6a
7uoXX8Vc90PjtBvIfX6ynIiwI03rS42Fy0UyKvZtFEeCEyk4xdHZhkf9LuVnD8PdosJdKBhgbrDQ
pUJf0529ESuy3HrFE1YTZ/dCPqCuyYM+AnAXhaZZgXZthpT1/RUZP5r0fIs02PMsng4VSYadye9r
4B3LPi4MGmdXlV6NNpAZWofOdYv7ywKuNADJmD+0p4HkHr0hbt+q/Ph0s+/XaMheTbDNbiCxAZZK
GnBk+Wam8TUB52IeSHdVmlD9x2gho5OSY9qX3zhGrMOONk7pHYOxkPOb9ulSM6dvQolAudLSLJyG
fW6TOWq3//KrE2zpx6HgCD/r0coTnTEu5tHTr4yTCmVy+htiNuxAN3Ti6lMzpBGS78mnKnxrqrqr
cZGR/Ur6tZ3g6wZssI4PZGxygl1TECVMh9UKp6UvH0kynFuMgYibvne9D3bQmus9XOREzdlswi9S
m37yUAWJrN3NvdAkWkkoTiI6BePMu7PW668Y9o44q/PqDRTBSpZGcvpNdBuVwdUbPocusmip5on9
+SRc3xYQGIbZp4V6W5GZuVulMj4YVkh8xg8YnMyiIGxApbCDIWI+ephML4JWks8uZ36us7kt1H/7
9MK1JkJTRCFJ/j23/VGpcE822zYUwmYwJF4xitC/sNoRaekXS5Ex76E75ySAjaSYe2YkDWe2CMOT
AH84i5gPREsygKI6vAF8lFsrIleU5WtvUcFWevshN61kAdAy+5370iLY5g5UmNGsu0nxBf2CNL6B
xttNIHfQ5ztfIzoFG91aeWOPcvUK9OQ2Ykr+XdvcLTAitnoIDXMF3RxpJtDNdXvilzwt4rbjPkRk
oH1ybneFcyNQ79pCawKECq40Co3/3dPnIh1GoB9TmCUV/TarThzS1a23q/D0rTa9aSsx+C9StIod
O+/kV9eEB1U20MpDUY6SwUhPkDrJYmu4f/XNx7pvDpvlUPnDJ5ttZa3NXLta305STRFFpGeD6ZfP
vMM+MkTsGLJo736OI43Cg/pTr4OSTgKT9TD/Gl9StBni1N6XEd3fFSw5BXwtLBAe/MCjch6wp7XY
PNj6PwFkjHB/k4UKuJcFSrLtWXO2nFG+n8varr3l0qKCALyB9OjDqWJ9GCBYG2Qbj8gOsscDL8ov
LojKlIDujQ2yP6FU7r1CNug0TtHdyiFGjjBu3Eaa/9b4dYWQ7YiJY4CegMb4Ad4UyCHRATcJwkI6
fRAOS9YWar6NTa23euIhRCNTGx2Vy2auU8wFNftZ/AQBmpFsXP/TfQTYzzSAPO969MkTBuDk0Pgo
Axlh4dlEGQbNjXyvqmCOyIoNuRsS8e51elgshnppQxfIpG5MDbX/mTQIor6g1vzfmySuBdY6o/Tm
/n8G2vdS3YRV8p0nIqW2vpgpstcUJHEiCzKPoeIAF5PL/qG4PRqoFtjW/fn3O1+rW6qQXif6D/Mu
hNJK+WjhVcs3ybpY4zKrq9I4TprRWwQCqvXJAP5ucrZSvVZuBGMFNj2IiD+PKtbJZQW4VAk5G5c/
LJ1dKonfQ0OAElkB+JKcwl11rrlEME93Xn/BpvWRPw11LsiBSjvd62gTvXv3kGRz1P57k/7F62lB
1mmp0mkWNGhlzG0zZl5bJ5Z6Bf8T2UZajOmdI+8HQ7SOBCYm9UTsKFsHKacujX769I5jWNuea4WF
VAgKoXNbTEqzb1Xf2+rO7wPAWUnsND9gxi7+9D4ED8nIXwbpidJYTdycOsYNNKjw7Htt6yZNuVVo
N3I3h5xcF3JhA8pCbBqOprxoBFFZWpKjkK7ZoyJBeEn3qDG60h9vhintiqwPojqWRW8rF6e274HS
zpx8qBK7rjPokX5Kri6BMjK0aQNoFBqud/DK8wUXkAmSlGEC36qbnwgVbmXHM6OHMkSI84Ej5DtV
XMpVX9+WzuSbvkDxl7koTqHLKMjQoWiQbFJ/WV55nWnH9osLlYzxFEv4i7CKLHlHIdbMbIzElpqN
6uSQm26oyyKE92LcObotJcKsWUBiHv8dJnZPW2d9k94VVnGfxttgoy/ki1O+Wd7pCc3wggq5ruB2
kMquUOgrZ82fDH3XrR0YnJ4NRcP0D7hYdwVsLkftqomo1Cpy8VpvLuqEJQNiW/gSU1FFiJt06RYP
qPAG0exw6/pjSUVDMg7QgkirSEEHDd0KRX8BtM3qpdjWyZdF0h9fc/w4p0OOJYHQCb5Nx1NkoOzl
PekOqVorpWAuOS66KI8iGEbGvXLEMO2eEl/NTqxTf8WbnM1X6vJsDsHlHCGmuUVUKwD987IHYGG1
YTZOqW6ZP/82x2Mx1Rzp//weZoA3HoJxT8/7p42aqDfep+TlggAMeoVRkkdV7MoaPcbpRwq62/yh
Y0B3nVvwPOYC17jsSqfelzt2qxCUdLQir7mj34O9XUnsC5XQQyRi2QjtVZU03gMtiwCw6bPfF3tq
dfUW3rNzPljB2UOOQ4mOvWHxNeEyHhx2WVz+nmHEIIcBF4h3N0Dfmc7Aiy1VBCfOmc9JRfEypyLA
+2H9e4IhfLemDxFfyYT6XMYMnu8GLWSmxt7xXa0RP+k8v4V64rEwScC6Js1n2ZKcgJHBKIe3LY1L
w+4MHq4GqW5CmXnMB/6Bn7CVJRayrVh0DJhhT3qN9rDsVJoCKeAwkGrotBt0dLuuPfC6UaCICRvN
vdhw3e7hyA9SPorxg8Mf6CI3PZXS96+ykzfEdD0lydIqjo+F5+7E5Qnanle7rT7BOKaPeXbVhZyx
4FhqOR8+XJ7DLq/uURJLpTECdFXZGJyDI0nwm44//astovCZfJ9VRW78NdzhQfu7C7AkqS9A+H/Z
xldYnmNZ4+C+uK+WhZhKuAIB1oXW/bTQ4gDKTzQEePvWR5SydMWJ0HoMiqy8Z9k1r1kOFHleASAj
z2LkH1jg9kw88fGGmVtWzEizMCmU/xkZgoyWjtnja7hwhJ93VVPMEGiTKuVAwvoc3EImKgMB/AUx
pJFFGejuNYG2uCoWCnFoozDYVou8B1Ib+lknyl4C52NjNyPuwz6VGkY+ZwqTh1ibOUsogb0GlsNH
pCGxmvFjM41OAiLNqgMvUk9N0MwLzU7gVD6U6TxjkRh9iWnaCp0srmb08XQ/YcBiNitPqrPhFBso
w7qxsYQV64n6Ku7mbRLLdkoOhNejSSphaqA7g1pwH9xh59Ebd3Pl4rrSuDOpUVCgLRT0LMHz67xa
2Vmw5lUPlY6rDbiHVcpeXnZgENsn4mwTgp3XNtj9L5ywnowVrldRvAuZrbxT3p/kjXaFIo8z9BX9
dAX23LGUZA0+cEl/5+C8/+/IELgMeWFe53z06osJjO4k3jsYzQEPTrTG2VXKU24MdsWI1NuihYiS
ubdFvKc+wbPHBlhdHQFepyz1uyvXVHd7XoWN7qEu2MhftyS4uy/jMuPdrDpNLYQgCSsag/R9uV8+
q2H+vDYGRIed3OdogeMbDCkwXc2gw877E8hJm6pTSWKJedPjZPwPSrRLOf0Zs+8Be1PyMlIJBshT
aH84VadyDblhIB6zRgkL78GQx8rg9a83Kek/4CrSc/ojYXTHeDoZglyPzBnnbuqZ5FWCcyF35+7W
0msC2vK7Uqd1sjPdRl15wmMoNZ3mDtBl5/D1VVYAqFZy4K4uNA+GnKX5mFpO2Rxbevfx1FSxdce5
ZW+LBAiBfbXOXnrSzQP5O7E1XgYJMWgKWMiOhsBDLxUkWF4+C2uyHd6RpZA3/YDii3P4Ig7MChFj
nEzRO7jzMdzJK826i/DkSjfR2AbUpC4NWitkO0i2pgDCW8hQpZ0mml1kTUh41jNgCQNjBnwiPsw7
BVK32tmZJh0Xk9wxujCe6QOmxWe7uNc3ADSRLblsT1LjdxxpCinLHc/iGSonk2CteRHx1rjxTXkm
Q1XEz0lP9saPmbgDMEc/lLqnKoV5uXtNYsCZr9S/gaGDWZ+aYoxSn2sNQjrjlqWcXDUCt7m7/ti0
tfCUEYFP0+XMGqv4bwdc1H7blKhLrNtJAspQnoA+fLAS945lAEqe2ATuiKunextPPHnH2/aGyApz
2A6SGqZvGvnhSasSKPszsSWEL8B3XRMqd6mJk4AuhOM17M5zjxrjy+dqdvTGW3Qulu8JTSJC6NrH
p+TeIu1cYqHVaWGXhXHtMoV8F59b/QbFPYBkoIFKUOOWGexAAWpaP738FPyxOYMI6xeaE65yZp72
mh3s6fNkDIAuJvpRWyej0f8axeTmuIw2g9UAnL3JLW6MSg0NFl81wMzAzeMDLKgEROW7LF8b2PA0
HydgWZbaESFrNxemi4ev+XD4rUuaNZiMeZhbbjUr1LjgCV3Sc3JGAMZQdFANp413ti4idcOict22
LA3It6PR3p35lPPUsg9g454BRnIdq9Ir3/k1T9/y3mZnqIGfpVPBYjw9ZnHamkX5g5m2dPtbE3+d
SGajOWK34wyf9ay2ROrbsMn196jXpK+nv43YUmtI2bDFfFahrnFZ5oeTRPDdmXrsXL76hN4CrCVF
7PHXtM6JrmnK3eYqd5LwYhDLuJl57iqb6suB3/y7h4qbOVEkLpVFkqeue3Qude01wkcIIcHHFK/E
HgdD1m3YOrAMOhwAVVlKXTb3ZvQ3T00vPGHv3Ugjfr+s5cMgPGrsfOHh27c3svFHvAywvVwP19yx
ohQfs+XB91XC4rWYrTeoiqOCAMy4//pHsoDk0fotc/rxpidYI0dtezi63nWlWZtf/N2hPg5u1dDJ
ra8H49oXOjwoIaZYstpW2ivMMX4/+EvV4+whwonFwhV5EZhAZjGcNMq/2E3+8B3pu4z/jH9Wh3KE
d/avQPVTFWavgNBlvwL29XpR4m+1KeR0llcAQ16exXZv3x2873avWd1eiilXfZRIVtnIsc8f6yGW
ASZM36TlHAtaAknsq5T7vrffWbHd8YTTiDLZ2K2C/FL9pPEq4+scUm6vsSQ6EBREUOUFrbrjhmGa
JUqH0DLUYIJPSJ0iUaGlPpAArOg2+DvOsT4n1itb5FUreHmwIwuGopReY5f/ktklNEWjn/X4dUJv
uu610WJaZhJzGUj8nXfyEFU2q2+lOtwRO2xntMMYCSPhD5wkgBEVdrguLKn7c9HsZwM4MAMKiuHb
gUltOI1yqdNB+Duxgpr0pyOGVMHLCThFmTwPIep+aMTTzfDei/V0uPWPsSZ+FgSGaEZYYDQiWW23
TWVDJ23QnzOrJbdATe23qdsXE9cYPyTCHhfgScMR/EYxAA3/r2zE2wlRkwq5B33T09fI7i7B00LR
wfn2hT67R8bguMie25nQCNZuBm6g7C+XynGtwKO1EBFXE46hbNiNg1PGjT2QEK3DG7Z773AF31Fa
ji5L5ExgtnL4zEaK8qXcvZqNUzvx8C5YCKX5ZwxCR4j9+qabpEuWlLUh9bcGmvjaWuQ5aA8wrbGa
pybSuQFkOaJsze2u2ZArUgZgQW4Z6uTdDxakcIVZrTY8XMjPdAnrYylnJA6hRLk0k59OXylGLjOH
3iwAWt3vAQLIXaKOnaogRJTFD8mtVpmYU7B+b/dUIiMmxZGG/0FMuypsKSg71VDlixipU8DL8m94
+n6kKMalNaomYqL+q0XlrmT8lEP4FObDTgNUAsXBlOuMO1MgFbU2uyfsTVGIf4EV2U/ski/t+zni
mt3KZPoKxYohdI+5mpzoKvDaHqnybHcneZeCOPMR4hEmnjCzwHYhILwDrTm3GRQnCQuSNxVATC0A
y63gtCTVTcPapH/0z6LbGtdv6npAxXnU+CGQX/+IS17kDcjNHxCUen8cED5tBMoAzJx7pcMIneaX
V2n8Uwo8mj4ql2yEy5Y4zxAza44lx17lSDBgfILZ8fGSip+1E5a6p85aRnmhHe4HU67gLVw15SL0
WLJWVlSIldImoNgNN2VFrak8dSOfjvjGCCXQ8qrE6nVu2RF02AqAaRWB8Di34She5yRw4rT/fucP
YYFGd6UZQRj49zMORbBAh+orFOay1OSMxGcNTdawYEksCtzXmK9ovfFsPuHUG1q5KM327dCRGBzg
OMKNo6E4b50LLuhgBBOj8aYScVP7SCVachU3E0WC63xJTcCXhyEUPQTRX8hQUNcUAIwAs+7fHLcI
tmWREEqPI03mfZSb4lVoPfM/rpkNb+j/fIfXWIA+s85PwpX3lVP36u+KrjKQZ2bWiHi8Ju+qj0UM
Jn3rHyCaalrdFneeTvu4Lwts1jpOa0ve9BTT5cSIVEmobgudh/vCoP/0kbFQkb5tZbqBwxVcrZlS
JxmVKzQxbqnsU5LiCZT7vNcLrm98yvhhv459GB+ejY5CYLN6TxtGH489qIJLr5LIL+mHnV101pYu
OyBJTOLR+9jg+OfFIT+QGaTDFKn1eqh5jbwJJuelvSp8x6fQVvn68BaM1ZQ3feoZrDNk3+GlxYIc
9Q2OJv/gDT1UlU8ye4JuLyjTVQFJEUknLNJTo2eJJ482JrlsSQyVqFm2NE2l+eg2G5HCm6PeUSVB
ntw69x7X/WITotIOoYviAKB7aO6qwYn545CIWBHN0Bm53goAcwiNnW0iT4/c0WiwJUeOjdCgk8qi
ykvz/Mh3OlsMFeaascAqJy7va4fADMrbP4bnI/2zV/MztxjGa5C2QBxUDJi1bY0AXV7KPkYLv2gQ
MpGxJSCn3h0z+Czg15+haN2eWixDRmrPZHHG4VosbJw92TbLfq/SCrAfFT0jKKZSgNRSXXIXwwuo
Pq9lO5QwYTVIxtLudEjiKeRw1SxhTRSWR49BKaZYsb0DtOhDlPUcHgkI7P0Z2cEZi0RkT2hfRKJL
JNMbHlLxMF7J0kANL/6RQuN+vFWHGsaL3mxZ8hLowx/n/Ce3Sk/sQtQ0MZIsjYnmRy8Oc6xFLR9z
EHZXA2FkaSPEvKUtrr1R6gKQYs7YDJGqc+ZblRHYAbrEwZTRTkDsh2JJUJlm9TfHYgfcarYTmrD3
M5HivYbNkR951ZWSncTsdGTei+YUr3WpSBpSRORhe/quUSQHxJLuEvwK8kfOHYwYBAvR1GbXZoha
o8UpeUxGGiR0N0WI7zfJCEffWy6Y10dH5wso8EOQz/O4suMgbCp+huIr3GdoYfcMaMaYjEFHTOOd
Szb4pHTJpfuaeCWPnVHPUzJNJlx1nEfgDgPsJGhaHZAh/SqT0dCMq/aH6dFQ07/HSHPt4tU9XUHv
qoge4haYa9t1L3zsS07+mzv0OtCkatJwNEO0Z8n0ut3xyEpppduZGAFLlpeHcR0L6Z8c6NPzPlHJ
WdwrIJCCVB8vNmVxuBMPj+I105lFc0eir/qMrahVY2K2018qmG60IOllQMgQXWSqUm4Um/jNhyfQ
/AQ7yT5HBkeOso1I8wReCWea4DS1PgJE5bvdCW1Mf6pfaX03z3HqcBaZ3r6vJ4eYApQd06nWI0jk
QEWRIatQL+NO67Svd3aH+Qa8Zh7RPQOSVy6qEYQEtDYRw+G4FqYycaWFGA+LXOowwrNPxmUfcRDt
Q0RepIb+wFRpUAH2RN4lGNOiu7mG1BFv2kY4QmkTMBH6G/RRMtSyUoQwp0LTPObNQBnNr5L1ZPpr
Q1U81PB60Da49X/RyT+ZtXJqn3wOW2L+jPbFCnVAcb5ZUn2m7WEgHQTjgXSL37okRt5oz9ovHGge
DmwAamkefcjQA25090I7xH4+CNBa1nvxlKDijVYpGI8RGjbmqwhDoF6k+bUgSDhuBcdj3ezepzM/
BHx47MOPkJkP/AbW9QEJIvDFsdP9lB7hzcomKmcKu5mJoVheMPf37XBAsfYfRGsKfxgYWAADw7M5
jlaSAHUa72+KjQsLEL2OjSza2+cB+SuJT9dvjYJOq/sUX7TGcoGqnsncyQx1Pb4Tre6W/uRwAtxO
V07tkZVnpILlIlpzH22pPZtzn+t3siC0QCZRiSdZ1ZEKT/8Wkk6BbGeqXssyrwa/GOELfcC+GK1y
Z5p2l7KlpWWCFXdInzEeV2CJ/+Rt2cppXTJ68I10iCPARPWjHUz8LDloV8JgMGeAjd/sr7KGTns/
lOVI8RrOJ07d2O8A0rNezGViZKXg5viFR2WKemYN09LDtcpEzZ+BEzPnt4D3yKx7ZxHbSantFsbv
VqM03MZI3pL/iwcRkd4ZL//jEDeW/9xPQm71vN7zVybM3qeiFwfenS3iQJQumi7s1CyUYfMNdXWY
tkSQqLYwMxbIXYN5HuBCuoR/L5+vWpMieRp0HZZWQxjS4COrQ/bmcUketG4JEFoY36IwgQZZnIeB
45oFll04AlZ5yUnN/eqCLC4YUxO7+Jl6KZ77p3KnA+uTwEgF1ahKMxc9/KjgVLLXxbD7k4PE6Ahr
cDUOY2sx3rzA5gXg7Y8VieFjjpbWWNyftZcADUJZzygCs4keA/+haJDnO5ia9XqC/biUBak5tQBZ
eW+qiCe2yB8J5u6gPuvzA2bD7M4nbJjjjt7sSVYFDQ+TKL1bHpkH8A/EC9xfgO3KGl7MxdVdZ+cP
E9dhlrkmSP7+PK3iOPilagggPzaqu7/s4ZEjxhh0rRqrVG9Dw+GRLy1P2tz47FPwjPCQuKwQZAUH
j1JmE+CMtcwsm3ZHiD12zQQR2JmyS39rLwrzAycio9HYuWC219BGrH0tY/+/oz0Lf6TdanWOwZUO
71YU3h22TPBVWlUioC7PUHoEfoHGCvWZmxpWdeCVDmvM7E8Xov0HkLQ41cx06FYutsgGY2WL6Cn9
ciuY6QtUrgTBSojQN/DYKq7L+18Qh/CdTQIIQTk5gPJQI3qNlYMKo/3uPjATo/fsBgtblqtGJyjj
GiuUCi6bQysq9pRe568mioXT1jSm/pxQ6nwCsRLpMv7YaEm6L8c2wtSh4DZG4OMPMWLhLLVhjhfZ
eioiXKnlLbqi1+0XffzU7Y9bmeYLj9Lfw46NT5KaSkaLSmZ9YzCDgwT2dogIDT/k6Ye2CjwMY5fy
3CRdyhEY9RvySZXruAyNTQp3zgmv3wITmosadHyGqh4gka0NdXkWfjwmiGB5L3Vjak3IyLpk3wt1
+ccFSmmyLunBP71oQr+/bVpYAoWULclrgcMVuxQvnNAxxmmk916wdHtOYj/nxX2HbmJx3qOs7gKX
DnVTkLPb2DmpQvcaFLyxuQpi6X7YCDAIBKULZ0k5zZRXgTITZvNSDxP8vH7GEEuuPmXW0P3PmKZY
aAug1dK1M1aZPSun/9Hrt8bdL/CLru4ue3YS4nwUQn2RVLkdJO1AhFyuFH/J+q+k/EQDlKhgG6Bc
rXSql7Yj1yjkXLM3kNb7AKkMzdzuNddKCy0mF3XxEHr5JR4XPLkqCZG1uKXS+i8tq1GTadtdM6KL
+bKLFhDrd4NAjp6qFKWmuMKlcFqZA97WVHaUEkQliutJf8s67Iun9xA11fxxO1l/QQifuI8FTVSo
D2pT8vttRM9HsDQZTCX36MSjOT1vIk2OvO2E1yKGtGR28Ubl+p1T/SZRyMnx84q2PoQCeM35WY47
F3uYa7uAWPeG4cVCDlYEHSgHitd1XtJJbhpzN2oSdBI9CXuNhf/XaRuI0Vk90MTtKYbvbj//v8ja
o6f0SeJ2iOwJJBR5a6xTjWf9LelrT8jYrPMbeUf6yytl/pKj2G5JJPtBynhFeMKJeTWvm3e5kTEw
tWGlB6ojkqSspAmj0tqMLdJH/TkfuZzHgNupGEi4sTJ9oSeepC64gCG4Ml6gLKf1tqfZEiPS1BrS
QRrW6VBjwjAzBUtVvS75ZtFDQOhKXGgWmSMOnPyYDmLLfA69Lga/+iPKlLDM4KlR3fQUCP5xzyU6
3beettR1Rj7m5n9sik976nk6KURiIcwgB8ZeDYgPB744UsfLj8z1z/aCLj61sJXDnlt5dY5jAec2
Eh9+mQJXTrrlMSWdt4OyN6tH+SzDQvCRbAWHWj98xw2qpRZsN/YmuGJTMml2WNvqAVlOoFFlVogi
XL+OUsdU9ARouFEVi5nmp5PZCjnKg5gRF7vUo/u6CyLu5RiDy9O+AqFGDlR250ShBJVdTSnCKDeJ
WcUiOMKUCirgwRpUHdcrj69HJUFIgAz7TEul2WiFy3kLXdTZpA6U1TcfQk5grXG7KMoZUxffpKlF
/Z99+wavkrLuRkhroaDH34rlWiI5DHiI9/7y+Zy1QvFtCuI3pLKghtnlTkXV+i5Qn0SYjhaNm1AH
U/r+9dwZxDAceMN+J32OWgmCkWcrG8M0NtoW3VxmwK7s+BwR0Mqe+CpZM+1TjRmG/oExXDgBbldQ
bMdWXLJLEWin0C+yJSloqRmeSni+vyygq3aJqwBMf0EYViwCFMK+H1kEmy6x77z0py5ANYmp7arQ
dfisMRqlod0fwXXA6c+ftZz8IpyHaaHY7NF+erLxpaRAYhrrJLGJECi/X1IQCJdI6+DJylIblgGL
W6Lwpl9zRAMAHVmlHnsk81t22bbyasyR6QadfQo35sC+A2x/s4zwaWGH9n8NUVbKXU+Tcv5wpAiV
upk8g8bgp4DuLTYqkp5nfHz63VAOO0j9vg9bfXRFD139p6dX0vJ7HuzIiwXFvitH2wh5gudpysJN
625JJgA6Fkn3cs8kYqa3SG0oq8V7F2RKm70Ayuw4hxHpRK9qNm8lcNbm+Wx6QiU7zPlPr5qiJxvx
xJglzXxzRKfda3SJ8xFs9JVFy6PrR7uic3fnLQbNA/DTKhyJMCiLIrXV8k/zQq8mRgZ9fz+nFzpx
Ks0x7JzCfd74zDTCzXecQfHb2T7YI1FmLiX4cE7OQEGXYZzeQFEkM0OsuigwPolGKSdOcAf+93Wx
Els4d6Hhi6iPoNaNYjeGtMx3v0AGnqGp6bUkJvx9GcPZU+2s5KqhTRbpd5gRiwz0YcbVHOdLyQEe
QXx+n1ykzr7prKIwN1LP/Ef4Yvp7mX/APuZ2VT+lw1VL11E4pLoN5FHG6vMINfWzgIAb5ALA6hb9
lRbVQB/j1ucYClOITRQE/dm3QkrYPk7Z34G2upQjpwA0VzImfzHB+jeTpUlyxjntbRtPB0GbaOxX
iO1kaSVj3GVRj3CT+PwnmY/mHUw1tJv2DYP5vRM+3m3gtmJU1MVck0L/KYsqx5amktSkwYhbPeNu
+WcQmJU12MX5uS7ocZ2jqOjuRPDT48hDZOa93p3+79yU0CcL1ixRWFKshv89oCjmsDXIGyLqhYIZ
y3BZ86c9QBD5m7Pilxe2ThPWHwwZ3ImhiHcSywtUAfnwoyXFAV9hLdd/ECoNzWt/g8PL89e82Xa0
ZZssYJITybUbnwYfffUvYrixtmt5jhzMNaEo8ky950Ag53E55FdJQp+NgzW6jawbjNOrP3I5ZIlB
n2Bb8vawJKPAbMh9uZFQHD2FwOgtSbw6ZyqYh5e8cUts+9Z1Df7zdjGlDrruXXKEWBjf6+YbNQav
J1aR8OfWylVGNE2tya1Z0eQjcqNCqe1bSGyeCZzxIld61jcXK4wA51lIiS6WIQxBIC0Ifedr5sDv
vCGoRvxhixMewr0rifREdvfgLpzTwfrzgpv3avi5JQxv1j1FBpcHGvzCqZwVr5J1T9wZgE4iV5sQ
fyfIk0ePaLsrBqkmHdu5FYlVnITg/7k8I4WRGvH9g9YJcL/Mq+rWIO5sRSBsdg4msWhZ2CgSJ8nD
Uh8SuiNu1di2usWhdEQ9EFtY1hYLycT2uaN8h/gNAI6T9whwZbNsnFMyFrcPRFLRlnyK0HC4j2kY
dxRSp9YTFrkqQYRXqhDZDbKR/94o7a2Xg8LA5kunQFj/Kd64qjt1gXv49bCwdGC7QURNH09p1XKX
45KWi3UkRANZJmNskzoXdpvrP0XcvTXDm1E3xdzPpDZNaScYXDTxCgwO1u5yoMNRqmXRhfYC57rC
qu5HHu4QuMxz1c8G9mvX3wKc6GVNyKvdH2azF6wKPx5+oS+U3Ru7Qnfi/vdLcMiOHsmK4F+A6CLc
bJFtqdbKduKcz+APTYA2NgxrPHCu9r4+q/OBTlse4YaiBqyuGCq5FDFO1zUAko105spyxfZLNvrM
x3YalP/Yyyqr8iuEFO0IpKk+hG38a7YP5FRpc4Rq1YdPcGCogGkVG4Lr2sliaYeJOkk+DxOkcNI7
1nzX09A330/vnOXmcZqKKJ/5qbFaUr9LgDxAUPjAcINMBhGhr2DbL9mzoHyVMFCdF9ngo/sGZ0+E
w1qfnalZfM/FjemMjzgsBBLthNlRU/cgdqPJUVb6qbrlHhNvcBlAdvCEvHlmfo2OWVLvwtLPX1Mx
c/NJsPMDl3GULybu2KIDOzASgXy9eLd6CNixzS419P1jXjz41GTZMyC2ZZYmRZAUFCDHh0lyxrQP
I0spRWtFm8JspxGLyvz0ytlih6HHlP5ibzvfkYGlcrTHwaDnJIPyzqu82g28FBXfLO97ayKwMQQI
E0Gco8Ia8sOgNhz1CNsmwXIrLtChJZfsAc4D+fNlPnLJrJ+s9Lh3NKehCcdjk4Rlp1AlRd0IWAe2
ES8tMIjcrbaAvjSLQsrnqewhJ6nTwx4Vi7xKDJRLdu5YffhqRPAYG78mjIHOrYQpRBFU3lA/x0A+
FE4ZCjaugTfAZcM5ycfh4r+iJwYYJo8XF0TXA8exaWOMPOCgQd3lT3JWoDoznLDhUj/Zdw4Y40IS
LTxWnDOzhqQS0e/fdx1bpPjcS2LMNOO5EMMTZaF7nl+s1osRgh1+ftk3++A2Ozw5mkI1bi9AnWQK
WiUtqLnAcRKby7gMwo3+gLuyLnrSrtKO5Bs/405+Nx69QTW6y89id5eyNLsK09ychPpVpCa7Eyuy
k3An4Gs5O4qTeO+x+s+r0ujXI+N/fq/tK/nBEYOps8B7ioQC7bL7vS3ThFs8TbdzIryNm5C+Appa
NENPHOsnQMFjxGaZcs+5ZfiSm6Apfgt6DqOQNUGIe/+7xDKj3FzSmna3t9poQ6AGAnHTuORLP6ky
rIMkmy+l+jhf5n9Px80XSEh5rdXnLZeQX0vIBTntyhAd6EBuUCzhmIAG69G9wvWggSTiu1qgL1jd
7oWIMCuu6ZmLNOShS3eZ2mC8U1DcFtx9p3IOD1t43MDIszSq0LR4Vbf3w6DxAbYoy4uxvEk7UPH8
mA1pQ76CoqDdPOngVAV4k5LZjB3EJXIQIE2pI5RhfKytc+iPKLi/N489MF/r9lebvufSf5CfdSrH
ecFssPzcEDnFevg9Q5g4oajruFSILKSKNqP8jIbU1WbrKtIRh1aI+GgxXzJCgoGRjMvWp70iruRG
DHlBmH3JOgSyJj1UPwBYbhwTkfn5pTcy24kVzkRjNi8wh//WyRviJa4fI3VBySgutksOJQ7VpAzk
E6hryzkH2GDhwD0hE1fWhdk9FXfOAriaX8Et1XGeINHNToh9Y+fFqL0mu+3qCJzlEMHVmZd7o4Oh
c3erKObPtcOC0ZF6lauhOP39HX2c2eWB8LKH7r7cNri9taHC1L+g2tYKa3q6vpOZ6V2I0yQUQ1S5
RG2+dYBLNdiKQSQkgNs0E5LQj1DM3qMPeuLSxgkjzrTF/EAs05kycxk245HOyjNi88e3zlL9ZVZn
4OwF/H9ix4dcDjVz12WraLpb4d0FtLJqiDaApuT8Vw7Wd6lfF7hmNjdiBxaovo+vi7zLfMBOmiUd
Y/Vazcdic3jpCJfzjJlUDceRlu8Y7gNVsBeahY/fDtTEZQ58to7nKcwGNJL7oL39uEcoKY9R/Ykz
HFco++OrGOXr3Y8Xbz01XDRDPGr9oBc2RGgQ4QPdPQ4Rlu/8mYGXi3UcCvan+UJ1RpCkE5j6Ohtb
Pj+xx6DK/wnNISSKg+uEwTB0etzlDlmf/nRdJDGdrZRIVfXgvg1Jv2E7DEPYkaBXgsvzXd8cokBo
Mxta5VvOntLwpK5+faCvDk/g2VQn+SrfUzt7nMt4BC1mftfN8icpDBrPdyqobGAkaV8OhnZJ4iWc
ueI8DeRcSkFjXN1TYfnIm9I87itABGypoSFDhVQEa/qJE6DILsO3G4tuUi6KWHW1+hqSNWZGiTQ5
ogBNejnMIk5fRuLxtjdcIjg28ygfAYbkOdOEaJaYs+xr4Pb6otmjkys2MKh45UYmhEKtxW1jvGq8
PCHyFKYdcYwxj3Jk3vjKXsL3fkAjTu/SPs4aShqRGAAxw/PqRZnJDVU6bxkShyh6GDpAdrdONNf1
oiGjKt3sH7IrCnd/ctoy174rl2N4jGbGKZIfXx5m6sPx5yaT4LAE4av4tgbIY8jNM+xrPzNhOGiA
6WuK4zlqdeaeZzN67VRfs3g5Jy9aZeovQVPnaDcynytUpqKGP9Pl//k5QltS053o6cHBP/rU/91D
B+QjW+wwsc4J9TZsnpHDoS708CrWiUiXJLLigvaoRFKO2EtgPXobcs8W0B/mv9ZFMn2/m1amCYoI
rIsR7ne2A2Ar+hxWfOpIz9AOnEqN707rVrcUcIlE/oMY34j1Qp9W5Wval9Kr56Iwz7cesI/4h/wo
SR09oACCvFk17KxY24fHy07wBmvXK4VFyA62nmVSfbzE6TWXy2vZVjNWvP4Z5GqP0lSF8cWBH784
o8t0u9WL0V5PHJi0xRwaqSLllip8m2GBwSd/IUO0dUGEt4C60RLb/i4DlbezuEj+uiq9q9DDDOpA
vWYk+3rGOgo5dPu5V5onKvsIMtz9K6Hcf12CrWjDIAGbtuvwwOiRwuAoEFUFWdd5BVXlbvULgruJ
za6gR7auhRRFDfPzbnO002/poPcMfjjkWRYW+qfhJIFz04VUqH0hikNn31SWrTYF9RNdbarWfXPK
YK6np+FxnNsGkEsER4dlfIMhZKdUGTG45lSvl0JGWO/Vyb307jrLu58Qm/er4iM3fyZCY7AuS/pl
aDXQ/iyYHdDy6x5OsZeUU+XxQjRSQf5e3Vpgy3AokdSvY6nalZPOZXxLHqW+Z2Is3St5tbdcp0xd
n/PmjyUaTAf6NioGla2tC+lYPpOsi3MvxWZBTyc3HgP0M8Jvb2vKu7V30cJshp4TI7arMRf763IV
aGMvZy2RpqXrh0YG5/gz+gnYMjuM+eVfhWETF6ool0uQYJlSZngzsS2wEKmes6RU3TmyCWOSupLO
JEpSNugXk0JPSqEEhtMv58aDYoCp2QpcWc5NsXWo0EHWP4NfiXZ90JnKOi4M/YVh5pBYJK7wEsC3
FvWyam4fkAiFb/Jp2hZ9RIIQp4B9kVCiQ5ebJFm1ulPKELrP45pL8mkQwda8SukhKose8sCl0qEQ
AijpE56ayUWCjX44tn0DGwX9UA3aglqlTcd8Twq7cKvxGU94iSeokx+3YpN0MAxJd8JoAi0EdnYr
t/m4Mnswc8egzLF/YeVegGjMjb8ix3Ki4J2L3hFIdT9ZhzEjgMk40HlX8AkNxztq1jEC0D8Sd/yr
m2oGmIQ2yyOmgORESr2lXZ271wJIs8K2gHY4L31fZB8//NLfrak/3AfOnqHqxvAoxU/ehKPSYI/A
KjqfF0C7DMFdFFRIehPGAm9xsNzBGq0MOCtaI+5DEbGHeM84VI5ERalI1+XMmMn+eLJoWvEq/sP2
hum8NjA787BBeNukqnmF8hmLFXxN01rgBG998Y33yJxn4jO1sTOVMIzFHEUO6CXNo45K3AjZBtwg
vqGU5b/eMaPsfP10DunFa4glIERBGFQP8mpe2u1Rml8hkp8aE2KtT0NzvnYKkePGnzk04JS4nHP/
+hISs8+LxjW5zSG7BONyAMNJMaldI2QlA4wc2zyAuOk5l/NKA764AiZLF4KevwbrCef6iBEa70gD
oWJZjl2TMbArHzp64SQux8/e1GxNYuzWxUUOKjiZvaathr+/z2mk1pyqIrE7qKxCl6BroNjsxvD7
TKkyjELQ01G2I+jqZKuFU2q6IzhIA20mZWo/65flzACVn68NJHLunB9jy6mz5Fp1lAQz5o+DC7cY
fIevvWVSsFJTG7ba6XQgn7xa2Kc++X3KXzuvEH5TVrv5H7Ew2wTNemiYJKaXiCCGs/AiHAhkLkH5
9xNFfAz/7ixjBbz6AcRmNAVHVGBFMVCoAC+EgpuqXrF2S/rUkXT6r9WDYCqwtxP1Vs+xAc7W610n
QGxKdJySFMO3CKQitOlFAsSGtLGR+z7YSzKeHkVjF4fgR8WN3vkM2lrdQH4uKZvaXKTodpRetwk7
gAseygVuJbfSDzfXb8LRQEk0pDZUlV1qPC90VUz+FvWTQwMs4gsan79zA0Oj6eEnJl1aWjywGVP8
J/Erjo95VKGh7nc3rGgVzysmHzehPGa5c977XdhdAtUn8vp8Vx6anZyM+Xt60ka6snQxbUjgKVx6
3LYvBvmoN1H+B7nxCyWK+4Fpo5GLe3Thjj0VEdlASagjoEI+W8HAUfbQn8K9t4qvAUsKq5eMnqeM
CjszeJCeLZWZoDIjrWDUOGTVcZ0o6LS+63daoCTDgVZQsODDH9ebgUjujUr0SXd+nSt+hrsbsXy9
eHhjvGwxZJz+esFSsN5qNHCzRB/w+/rDCgxxPaL+ajCkVo0ERuyN36dxTKiUBYLegFH5WghvMXF3
MbLZ9tVVm4ORCx+Nvr4cIkNUJJm1AizHF4yLs+YH0fmTDNZi6HMob8xTDp1RKtKPZMSKvQULjwhA
E8D+M30JMM5VIxj3SQs5OQAV8k0YaQJ6k77JAttYZClzBkI7Dw7l0msuNIYTcAd4iJCLqjpdLSnX
i6GvUo/N7GZalkcnC57o4W09twBBjXPuKHTLftuZiSRE57zf/IXtWbuTvqayJmtevAqc4R62+/cg
+UA5XESsDZObC9IWsFkcCuPWyn8/NZequS7yoAkTkqHkFyjKR29bB6Anf4JdCp1YQu0CtC7LgHM1
hBCAqJq4xGMbCMage+YIrkX7zm+GSMm83amdIPuptoKMqCbNzLc1JvAh33rAqF+QXb8FZnlO4p2h
nrmRYlx3Xn36+YaVZZO7kDaizEO7iFlcSqPeDhBHeVas5dpIQ+40LT9/D3nAblgqY0lN9qK1lBtv
7zz3HMNejcYAz7wI5Glo1cnPR8SVHuk5h3BHzqmw6sEnxMXXWZz48JvcgjMy2ZzmmQSK3CSnspoj
Kbop9TrkQAgVhbThIbJJhzgJiQ1PfB+8OIBGlqTxDhzWmxEOZMmEM+JcBPqmo1f2ogtwWn4BN93B
UA+XMRsQeALUkYF9RGYa/+rzFlCbPpGmIYBmujejZ8POIX+HK5dhBOSTLkG+/OhrGdKgJVyRBNe2
sEu2FkTOGixTzvQyiv7eWUse0NvYZnqP0kQAfh9W7AGZcpzw5uWpBq63FvHtHehCdXYoHRVtEsE6
s4JP6fGdTJp807dsRpAnP55LyZ4pkCEdQKxsl1KtgudQAik0QrgH0tiuiYupto/u1ZewvpBaiKk4
pQKrpM2L/ieFGoEAmEV4L5OJaWAkuqW0BVbmKEdLrzWiVKPUj+xoIvZB6RnVFlhHq/9jI5OdJ/yp
5qm9rCbCSgrDKCeiGHi28KY8kN4yIT/kYoigaGuj2VhjXNEa003filsKuBNPFCiS0PUPU9cmVOaf
Nnm9tarcJ2RGUjCchX+iXgiyN5R430dtMEtMfqQbwy2f0xESFRIi0iREyqo6X/OjrAVZujjm5TWI
KZgY9FLm+qyzW81xPApNHC1KHY3hjec4Y58w1yoX0lsh9BT8qv3jIuquTS0h9V5+IcCVl2JGq3ZQ
fLNiVHWnZZSmpsdYDSWWu3WrEeFUZVeE2YEGUdKi4R1khyjqe13EtMupHGE89PcBib+9GeV3eJdu
icqZPybNik7D7VyofN0MchdsEXzVQUBQvnz+HIZaeUD7pAsEsrM7QdGtaaUZUJQ1aTebS8aqnQ8y
SQ8fY9ziJ4jipLKb6QSB0CmPG8cF+In4JbpjauN9Yiy5mtCbXuPNXBk+Do11mEQnb9tbsGqjXQe5
M0Me3esY14nUHXxvjfOHeAILS8Z+cHov8JRqYH4h/wHe1soxQVJQuu5HU71ZeRo92wce0h2ubcRG
abQmXyfMe7xQH57uLGC3A5cfbkg++n3jC/ga0+3meykgt7A8Ni9QKxIXpdeivbwb1ksSa7VQOYsT
AfkYMzylIn3wct2GFNbHuY7n4zmYFbbjqU4UPNosULhNi1kk5hKCkCZ2jqonfZb77DHksECUEfgC
3NcHzyuZcpBz9bKld2IWobIAomkdRcKGMpWGp9jZjWzg8ZLuO8hsOMza9D2fey9LO2xWLyeHO3r+
jwUMkR14+VC6LRXHQLugHUoo8mdqm3rY2EDmALeZHQ+0Yev35bwRc0jSx88NdVscc9kLZ922w/6w
ToT/xMcJxCrk/5Ixi5NyV/yywrnG+ujzZ98bEGI3KSCItunZrIAQiXtuGsau9777w/Lbi8HB8xwe
sTkKNSYw5m2o8Egqw6yzf5n0qyE3ECeueM7E4Ty5qDV4TWI8HuzPNveEePN8v+PYVx4xUltIoGjM
qZ/4o5qCJzzo/PO3dcuWjr1FeRbQnDd84AvSWM+8Rc/jdI7ndylbl8Ga1jU0J6gJ5mnkzrM+qlg/
KLHdKqVuPB6eCxXqv5j9KTCEAawz/4Y7WQEvN3RPgk/zS4n96ALNQTdzavt2fQyD75Lu5vpp3gI2
F/s8rSeAb97VYHFw2fGsbftLkx6GS6lCxNFAFPs6iFtktFCCs95MkoeC9nZByE9bsvIjIDZB2r2U
DltpoFtnuwuRNwM+btNag62Rryon6PV1wUrhKTHZ1KvzxXurWvXjMavsYKwNjQ8LlJsJhMoT7QK5
Kcw82FWi5U9esrFyEK6HMQnv/hnUZz4w6CuCzbzC1uWRZNB+FYpaWyvUYK4DFZlWKL5mdBF38g2r
OgojPCvehHkPhXzMs882ikUzyu1FcCLHT6/9rT264cQoKaaOYt27khq6wMtXt1laNW/X+I9MOERk
jqDRBiYuK8MnrwRFlzsNicPappeSduw53rHhl+vc40uy5EWd1hwpcJCzytkgIKkevdqrGLIMF7un
JFsE6Q7yyZ7jfVx73pCAQCv7hbg8BpEnDGbD120D79xTairLPBOeano0n+dg+1fXhh+6+XB7BFBD
Vv7/3FiqFj4UQosw5iqtVm99Y/x0E/0fF3bg7nsWQIkYHkUqCe7nhNaMsKlQPhGRWGi/0B6WIqGC
tqY/rtk1chWnCK/WiDePcWiWM7cA+gQ5jYuzTfrOJI4uMc5pyV0736DoRaJwlASH5x+TWISXVISe
rHHG7XLqwslFUHq3ZJUgYRpqAASnPr0NgQuYOkO7c2kdtWf/MxVWd67OON+KU7wPYnbqh5R7tXiG
9yV5wEEMWD9DMP+UItxXUrESKlXrGYfnD/4CRf05QC0fLgsrmU+0XQyoKcoRGyBHZVqPIWA959Wf
y+0NPPQXnv2mZ+SCbpIebu9dgA4nQZ26k4Tly/IvGSytw8rA7ARjaEr9ENyGd4Bdf71FXL8NMYSV
xvjiZak8qtPm/jcuXNc8aClrh/xH5BqQG+ePbmlrwrc8TvduKD19zIw/ZwCk7DvFofwbKFigx+21
9sigVpM4rTHBK53QLRnhs/nwj3TRiE3nY+YR3PJtBqKelscWTaBgbYyBOcHhpKF+0FxAEBM+2jf4
wPpqk/uHbWrqgvqFRykcYfbBjrK9WZXebP1KB7hKy7ZEHbTTmh1kLo8rL47nowilsynLL/bMZeEH
syEefR4kdFkqwHBU5dpmoJL3WgCwOOZETtC+Sq04HKSg1usId4B+4usHu7gr8SJwYA2yZ5vEP2/Y
uXns0AHH6cIVMr3JleCpF10+Hv3OgC95jme9Tq9oIkxNN6eXfGZXZCmGQnNamBxMuwVLcPSqaOBG
vdUOrEG2gZDsbhRcStBI7Nvfb+Pz3rsW7kT89SHGFr+pxC9jbvhZZESBeSq/J8urTubgDxtjpz4C
mTB+S/KuArQvPEKYTIZX2Dt08l1w8Fp1r+c1L8rWrCtOfnhHmPDZS9Q4j1xSFVLcHuTGgBsqKJFH
bfyFQAMKwU1bhYtCKbcOPFC+mLF6eqsdYl6SKE3qqAlSoE1XIZArPSg6hsNz27cLsk3dplnk0as3
6+hZuBY6SU6njBMot4Jewq24Pc0DThxbFpOJl0AmxhqdnVqR94lBFECLTdObWZ+P2K4Q/OinzB5b
Kv05UWmz5MjzX/JqKwfR7kUM00IexOwditz8NIsEgsJv5oRcsfZ4pS+mUN64UPJhxLFZvYnwHWrh
C/b1OqcmvDWM+OPOuIEo4v/4sgkOsukIJrs/9u2x8AL6lCcOU3OWBgr+o8J7xeL0Uaf2rrPg5roJ
GfF4C5fd5ebeLdv1O16qVc/UjiSocVNipzLnlCJ9rP7pVaJE3PMe+uaa903j5/8iKjkC+Uclta/n
icJglAx0g9H7uIvDVjUyvz/kUDCKHgeNKw3g4weVTeORz+DbQQDp91QDcynXBY1ab6WGYU++nApb
ntemX6EaLJkhG8nzvzn+QyIxdJs9icxuSNhvAF648REmVGVsWVCoOWv1aAPz+161s4DenYxb9xfB
MpnZbmfoHIQ7KF3Ww0yvX35zV8x5DM3H2HHohU6nBbSxpFH+rmA3jqMtnQybqK6T7Q+VWlnrpK84
CBiL4YPXl/h5Pc2+J7lCZR86PeCVZz0rkNxFizqfFiID3HVCV5efqmP5tOu1oVMN+PYZJlNQWrix
/Cv0aeSnk+YBQ5MdLSqUVR355kWXffjF+ooQG+iy1HxwBi2KQRJOmPWTd1D00u0+yRKsOURLrMY1
G3vWdXT6T4P+cye+nm9X0HuxvZeVLMttmCjaxb39GctDCKZECzGEIk4nvGq/aL2ivSuNyOJUlROX
bZj5tolu/VJmf/9Amo0J7bevYddBVCz/oyFuFuwqsIVpdx3EIHFDF5Q+Skh7MCwI+Dr3sAQYv1pn
EtY7Yrw2JGZJ7hfvTrCb6kiNvVKpTP3Ug82Q2pBuaUryZpX6KWtpOrFf+jbhXPXsDzPD9ba711+C
u70WCLzVvOehJ8VI9ivV//LjcDAUZPCpGP4QJWJTPlCWeS77Jyi/Ejbh5kHAluGPx9Lk8FC1qOHf
/iCo5828XLAcKTjM8UkoNskbr9gQ4WaKO0pLniI/QsxfdhaXxNjuMYp2HevN4xCWWSAd41benUra
vg/qmi/YgHgbI8Wu+5w7inNtOhKBKe+uqeN7Or3sn96sa4kkHEtawc68HtecuOvu0On8LgpDNfg4
t/aCbNYw2E1gldyP2uwFgs/qpU4c/8nqHTjjiqmm8GtMJ3KUwidszJkhBU2Cp1ETVwCGHB9j3uhb
yTWs2ptyAtBOn1jGe0L+f2PsXPQdu5ST2xK0JIUX9fX3+ymxQRdrlCO13D6UkOeniUgv6LzCxcxW
9kKyCZ9VSks0wAM1Xs72dWRzmwMMyi/Jz8iOGX6NngeAq3YxF0A7Rsoxox6KXgSv2LIgGNjQrp+1
LFvzVz5rsBus1OCNCIxYywqxra1mqAEEMLjRVLk9xrlVBFR4QzwAKHSHWgFJeXAPF+PLldCW8vRw
9q7etFZ6NG0MsTFd06bUi+xrGxo+sxizZMX8wuPompiaL7/xXEKYU6oGMD9cEugVd1t9cyEom+Jr
stuEsE9LhZWsgkDc5GwNe9JEkk1CjHIBSZ0rcIwqpmBOC6KrCX8vefAovF+rc9RqslHQ5cso9/YT
Wk9O4GPXwU0iN6iBCFprK4LGwesLHIsrA4KzLZJiARBCo4OOGAU8PytmJFqwXBOFq5aKPqzmJ3Zc
pOVJVxoUmAt/ys3fHeS1nOGVl8Ijh+PpLQAiHfR5Jeg5vekoVIVNJn+AlMiJ/vAX5krOqDp8SjQb
TAwbI0O1/FpVJe3yWJYO6wFLRzdBBCbZ1ypzoivjGkCRM6YYJ992b74ccbCUyYid+Hw/1a6vNvkU
+A3yJrAKtbTxQmHLnmfPzpABZb9hOdGW9T4VPQOD1D5dah8WUUVGZKLFahVL68AMU1tS2nVyFqTS
h2O0sKEcc9gUlUa5S5MQHmds3MQrVvq8iFafHiyT2rqDv36ycWczVFwdfnqXHsp0FLbwj3IUDkxU
aNt4vDGS9+hKCFatoTsuS4hvOEQGQ/8TtnVgBV9Hmyh6icOqHb88eVGk/AIkH+IQ5d1W8IR23XiV
7jSWEILzBrmRuUXusJkSShQcb/l2Z6/4J7mAXVijSL0Oyg14JkXtWLO45Xe70z290p7W0fEftt1p
XGJG9MiO+sW0qLhRI66psM7OOKO0zV9dkbguCCwcYJVSEGLNMlWa3jXtysCzE3aUhp19SWWw2/VW
W2wyxWdbimO7qBmaGjgURfezYsI/BtPA2bIzGbHMSZ0fNB5kVIOhda227m715/pNwdKFAf4uHFFj
MnoSLmXnRDmQsCT1ZQ6XZL8S8GjCIhMoFW3M8PKhGPYENH2PKboUOjemRBAgt1E9xnj3nKJXKPkS
+LM3wp/x4bJ7yoXx5bJPGUie2aMSqcY/M82kS8mQe8/LF0SQgRbbGnFm81uVjqJPms2uUbHwMEHx
hgdI1enFcxvVqMqPV0wJiFO2gzRUxnyYuoTbNa69Pn1BS7l3QB1tHNsoWMJICPNl4PPPIaPkL81+
Gl4e2ZBZuruDiBdcKU4lztyor3BYZtZuBdUE5Y2NMHpg2Ov8uFEFr+hoAWsrbD2De7NEokdQLmlG
xpQzM+ZYGVy4bmUjeQVe+6q0Lf/KSY1HH2aXjxXLYh6hTTSygk2XvyB+zfT2Ig/baO0cU8iybWBl
aaixHYWlwLyrCKUbSCUA6Ua4ITqiCDJRA74VI7tfBse+cjjqYutiK/ZzX6v1K7+Xpe0gfVHQrIw5
zWktMe8D0jOEk2Js/QUWT+jSPXQLbsiSGRT/AA0FQqoRVPKa7/Aeb+FSPZhIH9GU2Mh2Bp32DZEB
enB1qfKOfoaUi3paDTLwdwmyEHhX48g0EugOz/g8n3EVRendJ5aSdKro/smFtYXlo1QFcwWjY4Ao
V28EEW+ZwMyg1Fn4DOe1d+/iT7dAnuJW1oYee7tBdwqV6zZe+5H3kGz5HZ6nkPKTEdlabTojhnf8
ZfuFAYJvJ7FQ+TCgMBHFbLcqkbx73cdrAZNzs86imjkUSc6fsZ53gayWD5mrpC8wVY5cgINvB4qV
st46Lv97YEQcoKcj8fOFpuWnaKjdDzqwLCyeFc6U3daBpaFfBx3JFoMUJc2mAX+AXmgBSlxK6PH6
2ISBerY7euL7lFsmMVxAMr6QACvwq7Z6hcxnrfmWg6qUXyBgI1Gd5QyNGzbtKz1UxGUG6lwA0TqT
AY/conasYLxt7jXWnI+w85otzF5V46DNkrbsJfWBzxm9HgGqoVXtxNWQ8QlUDPpvVac01ThAv1ST
yJo6hBKKems9LA7mz9pcXFbIjgNpQJoor3zuCUBjPbw8E3kJY1gqJn13Y+NAxUOxxk+v9mBqmno1
YzgOYx23b9nSixzHr70gcpTIN3bVtaJkQSt9Q2clqoRLSRXIYiTo+xL5X9pR8g0vJCtVgPW/oHlj
+6HvN+rNmirgX7o4G8GY/7X/1g2hSOMgPb4b4u96vFmWyJtAqrCzldO4m3u27InRIyNHnc0X9IIA
0k7cy3V+5Bs08M2LXmRB58aXiVfOQBJbKQIP9mpJO+DFvj7Wky72lOKCcpocpU0Wg78jegBBrUqV
nJpG8QT/NbPSS52KB6zOAnrTkyXO9o4YPBlpoF1YvAT7qL8vJtn1CSDc3PVY8RN1blPdJk/xbZ+T
+9qdExyJeHG2Jh456v8HzXCciyXURHWLBnXnxGYleBA2222EBwatEkfEmv5PlE6MkT5TT3FxT6Ai
JzWPEIkah1FtmxDsPi1taVmjmpAeRtE4g6SlRFNaWwjTKIrHbmX3IRhKx4YKteWgHUtCPR3LhBDe
L8FEzsw69PAPh92mRelEjvp2IEAlUC90FntSf7l3eYmceIRobpO4jltM++jSIufz7d0gr5XvUlSP
nGSH6hFCK2WvPhdV0Ym4CraBXyoztanv+qGu523jhhqaYTVU0OXAfrNslQBB0qsWo3tuJLpOzqFA
Li6NhF48sOLLxsYjN4N24vDcFirOiyR6/BCL4uZsenio/7cvy5oUfpEIBwb4LXyT3JlORoejpWrg
YJ/Kpks80SFEyQm7uJza/klmA/siXaaHShQRYsXIwq3lNClD1gP/JrsXaXb9tVlQmRdAr/Izc6QW
OCyGWC5mL9PnEf5ejXoJiz0BdLYe/6g0xDwq+w4uGxaMSXeDtOSaukU7MwfZWFkAalHi4lSoYpNf
1We/oiCeKC6wek6gIavDCF6pwXM4adF+B2IctZcP+dotV6oGr/xDFiWkXH1wY0QsBnp5gEy3ZZdK
x009HIonK8xo7Xf1H1QvqfJ54lCiNdkKtmuXmUcDAmuXvqMeCJU8Rs6v+AIDZyc+9v5xlRAFti9l
N3uJ8yLSG2s5/IbokhdrV7X0CFm6y6ih7UfK3oTzzZGP5hpdKb4eD9c32upXxEE/VNTq99Y64J0v
ao4onmbsLTeG8xSnHgqYkZbMEqWhDFkmAN2PjyCWrZRyll5zXA5pMUZ0ne4m0nuNgMnmd2Vw+yr3
5z69ZW9F51W6NSH4eyXRUSk2lj3joBhvmfaVawg1OdQLlVOSmeyusyZXtsecKlXYNgRF/YSlx3pv
+UjWEwneKJ2Wu/jZ31j9MmTy9X/QIlZYeNQt3LtNqsYMVe0NjDmZVzy53VNLAx95SURLj8UiAcWE
N8/Nm9hURzhoZrOzobqK7QyN4NziW1dETG/K8ctWhUQp5RbPk3bfJl8EBpyd2Bm6zpFozW4Q57Vx
YIKKvbrPG7kLvdfLgr8x/suagiDIJaeSBUoNt751x35kdtmxgM9fJLAnS+Rtra5JFRCjbv5qtuDb
BqpZIfSiLYYEiyQWjs5cSCsZgrSiMk65wuiDnpvrKdCXvyQePxI0NEFN3XjjGBu1xuF8snDgAJoW
3T2telNKEnhLb841dXyBI860p+7suzLSSGj+ZAjWdJ/Iu5qaIcI01YARg7aV2FieWFHOhbECxtQb
D9M9TrMrgTdmHRlsxZHRgnWJOjkznQtqvhZ4/DEMg0FncXa4kGmVU6ViUFJonrtyBWXVXgObLzYr
8VLk0T7qvN+SUMFi0i6q/0IHuSNjoQdh35XZcUtmXu5uGq9sQbGMbs2safmww/67Eyj3tWC7xV5Q
ebqow0iM7APDtuU32HLzGnd8Ef4HKbjsI80bhasZcyWpLZ78E77RUZkCZXHq0VqvE1OOL3jv0hCY
YGfcBolz8NE2zP+acQEwOpgKcCMe2qYH73DTVpB9Wtvze5Hey5i1yJ4nqEW3NE5eXP/y03GeHGOS
aCSiy12dCA2CfyzZoT50RYe1ZumzT/wnuHzkLjl+sVSJPRlpQR28HsXMgeTAR0cS3U8wutchoX3o
3HN805sUhrtcn/PrjHxoI8FpyEqcsmTPYVom/mDb0WrQDzRyt2BiFKTlF4rdbNpfysV7l0bts387
kFWA8rSK37fWgCxLKaUIGeI87H74o0eDnRuGHbu3H50uKc+M8nwhdQ1nd3OG9fKoT+okaMGsJFpE
YcOOIK9c8vB6DEv/U1KcxeM7m3+Gyx4XRe/O5ok8i2Xcsps4BBWgEIA5yPB1tNJa7rJ4o8+Gjett
362PH4GuSQLWFA3RY+EMYOCV+15e8wM5WSTeWU7GUaTt3SstEqY35HVoRhFX1RhNhW7STWIoCr8/
dbnXot+QJiKZmpbnRmEZphmF9SX1jvUpnVqjSI8UXKo7DNqQMJBrd1E/qEPS8h0DCl+uDrwjGtj9
0r0CpFQ/CHMnHDPiugYDlRawZtA10FMAoXcYcXei+fHeXGG9M+SsKx1deINde2yjLU2WlidCG04o
8h65Hhlh/3ej2xK6bZzJP7/yMByxOr38EaKgNLe74wvYC92/J0FoQwAhzQtQPsISYnVpEXZMYu+3
OSWWuwSnJPPr/pMSwFt5cClFDT6+lRBORhKBaqYocYpAiNNwtf34yP8CG8FOfx69eYMWF8oGFpFA
l4Id3EkcGInWtue3F1VpXvPYghiFxAWTm4I6m/OgBxPKEmPyLrtLogjj8cQ/jY+gdM7WoAWnQzFY
ECvPOnF+rCiL1KoRZKXjQargTQVoaIeRYEFpYOEX0LKPbS24YhQJsp0+wXAiCE6DEolI4ZGb9394
VaXdV6m1b/XqJYmo09MbgydYKZ3S/R7s3cbi2CdPssHWpqCzgEs3FgFY1H2oUyVqzpOkKsXVQkLd
pieb9Y5xyBvIjCGeuINSHcbVWmFK/CY9cOrALxUlvdZQhDSimQnxlBCH5nlxoOOQ/qwUNUibKYY4
FhFQdRUuIHbchHeAw4hvDKRiJc5DerKMuyMIxQrxt0EHAFZepDgumvmN6VAQA+0H1B2zrJ4YmXMj
tYEzUaN41GmaXlJuWc7J+3PB9jN6wFtREyyrr7xuyPwHZoElaEq+jb3IlQ2WBiP5uHpFuLjZJy8H
aeq+3Anho0hs+Bo0ivN4aqQAEGm4wWGTZamlQErd6Fxh8OaNkwvPL0FZcHAO2xOPsL4sG1kjS1Nc
1IpH5DtIbHuWbhHEvd9XU5VPYbTMgPhBukLavCGE9ksNtsXIIRckkNwVynKWU2eAb/P+ORgcaKPG
6mhYVEagzV3c5+YFggs8P7ymu+MxndRMgmv7vutbKHbHStL7SreE1abyCycHkxyrglYkSbY3b6xi
xeVpe5oCHan3qVo7LUFdJVEyoZEa+yu90DhRAiz11n20nxTZW206LDNT+lcHLeuqtaYfHS3OLZr/
Cv7DYjjCKQ9b2KcQCWHdcSd+SMyfmZDDgtoq5rEjciWt5NL1Te/Cl9ZKynJp2mEw9d9rKKKdoAZL
Z5ok3q+M5E2AXKeyBUQmi/ivcVnwokUKMWoIFLQKREz9AZtvz1hBWWeIq1cfKv2ORg78tcyGRk+J
29htYckau4A4QmbwCoS4HHYSX3s1cHGO6pvD0kFM8XwXGGfX3fG2T5XsPvfdi+lnJWMpNzQwn8XP
cDE2bCf6dUjivJWyfvQQz2cn09qigGQYBgOs0fKNz5gi8I8+nQfWCDL9iIwZy8IVow4WuRJ4g2zP
llRJwIafKnxBCVm+URnhqPQyLPtE4Bpga/lkjGX3n/etgAuoawxYRE5yH4wXfXrzTUOGX/kAGzaL
auCekM8EwGhjC8ziNmWj9IbkvM9uJ3lDk022+SWrQBX3R7TNBxZNrxz8dnBUKLDMyYrXnk8Y5l8q
WUptb2jKGP7n27Tz+Hmh9L3ypquj6sE2aDj+XqMSZGWlpSg2QMqIWVE1vi4kXu4pmwppScZ4L2SR
CbVkA650j7exlYVC8cKncCEEiHIBbI6Ja4byoN/fOxgCnaBLoPGp6ojQ92fGoaZ1CVF9Uh5fpRxq
3bFf3sjT7A9UTNVtAeYL3kDSNL4E19j7xY+K74U4Y4AaxYjCxryrP4H9PGmahY5YywpBuyu6z1tD
bI9LcIhI5nWAYOGMI7oSkidyZK9RojUpVLtB0pwDUt7PeAXzC+sHx3Hc9pOr7o/to6DTfIfXirSQ
aZVVu8tb2yHmS5IXygQNpsKpDMUrg9MW7wPr7JG/6hZ+1lNSjzsUvkvYrW153z/ExpF591EYJe7A
BaKhYxcMclCi9huV8309CKBmkfBgr1LKSUUqusn5sv+qnuVPyflX47z+dcocijRp884ktSp7yxaJ
AcnvMOGZuY2nMcFA90RBGPO5P5XrPrWkj/fDfnYKy346evIGFKVwcG0SeH0ISgkzXLPAeqO6QKZ2
YLg2o8ho4JfPG6NOOIe7S6NoRQEwKr0pT0JoMymEu/8ldpgobrEj9OegGsloTN5DL3vWEH1p+/yP
DkJzvtOnkU7jylF/Oc8pHWya9t7sp5PouhUmAIWv63djbc9rO53pJSjTLuiaPIN4usfjyTrDY66p
o+i+U05kgGLJMK8QB2aEfTwSgVpeBaG28hRCWAlg36YDkyq6hlKiGNoz1nZyQf3nfPluFrVCcX8k
jq6VDEdyIKqX3qhTU/vbkVXcITAubIn5WPXKRiShKObqAcSJfgVqeGQuFb4EU5LLOEpbvR3Di6lV
r7SXgJKbWsjxw0xffXiOlb1qNeKKZ4NQPViHji0VbVcDxuiKSjuf8U4p5iUKLEGnvRPZUJgQyCVj
7IBDPqg6Fih1QjEJ5oK61CYc0M1O57RrdAUZFkLPLbqofvbutVAkyMWyT8sywgMaZQMkGdTW8lE5
hwT/QIcYzEG+opmc4M72bhQNbBWLTotGrFtcitldRj7GLEON83gysyrR0Mlj1XkmnAOg6aiV8TAm
CAndGxKQDFlh/xT2N+Ooe5EA7+tywOX4ZjpbVP/YSKobyB1xjrY0xhuWNhkEJ3LY7wHIP0nwquZQ
5F2GgPO3e87AHv8m6sKMjLgBQ5Wn0M5asFPLd1zd3SsWKkJUwl9SQKaO7Ia3BcBq48ctT99OJjKR
PNNw/BK+Gye7lrCoY3KsHbG9ck84+uVUb5kKg7n0wUWjsZr2uuVUy2bg8EVmdnlwpZSejvH3Mzxs
l92j36BPuup2d7S3uGYSVmI4zajOeU0nNQ0uBShPDyJ6gjHFXn4fq3/nZSjUOoBL7RH68YKdFlPQ
PcFRvw4oDD/PCOJoh56pxGpHrFopGvET10PjxitdXR1UV014LMtANbQrssdarIq5lyGuDrHCbLjl
knjLGyGQH7RMHg/45QBcLnTNHhTc5L010CfF9v8VGii5CO9VFydIP1ELnqJL4QKrc0Xhp1KYkaLh
Z9z39i9cBfaflsRGspFv3fCaFQ2qWUlDjOuCviBUzX1kkZWHdCHHeUMzZEksTN6qU56W4XdMaahn
XJ2eILolRrf3Tw+eMUYw57jEz9eEZHfhFkyNau+RuRuv/C6vdWZ5RILOLn6l16CA4WV1MCRchUbF
cHxJ0JVHF4xFfxbxlgjKZ0WtJB0rXN5iaBJUe4nBhlbX44mrG6mRwcib6XkWSc9mlj+pY+p6vajS
53UETZXX3UrpaNrxrgGiUerSnNIK1fGxnfAaOAOd+z+MgSr3DAXb2q9M7NFfnMFF4gIT50FgmYr7
TuDyu795g3LJPWCMO1rLHDbH3RFYENt/P3g5Ur0QGajJLErmuS8/VaHlBi9TMUNYGg4W7sVi9BHS
mmjmbp7KNriBaH6IrWEY3pOv/TWUJhG5r3GFet05vzrF9NWuV2BuUoaTegteOF0Fkt96L7KtomOg
a7TWbJR/cxS6+cWZ+JqA+tr2tzKpCWBDIVAg/qKnof2+I829p/BC/S9j1WfWNcFoI/xbi5/hBAaJ
wA0cd+UmulGCEyPL1w3PvvfVueLtAKt6fyJ5i4bzZntOPVBS/1h34CuWEfxgNRu3e0cb8vnNVLGq
RGHWvkUC0ZWuGuRC2/uHu+Y7ASIOmcbKw+6FTp8mCLGANE03zLbjHTRCCBER9KeyghtfTBOn9N2E
E10moX/JHb427NWgetN5GF6HwySYY9RHmVdTqikIeGunNyQ4PWbXI1BjMT51otcsZhEWgjvtRMFU
dIswWkSshWsaQZVmJ92JEZbS+wyRD81H09QHI9lUtZCGM3LPhDyW0NoSaHaQUNxLeM/I9QHFOy7o
k3twBXujCxrzTzg4kMLGj/EhDUwAP4slvYZBddYSq8jZlh3AY5bPdaQLNuF6BP6nQoFTzfGJGdzf
Nd2iyXvn6RAWmA0O2CaOyd0DaK66iqMzv/4p5Ig9B18gPY4AmZhDE1fS3Gva3JExV6U4Bk/g/mUg
wWAzRFd6/n+KKH3fVUyUYE6OtMk6fi3uZZ8+9xJjhRLYbVGUhn9tHLRJz47s/A0eZEtMuTmy4iXu
F9nL4gfsZqAYGa1Gd2nRgg6+Lg4vN+erH/6r5GHJYUCIhL6a7nT2d7aKXpo4YI/GPKjnzbdEP5lF
q5A677UZXwNQTCqQzPBvwcm43xSvgX3gzSYaK5k2LKm/6Z3B4qXhzO6Nj5BVlVgC/8DqlM+CbLen
E6Y+rxRp8wdf+L8/owwOhv8rnw5rMnQ5yQIYiXOwyPEiPl8risk8lx1pNkWSdycXr+c3Pche+Pgt
vii6HnHt4tJzwXiZ95zV6DMIkslnODhdVmDHTU5ZrYLkA0jI111VO1CFu+To672DCjuvLHMfKI4b
QJuWLtelP98w+go+8qK34BPWHuIezoHMImgU9q5MA0p4xK/lmDO6NBOh2/wEhmzaU7hloNzVg6a6
DY+lvn7tmvHFRtnvyc4daZXweKQ1kKqlVrnM+SCSP2AXSg1ZK1MX9dUqztR2fzQuQ5llj0jokqQz
siOn/NpVC5DnulXuIgJctKlbn2cR+e2CInSv1FIZ5T2LNbRIGCuWyJExYHacQey3cOy3sEgyUgBj
1OhWq15vHvmFyK48bfDrn1PKoUcE0EmThiak1IBtl53LbAZIfZc5St6t7Uf05CCvUC67kKHAvMDZ
dq3fzaeumGHnKJSaO4iJIBbT3JPinh1bCCNLurTul5TvjepSb2SjD3JksQayYBc/4CYuBqJhbDPT
Qdn6xRJ6xfTP74yPIrb4nY8ARYHj4F1TUhF9zrpQaubvpCPSrFlmjaF+nhQZxs2PepuWU5nD7Eot
N0r4fClRryxznVyu6bcejfztRLMOtVRIo6fJGig62d3sqvfJEvbFNe/w8S2qNP6nl11KKjQzSHTX
VF5rqQurp9oYO33em/TbfiLbRNz/TJ4pPGQVs7siEeotDLbKCkL2ftskkuJTr4rVsZE+9NJrqUPu
KVwkrqOqkxPKrUmPAO2RgZg/Squ3YpWlVxZ7yDEDxCfkFIhWYzxfTdU7Tg61clt/a/Z1IDbk6WFR
Kbx63waNNBWnRv+4DopfMthQavBbNLPq9/ArLa1kseYIjlIkyXS+OV5qS6eOYoOh6OxjfJT+vz9s
pZd5mnINeN2UbBo1noUxcNNDa4UvhfIBSA7dJmivJtH0avD7ga5rfzuoIgwDkjAaPpNJA8DK2IBK
xcnwrKm6PJbwBqWFIP0BQyNdFMciNnFq8w2RsW0ZO7Tb7sspxXORB7GVWE2c/mUQ7mW7PBeRD46L
yt5U3iAf3hiM7O4O3rR2K9LQShV4QyMh/ZGxg63atWqPRTXLMJuoKyWfA3rBZ9qjYo9HFJDYuHOw
R+zGXOKYIijfchJ67ZSJzmZMQmSMzQo3G38fiSlxSmZH3PdKD63JvNBpaG/waCSvXHg8mV2xG+Ni
0XlVx2gbhBSTg5/Vd2qzTBwUPi4MiLakeD/7M6Kl54r0NLbGKkeYKFLkn1cv2CAqFWnB0timD93D
qlO8a6yZLatmIyAmF/YoBorsIP96Md34N+hKogCpE/9kFF7Tf6Y34GbscOeuRKY3HVwZDGTcZ5Jd
Ri9gt96cbjfhqOO2vdRxobxhJhked5lZx21QxEYpBhzpdOpYYZEtjAz/5+aGb6KBzXeCF4Phu4W/
Bt+jUt+EhcHN9XFhoMmbq+WLt7q/IYL0WaEsXbGo5saVVnELCi+jHjOLjzPt0xYqZIF7KTfIWDhn
4UNPyLKA2de7tvvma0sr18xbkBmrlZU2k9Gy7LfzAbt2Va9A6GfdKOO2M+SHtyywZl1KwY/UBCrq
MndBorV8K/r/Qo+R+tyiSSnNbt0iWRVdBKsjL7EOG1/W9b5IpZum5R6IwzaR2ie2IF6eqh5+WBPs
LLOS+0iol96tjUtM6oh70dBRyYDCrJ9ZaoJWxJopMIkSoq4IZq8f/bOEy+Ari9S4pw3oV2sb/niX
9WCgkgQZgSyX8Y95pYlDVmVql/RM7t6nGTFyi7Bf35WKQH9Ltmea32kMkIUehZRfMqfxUC5hLOtk
eXzBDihjEMctRO88cYSZ+vlec6HUwJUZucn9V/IR7rk1htf5td69xvze3l3fQbcSpHmlqN2k0ZPm
ILO5fgBGtzEiLI+im7lw/H4aCs7/X3o8b/OpD2RSTmI+tU0RBek2YktCVaT9L12huExw/QPZveid
mt4bVNClKZDZLCLhUk28GHBxiqA8vT/EQWaSOnb8AztMROTg97t0/RdBDE13U31Jo9cAXN5KGMYC
QAKBBGvHS6MbhaHKEuAM8doOGy9UMbgfpAEgqmAHc6esUbX+Yba6AwTyxDrdU8lYOm4kcC/dojzL
qDIc18E/V/6sK8DLlD0UOZ25khq70eYxTHJxQ96yaC0+YJPZUvLlywmG5w0wYShw8KK3y4ebQl1V
r8ZKJSE4Xpbq3Arqxfw2//QK4yP/tqHJgebB1eq0i3SleKpcmsorzkW1LLviJP6tXvN3JDT59Jye
6GoYJNifBfrBl0WrBPhOwTFWBybknRsWdIsIvpaMxXypGGifwwlEEtZ7xhvk7h2D3A6r8tpJlD7V
d+yAv8bib3TuIlAPjONrw7X6Wh4EQzP17uBAO8oSlP1ZPF31nPeMPwOYCL0FeiwMtjIJH+4Z22ai
Wj/EQSRe2bU9vKSepSJYxxhpoZ+ppHpHXOr+BpQl17TOnbL4S8jEZS1pdRQttn4rOibUJLF0oXen
TZ6cJb/ePAP8ixR0iGYVh7n1WH/chQ+Y81M1a+Ac1a6tUhP2FXra1reVyFCFZWoDTUVa1+untfyi
AmRrIMNpfm5dfJ6DyVVhBrQFwPZQeZsPMcjCrjQqzl5EOyrSornVI/5BbtH8VyRBx1CjSmdCjzq6
+FKRPg07MvWtDLEdbWywZFChwj+Y4Ke/X3s64gUCrNtsxauqhFmlubttWEVJKbejBC4nLIdPBTfP
2XYfXEHJ8nPpN9IG5tRLWBWXyXlE1slKIjlmFLmUOQyrt+/r7zogRbRLvcl1Rf+SxN64rFX4MFmf
5IHl1mYluGd3Mi6rpq9AcYfEEXr/QNnXxdB/yThKgEX+QUoPWCOd2lce3R/bq4X6VvYup+kMDy4a
gp9H1tCzi3B7EhDhHwKNVCp9PUln4m9fkGKubXJim6k4DkHAVVEhXkTP61ORxOPsSUDGRnrTsUx2
NlJ/6WkIxxSGds5oWkRgnEXSxYqxy9fhvIQmRyH4KiFFDo1RmVoiTTdLMuZdevlkZl8zgzZwKNnN
WIPc3SL2ilrPm6cu+IgBJFKaUhdQcDr7CJkmXuqnffEwgWSBoF3rGSIiXrJT3ZPxJuU/0tnQ0j6D
tzaOCCnvt+sJAivBaeYvxTmcG91SEGQMxZ+DRl4xTLc3WFKZ97XISVao5DwBKqLsPWeOu0gJUCPd
TuPPrJFHOiUSrrYeua3K7dGVK7thV26D3VUIdLRXs9KMtDAM8ql9IuIH904U7uTmexEw7JbbKC+y
Lo7+lZvOBM5YIF6apMZoH5sWD60vdVRTUR1pGcUOquMElGIlfrpyW2cgLb0sil5iPjoEonRFvgqz
AmYZDkA8iO0XXm8GMp1DhT6Nj14DBaknf7gwcPJ3OiQVNWg3CmJMqLbcTbBje3TutekAzG7wtSBp
c69btqFV7VA60+aSL05KonDbVpNSYxqXuXpCAbnIbYZoI0DBRMb/5UdYjF35k20vt5P6+P33AhUT
6mrQMz+i8ybjsOZFXuJxHtaWmu2c+8JV5BPX1/8LqFHQbN+SjhF3XR4rgK7d54uoCzZsf3vw+PAG
0tUGiURof6dUtZwczj4ApYOStZf3iZDlUPXhZE6aUOm23iQN4q+y4mkmW3zxwxvP6ICVkh9qOm/q
IS4fTQkZG2v6EIRWG9Jbr3Qtt61+mFbLRL45ClK8RsQHgUWUZ9dwoHySmVwgYPuw7RYTfIFREAJD
1X8eIrGet72hxKc0j+AECJKJa5K/oV2d1O9CuiTdds13PBpw3nJVLbNXcpIhNK9zls5w5RrwUvGd
QvI149ayUf1Y9uUTqNLFEo3jkbIKdbzeRSs27Bb4c6Mjla3TU7gA1sfWSGB8yMyPmeNIBetLQAzk
mv3KWd/awm5XhXScZWdAoYzqj4H5s+JSfxr2+EH+w4gNaFz7RwVKz0xRKjnX6ID2lk23UXS5V00G
9LFVduzXEaRG6TQHNQe8nk8FPZuU8Bktivh7Q4bJ8EoIopAL6jvGI0mIVgTlPOBsYui2AhWj+B7+
9dJGjak6+flG1XFpJGJliYF6bmCgAXs4BUXTBE1LCiL3dewXI5igrw2gRCBd/pXEKfyS46sm2d9I
id3t0KgzV4R1jKS8hV4cV070cNYhNF+Trhk1dWEzDqBuU44tpd0O4/c6EYswTOxC6cCWuDrgbkxP
O3qXGio813aQeMcxEI4hZpfsFv2BODP3ls5ql6yfgE3C1h9ooTD6hsvhgX8/ygMTb4uIwn9MEs45
NcTaQ360Or4bMcSl6My7x0e6TWNHsU1CQZrubFic0pguaW/0gtY8Tf09hhh3uSEmA3YD8KWTkXwK
1AgBagMoZQeyOMpgSeQzcuMzDiNMk5nZmfAFDj674pPTaSfZO43047HOTn9ppBDI7Egewd2X90Wn
HqGiKiHQij9ycsU5v/lqAkE/y9IBwtb73Lf8A2/U4qIfrn057VsHISKzQo0CYRErkHls0/V+zR4g
pbl4mL7xlCawJEnvCZTzw7dEYTiUAIclTFWjuBJFfU2MUWsTvJTfTRDCrvrf3VTQ4NS69Jp4orMa
UZEacXEjAxqEPMg7sEyRyBk5pcqq6rHGM1I7jXUn5vHvIiPikR34JqvlJtoiBTOzAyJBaRe5waWY
kL1CGRuSmeUIDaW4MgWDKYBccQqIuLysAXANdH5KOSefjE6XOHjplGRamNZubESLwky+Nu3woGtM
16jWUFSwUjj9tGCC8mVJNe+Scvx+O9z+X2L/jkkH7tjxS+OQN6ZkOVSqD0YM3pLr9SVr1n3US3hg
xLMaAU9lcsjWmLFP6wdfgQ29WAyy1xw/sCBsVi4iyn5MWLUjP+UZVG2SyTsrERtNlOySe0+TIXWp
pWuZB1UuKK2znA/Ac3tNML/9YahnZNYjePllJnnbtKiQB/3mPO3zuhwcoB1ltCfAxuCRCjrn7EbT
09n8DqyIffSxk37K85sqYwDEkcg9nonvyRBiSdsNKx9jabZ0zuLBjj8FFCQiokc8CCXdQfDyyNe6
QhyMsNeJJoQfH5+PkkyJ+vNIoi/dvV6f5YN29AUoWt0hlvKYgtvMyiWtA4DM9OC3QytVxgb7TruQ
9W5Xf3KRQQ4xILQGEgTbnqZSzhg6FQuakx2n7dq2Y+TI8YzNaPF/bGKmlD347prqaqW1j2qp+l4B
jvh5gDc+XLFexMGHkJJ8AQtGcmWieSw80Ezg5fktTSxl7a8C4eEzmjP1GqFTp99wWfBYP+sr/5rU
A7vXJC22dZAVDHwpupHrr5WCpgDusTX+ccpg5gP8E21CbrBUtu2e5pYOcf39JG8d2wv10CSWyo4Q
IE08clrPeqaB++Rq9Q3vCFxFjJOPAdPbNbehtaZ8BqQf8rS2yvsmk44tqzlF3gh9wH8yGCGIl+9L
+TA18kg/vuvpQbYHkKoCzMRQggYSoE/R3cFmImHO5GDTszgEvxXgOqyjNEOR+id/Skqh8xCigVXx
eVvfUQLvQKvaWaKQJd3e0KwBhpklt7UGKptDR8EwNXbE/0NjP6oeOp5qeeUTAyrgyS8vHfdTylXR
BLy3MK4Bc4UjQwBJLlrEOyQiRujL8EywCELSWp11HUmDvXRN/mnZ7RphOY3WHPYRlnAoI0cCg1hN
zOt2n5Yq+VGYf5ZAINvhzqn+pHGSOUivFzspOd8fZlRV0qexOg7bfys1qfzROs5v03IhFyTS5eaM
SEsoaxaG4niu9qeO/+hORd+voZl1Z1HNPNUCxB/kvt2lIXF3TTCPeo3VeG+k8FHzCTaVha3llmTV
FwUNC/9cCkam4q3lYmml56IWM5sboj2KOZY/AWxQwJuTk+96fKyTNMVP/6TNkLUkjxraVQI1RgCO
vJDInvSBm+f2zSNMn/BiKRDcINlCEKpWn/9ny9cujjDpJE4MMheYm1nrXoYM22T4RkcgSqIgDYNK
WopEWtwDiVrYFdBKQM6WErhvHQXn1AKi4HcAWmrlNMnM71iPi3UKBcTol2JwkEUdxYSj8PaeanmW
R4ojCmafpBcxtk5k1U2WwhnOUvjmR2a5c5ngXCbrDLyfE+1GrU0nwf3Xfplfyro+KbJuszGpdgy/
JNNThyD29SHSDWnu34jKHv+pDb1Vj5S6BVbS2WKOLuZrtCQql0Z+XmxskMDOkdheF0OGyg7mpG1P
8O55I5jNU5LYJo2q0vQ+Kf5GdHRiyfYLWprrml6Co+Oe7nu7aJA8sNkzUkgyZ6nycuMhC1gWlStN
1e+7DJpW7X/BEK9qykA5UPvuRoeExHKIJ7vNjUcSN5wIB2L5E8E3EV9Ynv4g9mN9D/YVuc//8hVz
yDP6FP+VpKPgxo/cOqiqNtaOxBqiAmgSm+8OCTqmXxiWBrGPseVpYKi5yPiOFyO+0xmkv05Y6yqQ
MncFf7BXcbsKtuDM5vz1Q15/GzIzWeNC1L9SX9HEksJJNkqoyz6HrevEDsk6AZ1HuU5Sz9eisFA+
772SrEzskOzHDFO+DV8paR9FnUIeMZ9oZot/YQ0PTdcnk1vIJRWnw/2EGOm/Jlh+Xp2qiw4IjM2f
uMtYmkfDZv8TNe9y5KdOmdoo7dExNwY4N4wj3sHaNswHT6+4ATTI5nVq/AkTq1OF4hxUWP3V86WH
MDnOitIiMqI6qsIBZFNX0hizDEdJZii1NMmdfOHjupzJ/e9xc2frcMTWQU16RcxKKey7ie9LFf19
6FvvYNUA4U3tM8mKt7/roLHIPPEddcIU0j5Y8dpC8NYOhAYkWRCAjdeFxxN/z9AhYi5/yEt1vaMg
bVIcOsq8GXhp37ZwaSXcPN99YpE/0EpM38YXHUwSxh85lym+6Pzy728bQ6OyWFLnmB1TlrlnDM8W
4a7ZRBdxzqNIqdQcKUD71ZvvNL+o6FCmKUo4ponxbgfW1DCFmr/j1ZAopBxMJ3ljYR5aEUfhJata
gfd33XPWsQvE3m4kciIVq3ehWBBbjBCc90dYWBFGU5nKAM3Mh8Z2xQhBzl9IQqx8HS//Qhg8GKMM
yHYJhZyTZXmYZgUEbm71rvDXJf/MkoxIdgsL/I83Au8AiLIuONNHTDCZ441P7qOaNvbYc1en9iPf
6sRXgLWfdGrxGFFlCIoq9lKmOKlBx+SFGRq23Hivsaks82NrcpyVAWQ4zCwz3FzndfoVStC9EhBO
8iiXmpVw0EA8PuHq7qzRQovC4egB/QZAvqQirzeSigI+7hSy2Fs8sw0cJ9YUPUa9kOFmGwkBXp20
HqggwlxIXsm7EiXZn3kcEtl20gp4X8/kPcLqzOUw/WFe2IyuO0nfRSaUcs3spG7w5p+6NDShoMmi
5hkyv+UyWTgKXt/M8Fpje5ltyiKCTT+cdqr7wDqptvjD0P9hXF717UhN8mpDNhkaZ+eGFui8ezc7
55Hy/bat6AELzA62RZJVfC37U+kKN8G8rZWYl9aVmbiHfJrQoBUW4SlHIk8uboxsouAQPU380hdC
vUpE7zBE+plS23V/ekRt1R+wIDGqrbp51R6LoTGZncoS5TgyKSlrV1oDaBzAVZpjs3wozHoMV1dW
IRsTyNvhg+d/BKcp/AoXBNbRDrH61/yXaD/Pvqy1DwsmbJr15aETtNKUBStpGfztbqhDfsJcd5xn
tzuVT/GEDGLlfOPaUp6FxBXoabAPfsJjXRw8o7hEpTj3kAzSOud2qT53LlzrvXY3O8G9A7mUxH9f
kv3ih17UNgF9FqBwGR7UBkChhXqpCRSgLcrDoL0GqdzrCfw1shnzD3JwdczW2DtRgFMAnEnklDir
71DGV1r6kpHuiEImyVsaRtkFGOU76lTyWlQB+d3AkHwydZO0zfbEK5P5mp59+FDg5TdQYNp84Ok6
e2YQqj7zDR4ycZhy93/TE5tfHNDufjNRUdW9lB0ZQgMZtGAVjzhs6M923DJk8AocOn6uD2vSrO1M
OjKj2tX5PtH2zTIOFP67mOIH3GwdDVccnTtXQZV/rnoV0CHPBqz/RbK20x/u4zFJlmzGkktMsrnS
WvoTb0EZQZxkFnEm+uNr8yLQ8tjbIdQ9PSt9v1EAdF1cTKhoJAjFDvOO6/ab7fadneu5pCc1DQ8e
L0XLfCJQBamcaN9/1aysA3anQk/hcCU/S2sASTWw57WCgJyxt+vh/is2U2Mmlp0EjkbuQBjKfcxf
7X1t8tktWAkwN6ezkAbXPr6ThFF7FR0aSPayY/8JsH14vuZmZL4VUmxHTapa6tqOo2JoUPVqfDCf
UrWn+5UfhVVwNUrprGP6UIBGKKjxMZzq8Ndwb65QJs6nctJfw+1MGsMDjV9Xu15KayA5R2UC/7Mh
AgtQS13ctD3O9H5MxLrJfU5hIccga5xwl2e93ZS+yDUNpeXYrH9/LYHUAMDiz7J/nge+R1P659nD
q/X2w8ixpWGC9m0Y/dnuMi5Q7nMX1H4+Wul0Gd+XVTfWx9ieH7sagpHo4mxdNea4Ma4zxNnrHb/h
axN0fXAvnAd6DK8adCyvUw8ii3XM00C/pawMCjtnNB0JAjJdPJmhhAB9YlZVlJCPF9nBMvbof641
ThGLAHv17di+uoy2SQyAaEvBJK7G3/xRMrLCcyMj/HL5W8LLbuBBCr8NzE0ymz3Zwv12t4mnp1/A
2uK4AOBdzvVE8QxrLD7fqWZGauG8wt3OUFb8AVBCfXM1p9RBAL3UWtVCUa//sYwaQ2Pjj2DdVOTu
n+MD2NZ2nezywbEfjCMGum+L+jBarL4IqqWxKHM1TNM9NA2JXg0v0QhaUWk6wgVlpx6KUh/Fxs/V
EUe1Ny8PZ0+o4zOYysd1SeGVrAWMhlP3l5D0xKTHaNBxbS7BHiTNI3aZj9nR5pZNLZt9oyBzMJfr
8deyUWDpD1wrWWZ9bztL7pB+Zduw5HdHycVdsXedAdUcRthU39qXNS5i0NpKDmlGazZDRYn4AqCs
jQzdHkXH5gBifpOeBb1EYXq5TOOdnDlR/nNr5amM8ITVJ8FghXhWe66rLg7/kfFJVZbXBa7osbb4
tjJgQCVAMHRmHCxYlzDJcKmYHVz4rEo9VgkKhh2dBI5KTF/gOwytclQc5WM60ogTX22ROOGFtIav
lP7ev098fpQygGkS+FcAWEG1rvs6LruBKdC3XXLP6q8RWKpxl0r2k1/VTdxfSVmZfQ4/BtQnO31j
JJxv7vwd0P4k91y3KZWVlMwBOjtE7P5ohZJDLx6XdtsS6LVk+uv+mxhdtnN3Ou9aY7Rb6brOQG0s
fY1gHfDU0YR+g6/9JNmdBvEkQFlu7Z+VOJopRTCCEyV02xLJmZqTPwKeyblTRXMafQ5laRzkAMTh
AI9ccvucU4RrdDKbtxBDUmQ+wgs0wtodgEHb3BDybV9sjm6Yjio9GOYJQ5ywJkfuPvTXXRcD3MTm
pDtw7WJnNynpL7Il5ry0iLamZnf2o4qKRByzjVB1r37I4OUzwDS5+yzuyFs0wQXgEf9Z5Ctt4LNB
A2CHDCfWCC0qRmoBPqwNZYlosq1tJG6J7ztE63nt4Sil7IWjwlvoKdoMFFfhGMb0Tz+J7Ly6wRkU
hliqWnqVO5kT8KbORZsI+r2ceDdYVoU0n96Po8O6+uq9b0r+KzzVRITKv70xpjAAwrqrjDhzm8Bl
k54g58yra0lkMKqdcQUd2zQrSDYi5wQoJG7Sg3zfWbEWPNLObwnnZX5zSjyH3D5tVY9apBAJRU4v
6sgMcEp53K69UzVIPPrV3ht2EBIjRkk/hNbjEG0cYuk7Zpjh2E47hOptU4p0E7dMmlmrw+qATTxI
FZihvjKD3ZIX7Bsv0tphXj8v2buT0oAhF03PzfTFj9c6OrWg9ZBBAo2yvwBkGBKZOFqZkoxcZsCw
hi4creyHoKAXziWYGBp2VUTONwuMO6AFVDdf/1a5QgX4a4NPpMyOqXbCHcfeDC2soigjrq45/0/4
TjOzxp6CvebeJN2RGivImbpqNCC9/2NobCYqxj6tMBRLOYG7wp7CA1hPMWNbR5W9kdpMfI6knJ//
V3dQuvnDIcJcO0eUlmcxKh+iivATP7vE618YUxR9pjhf0SQbZuO6D6qFb/MIOcVQGLMla+bJrowG
Ddja8clFXHFgGaqrNXN7yQ6Zit66hffFAgwLUM3V9b01zDpdQ1ELMpuDc5Ofw+ah0h+ywDgbSbf6
Zx+qC9nDT0TQOXr0vhkLd6s4LDxT/RPNeFJbO3/kqkYI5Vw97xoQc5N+4A5d68QH7SR0q/yaF/kE
RRnAc1bC0Fw7WTA6XwMvReUPgAqKtUrPbVy7iFUHPx/qzAinvr4fM1T3g1JT/qSnibZR8x+24LfP
ohCFV15Y27SKl/kofTxpKYJjc0ZDX8d4w+b+BcQKasHm5RAgUAziyiPg+7ltVOSKcfo+UEMbdKT4
k0N6jniftm/V/1P4mbEvci6/AyMQa8tOjQ+vwX/dRUETNmsw00jVPFB3XtEBnVFbLvGOyWoc3GAE
82CCMD89gGJGWL6yBqTrjqs0hAH2opnMFr8fbs0dgTiLgd7WGlilFmnOQI+XPRNPW0P0BDlP1TTc
TxpyUZUq6eMDLngg/E8nl58Ai5qLYVXCc2CW0WFH28f/N8Z09KRBBqO0IPBV0/kH3g3o+BMiiWdz
4fbMCT5MRXy67dzGMcMsnJK0wQoczZfzFK/ontTLFvvtRgQ+VUP8vwSSmh/O2baTVQAuZZCtTW56
5kwxcNT5/OHc/iF2AReDHdNJ6AzeAVlJthcc0bKbZXBjJkECkZSCty0mHeP3b7FaT5zQMTPGsLO6
s3inHhy6gwle6PLWhaY0Oos/+LCNsxs/WY6UPNix0ZR1SjbUL45e1UWe6gJtoBJwH5UXFVDRhx9Y
abKOVyu1Bq64L1guXl++ZkLXnhB7AeHJlBTit/kxmvIgSdxb4W7VlpuKBMAqIYieFvWu8T1rcfXX
gW4zZzUQqtSosWedzkrftVAcHQQ7F8swgXIBiO4NiwcdVs0IolXoplsroHlqgBRwyYRg58S7x7Gb
kRpvoe3MCw3IrDRfJMM4NZ0C15WTVUYo4eQgW92iMpemtGiZYmrs2y71ULd1sBucLOS8H0xLabOm
uWdi4ox68vd02vpzVnK6zwwKHno7xjwCA6alPcABQxhYlOUAmulbvezTPA4dRsyingq7HveYVJvu
lE6FNDDIufDjq35XBIKBS0CVho25SCP+mYWwBlgB2pDM/eX5nJxrWavMaFJB1czrB/aKVV3HOLMS
NjSV1c0JBckkFwviXclyxN/ZeTFgKBOAMCTsC6D7pdPtYlTyKleGZygCvNIe07m0cyWztPY4sKoP
nuqDFWsmlrP0zbV7dONaTHoqip2AAw4pAYoCvypFODdLHUEWRhNiYvC8aQwIVi6UNqkUJmjHy3nA
eOuhPb/WzZfu/MVqpM0S7KfnKUA+IrK9KBmy+CzLQ6DvdGzMeVBVS2m6LEh8KJK58Gjc0Ek/lg5G
L6ywTcTyPMGUtfLdFSk8+oAkN+ut+vxpeBqXZavNc+gtHGeWgXuALenYNC7CLP9cFvshJtQoUAJN
pj0/CBXXIsezKRk6PkuapoyULa68w3IhBn2WTS8DAhNohhE1ky4A7qizQsotTAA1GbK/W16R/QUH
hmOqRXjv2fKsRItNSCzII+6CkrZiuyZs7dxJIBejN9Qfg3HL1Odwq/v5dyvzk2snte12w9QctAYx
+9y+0hOpKJHVF1oMYFwV6BTszYgOggLSR7sY/5AY48tCPSMRgRL7QCvQKVXbObKlkRJoV6azF7Th
qxjCF752uND8SinjiDFGS0bhm+vj9qx/oiuWOlLOCo1+3HQFM9BLpyX6tDULvn4a9TShco2+hyST
y/XwR3OfwKR8Bz6AHPx0d70ERHD6Ph2wx4dclMdPbt2/xhyMUIy16r919Mx8vtSVEUeSqb0hv5RC
bU9Cpf5rD9Sr3y8qG8C6UUUdswMl80RKHGcIFFRud7QYFxnWjsPjxaY2+PlfpSISjbsHBwD+pAo7
qaiP2+FvzxAOkBi6O3cqhlLQCucuiZ7ucdadVtJ9VDCNd41ls4NBA7uRPT6VuU0C1ivtgTUCKbe8
TI3nNHEGOYcnKGZnP7GrPQfwgweKwSjX1DzL95IWS+2BIXdph3Nf4CORfe7zcjpPHOHEiu8umbed
9d8OFCVb6mFC9zifdjc5rf5i4lwZ5g8K/FJIHtjuu3N/j9gA1ZDBSJTLssSfJC1/fj8TXR7LeJT3
UiIuJFaXR+mebV1bGC2zRFKaiOIm5IJPV0WQxiToYRrLJ+RRPyQ19lFloTdcVL3qDIH/1ffMUU4Z
DW7gk1U7hI23COYPIlNnO8kIjMuJFOPKb4u5JUgJpt3Ctc89dZzVDtFvHz3VfZmW2J0UA/zujA+A
oBaQ3wh+UuODpG1+kCCtcD1LZbynEZUGspmRJyu1zZe2J8IwVaQXWCgtQ8u4kKtp7d9R3zhdUUEe
CzRYfqeBLmA1iDgeJLCC8JGRry8G4FBvdpd2dwON+R70BfewC6Sofk1qrqBF//0ojtKYd0M3b7Ni
XnRzQ3wJPqiDaLlZ2jNhF3ZQpRLUm0GUsnH3j00qh3bbId3UafSGnV3SXIr8KS7iDnpaC1vthx3w
Rv5WNJ8f3g+jDsGwiCZTaIezgTWrFY3OM+fbn3in+vcfXX2wGjU+scbbPO45/SctbRsSqy0W5XtR
TAMx6vgGjypvyw+hiPodVdZI2fE0eeaoyygk55kFcN7gpnxZk3UoaCqoakhLPUIJJH/mtBDRLRPP
0IO6YyWOmX/DWMl5sBZl0cph2bBg1J7Wffi73hrM66JV2wzhKt4qiEphggaKChTbuDG6LV5fuMc9
CVxWAkxi01Jos3//Pgr1KXsp2niK67xrhnqQOWlt0QizK9zHblxlYxXdLnUkV6SOLOAISe50Otex
WEJRvXq0zGpDXNXnlJbBBsqAzAiYO6wrZICr0qQTyZKUYal5we7lGB4mPQfNA3cYf4+CMBFAuE4r
VXHsorWyPvEK9d5yi+KXTOG5wh3TrpAg34lSaMqgnzSwf/vjb+4EgH/Ldmb5iEcWOP/LKR6gMaI+
E0UiSGKxEANbOa6Tk3Onvuv79vA8GcXNTjpFCSarI6jbVN+M9KynZpUxl3BQPWiU0p+6iWh2EdS5
DyoYe0Fzc9R7Ixf5u8/hG/tMYulexNlkUVHKEtxmXnMkwZ3A6hGodHs88Zfia1SQbRarcyWaSh5V
UwdgNXwW+scky1fBBlu1YC96F574HUox2MrxrgDppmXObpooyNsKGk2unp5oh8r4jJ81CV91lqDF
4rFtrWBjoli7mRj03nmzambkeJNk8GgbYOTV3ujNk2iHHs5pbYHay+BR8eCcxHsbBL7O7yK7pSP4
+wn1uqTt6JviTdQyToEz52pnQkzNV/cZp+lLY0YFiZAaMNm34CqJYCW5xHTvTDSVxnYQ3XjVOgf6
qGS2g0jIbdvbOwtCrTVn30LTPbkDLPQMXhZ6DdBvO2ZOJmLi+sBe18w6r1f4/oezkB/wsRnGeCVd
BWHP6hQcCuPyi36VTZR2B3/LJqUzlG2tNcRb8HVHdwE3LyLhTI7TZAl2dmDHe/atmRFcpKij34Fj
LyVXXp/4wLI7M0Os5Td+7+h/NymFZpjWhcj6g+S9bxIWao5PyM61Y2ao/qxtYtg/sAX/clLl7yaZ
uSqSoW+P7/A4wVj5aofLKbuh+/9fM3w2Gq5dkDi3ynPlLvlHMq8idOEajygYUj5ibviTRKEbYfee
aiXhNH6hsExKutEXxpBJpZxnc870LgzxOBYm9fy+hX988EpGaJBsmPzgnyBGPv+Eq5iVlKJqEMlb
uOyqwoaN8AYYQ1sUDXF6vQ91CeHmGOJr3giL379wWaC0tVYgsql112q4B34meSjdVtI+TGEv3NBe
CSQEf6ORvqOOVwSvvsqqxR5j1yNKLzVGuzH5ZvD2vXj0Y1rwWNlMTWGNY4Ddz++J4QVY1xLL3hOd
4YEYQEUTA10VR68E8ZS0a6pwOvUe3j6Zr8+2PRUOaekOG0F0Tt0JALPGQs1P84Z0n7km+sVq/fIg
pTp+TCfKgmjd1CZTr1yLLb4E+NWx75FYFkB0WLIHAt7IIVQSyN8VcsQK2Xk9Ymnv36rvELaI1DUO
A8igKsJCjlqT+T2rkmhGKZJtc+e4arUO5zGnSAQnvZgX3TCZgDHg3gto+Obw2AQncYeEs9wlNwWD
9fovJLPOZ7bsYekZlvV2i0t2QI65X8xOiU5HraPNmCTwo6RznSRZ3tc6feHPoR/cFQHgqBEsKIt2
MX3b9nY6dWnhUABYLcE6dabyAysOMteGq3HapFdmuHE1V1HovnsKUHmIh8ik0iZqdtRG8iDThOWB
d/+tggLNBKWrVgk98SSaq15XYVUhlppzOK+mJtovbtO8Edh7jxfgQ7CTZ3TvUObHozefCjvEYftJ
Eaj5zKGFBj4GQJfGq40jkBr25jEii6Bd30WjdmsvjXsR6x07AI/jJ+3MVIKqvfns1GNg1HtQlei/
PT++gtzp/Z3kMCidC5iTHU+blA5e5j2JhfMPCcfPF27T2e0A5JycPFNwNVcvSyz4uShjQuGnPRG9
irm36qQHgDWwFlP8FZLDQG9an9elGUf1AAXTCr81/MvqMfdSQB+tI7MgvOP+8RkRbHwl/Bq3QG0K
MBFbN0PNfJEOcajznBptLcm8QKdthaaheaHkJesIH1LpvVCo/4nWjNn9Y9LSiFC608gQfJCXEWYI
YOISTeO1gqTwJW8bqLcEHBzoDit+8SKW1NY+MSD27nnSF7/vBP8KyVWEStefrJm4hvdk4jluViF/
RbTXjE/9DvcjIUFVJdE8qOUiDnemoq4s8Oa6Fw4L4tm2AYN5xldl7XbG+rtJ5qxZjktlJqLsWabJ
WRIAIdtdy9GIVbjSHdz9mIMxRheZlW66xfZy4hXryKXchAdr9hwvRP3XuEv5i2NV8wMbOTEunTdf
S9P80FXKQRknDW9d8fG2CTs8uAquxjc7SRAiKEob5zPHXFaIrugJPDddtqbMtV2AfeXihJIbGr++
Xcnsj2u2gpbOse4WZq9yQ//DTn+39GLoHObBE9O4W444uAiWzBPe6icwT8e83dPtSbGq6+DVno9B
joGJJBznV1PwzQAa19A1FfIbVAN81dXA0TcVzP/Md755ew2AKqR6qGY21F7KO4xvfF8Tf8xrbSg2
DRuhp687KX67J+lcWt7R0VWRpLWOeU+HDS8/9O38q4SUirMdOGE+3KAWU+FKMKrlpr/62jAAcuuM
wFSAh1gV7TrJOzYqo68yVUV2SGMO9ZxES1mVFhVQXu46u9uCvQtNzY5SwuoFIQ0mJQfexruKNbR7
OVbO5OfBfxe0sGs/ex/QY4mmLvvXdf90GRFxX0MQSeUnSjVHBvxgj07clnw+Le6Hc8WvRZorzOT1
cTr1/Zrdae5PRfR4VqWZ9aiCzfWdQlxHqhXXCsP55MxP953e+2Mbuz5/ov8xlclDCwrCE20dh7PW
91/1KaFtpLDUSN6GafYyONRB1mEH27Z05ky2Swb6YWG2wabE3AKFYeRfrkHlZJqeelCWk8LVvhSA
eMhF45nN7ql5vhQw6VXyr5vz5GMKKhSGC9fms3NDea4RlzWVZ4gQyEDAmYmqzPy0Xt5B5nfh/cXF
Kmq6BGpd4AyDb2mc3AJ5VeZ6h80/7/RVk2qdNna/D3Xg/V9+GxCG0qRB7A6zm1vEXZRLko7r8MdM
nvbtnnHEaxVGpGuy/OThGoXYPAgOWVKxL5KVPS7q3vBVzoSwfFulHvJcpm4VNc17mJr52vL8hEHR
SSwOTMEOJtuZ26mGDcJustxTDU0i9MlZm68x6/D2tNbnQE55rQM55yVLFz9RdhcR3NG/IQ9sKGSZ
BUoq6eeLh+9FteBYaf2kmJdCiWCCR3aMjZG8DLyUkNMXX/zlWj1nvanNzW7528Va9WQs5C4b04qn
uDKPvISU5xhhg61LIerwFqAJwT9eD/EHCCHHaFZKICjGpDkRL76f22/2JJh4HWiMCaIbjP3MQora
50rhuhzXGQDzDycXIvTHOkzJIRg9ub83rQK++sVfFto6JkAEWPl3OaFUkRvCVZl5HSGHhElT6ezR
Zbr9zBeA9mBrWOaB80aZGS3U+N3sdFLA29fMx1uD94kmxOyLUpdsvEpPurdN0VFeb1UYAItIl/a5
zsVuHtNBS97gyT5gTlMQ/5LauiIWFxtLoImVsmTtNLmTPVbWcGrRaIX1z7Na53mYiXNsWf2EeY2f
MN+TqZz2Om9PJdGJ5GD7qL6sYcGbueQbf3QENxyy06OVtGL4BXIGvAed4fm2IDuf2QQLM07dM8d8
4WKRiVhVtyj3xMuNQPvRj+nwT7N83JkSL2Y5GOxSCkGrnBaT71DkizCgA3kkxRa3hqw4dygd5ksx
Jh44NV+BgPIm4dOgEqDP+cKh557+bKoBWQDdbk5QmPRNGeN9a9zMWzYv8YUcfOylF3lZ1qG39e5u
nsjoT88waD/z2PUYkFB3Xdd02lr7QT6Bq+aj+f3WgikY82+zsCfu1+tMUtEfHKwVzL7MxBhHiAuj
Y4XwS+6Jbhp6jIBuInYo0g/Obj9rTLg5EGpzqLf5GhqnmMAbHLDygklMyaHaKR+JBhVm0dj+Zsgl
hMbbE4m41feNVzJiqXQV+AlNzAP70IcxE7JRJtEdAU0GAKlbNNnqzJ40XwoGwnMYvMQVDb5F9sJJ
sMiwcsch7kjDt8Cpw/4Mhrq4T8MxDXVyam505l/Er5Gh5zbEwTNtTZkxQ2MVA7ps1pfdotOckpsD
lRKQY9eDsNKYAT7GfdyvYKX9T7nRL2Mn+oaGVTTEsMtJQofJ9WzARVz1gUxM4NnZQGN9uZPC6bp7
ndAAJP+n+F54Fh3KdmGwVDb14fomw0rP597oqVG3pheN+MBmb3iDYg4233upUBE+Nwjhep1OmLue
IKSbNwh3FrbVcAxXMh5m6cZkiqGk4mR0MJ+VpZZANDNLOxD6R8Skcv8soo3JCxJT5yPi+yDW8BqU
p/Lp2bYXFM2MGdP/RLStfIT9HAyjq1lRnu/niCzZLmQaY1SujpJg8euM4ON846xyAI3U8oLtHxTF
dGRAzt4pcVwM+4nng46OhXwdAY78KjYDM7J+F77dxU6/5mYsQCs3P3OcTQyzHz6tVAgXd7X77JnK
uzYZ+jwZyWHg31NMB1WoInZEYwhz6BCvSOggQr8o133ATHwGpkI0OlPy7gXG6gYNXESAmZ2BwDlb
sgDRbJH0+kyTOhdQfzYWcKQxhsrzd4PVQBy7h2y7O6g57r5Vt9OEN2Ka9GpqPpmSepo5ICMMTFjH
vJbDduiqAO+gf9Gk7HIV+sJe83hPlo7EBePCZ1gn+TBNc2znvzE1cRXojurKXGM6cWGQ8PtR+1pq
fT37qITwvYZhWAyGBUOkig5d3VzSTs1ilCrO9KTCD7odxK6pLi/jSZUUBuoxwuyoW1PU1Vo8Akwz
dpxFbbPp2VoxkktmoqfkxFGsRJOGlh/nuljV8xoOPNEkyLj58eYYN4PIV066reQFe9qN+dH7Hz22
BTWb93HZVeNvs4iB74UJfXR+FG404AaecAa3E+llvIHxmy/wJd9M0gBdqKXiIl4D9LZaATWmQk2G
x/c/eO6iMdfQC3Ydb0PAMcY1yDgGXiIQ66VO5r9S6Uyd96fniEAEc48mytqi62WngIqOYKUqcPYK
isDYoM0PPSRRih45HeyfGYb3xZMV8O6/bOr4NLE/qydDy3oshIcpJoMfMRk05pJ47PlHu+sKRKZj
5DP6NixcpMktVDNnbwQgkTnWB4hE5+JKKNEpRP6b2qcvZehozl7C3/IzR2SThsjgA7z6Kzfcz56N
brxIBmNSYIr5x/04KXoUG9T7Z6DG/S3X3NG6L7d3ePsCjfe7waBi6/scC95J2+P1Odkb//LpS9SR
Qp+rvoKtA0V1GwIou/YDspwq1/8nXFMGDnldR7rofDXMvoPJAcNfQ441ITz6J6APlqNslVRbxTKk
T6SMTlRhFqT+49WTtFOqPqv6cAR9PDgedHgFyuJQtspJhKa/nk3l3ewSac741weg/eofqaSazSXC
AB5iVyRXAhy7qVUaS4qwKzd/XvJ0oMIMK7TlRC73bHykb4zADrby2fiiAn5vos5OVPksKk6iQuUH
+UKKM1wdum6HNmewyW3+0ZTDDjsyTo7Gv5sYyfEgjWT8Mb1CiwPM81mGVyIhlKxdT9kY/sp/2yce
hx3uTWq5OOmtyLuMdfH9U0FAG7fikLdOo6GRdDfaur9OTcE7jQ4GXMEygAYdXrnMXVmgBEgR6TFg
R7CQ4AztAPghAYre/Hx/GPimtsBwO6Tfeq2trDsZWNNiPB+7f0RyvScj82aowpq1GpXtUlkewi2b
y2Ax0w62C69Kj7epsbA2OPWMOSmr99JVenIUqQDVvecTjULPAy8SX0RpJG6n05xr5edCNs0ng5Z8
hjieAB7WopM6sTUNxbENGUB+4GmSWqT5lUyllimtmZhx1Iex33KJvJumHq30l5Znrmjl5f+g1uCO
2iuqyT8buRyWFvNP8+mmwddtSSiZRHYdI2lNFeCBY9X5ol+FkATVggS061T/InIz5fbnBS8NDJ/Z
CBqB/7ie8b6Vxth3XLTZOkK0UxCIE1rv0u8Qztpjjd/k7chh8HOI0U+l58DEcfgmxl/Q/1C/1C53
y+QsCSvUsIfZoA2pjPudY4wfaQcQuN7MaN15FZMqPbFq9nhzOTbSnlkZJfuMDjUeyD2rfjbeYmH8
Qdg7BK/eVLAT5KkIytJpB8M14RTKO68xMn466FPFqEFzNuTKJM4GbyWLNwUtogrPDlzihbtjj08a
i4cRSso7ejoUEULv5Ismq3eMn8BViRE29QsL0qb/zmvLiB5DRNW2lG5RUWOqjySGe0lGS2/cwOev
r4J53qOS9HmMQLsOE0CuZ8CQw5kNLObiGilEI9z8GibSwctB3WXfDmANKYYmJEzUStWXQ0z85Qmu
zZ9hOGFmPZt4i2AMlmF43Zqew+X71NnoENVbD/8+0b6RbR0iOqNKLsDc+7D+zX48f+7Hl0r8BQeM
maGz3rQYT7olbQC+LtenIv1NV1ayPeCYecyGqWzuETAvKmFAnaia9NR612gAnoQUB4tPO2NxfcRT
7KZWCHvdy38FKO6iDWNQXPdUmL3JLRYVDFQCKlV//FoLkCYtAxDyZKTiv7z356yEpS4wYEldofi8
ShfEA1vqAwfTY/oIekybC97YhHyZVAgAipSS3R+mU4AcyhFKWgJhUZTXXG2T8sjDY4KnB91VM7Bp
19Civr3Y1n2WThZyZTdmzm3Nkr4rillhEFBqDDQPk4GenfPU4Hs6EiaaGXYqhpZvZO8hk1z97NuN
qS1sHBkzch2e4BKVfwZ8uSb4AyXA3xVylzHfempl8tWr4dcisHfm1TfqltihHuO+y+2WVhFSbOSd
IznxYXU+oozyz7R+QuW7+5exI0NDCz8uHdTrk9kALsc5TK8r6sSXSlsMqvAlzplB64vAxSuMtFRr
nlW58/gS+DSEciMgGwtCaU6T74/Dl8I6ULDsnShmf4hD4T2otpKccH5CdjyicIVcLqqT/mzCjhZX
FibfifXiTYqm/byUdZFVCDtuJg1q4tLl1nBWY3osV6nTR/SaC8vTdcfMzuk/zrRFy2rGflWEx1tx
ViLd/nb1KdFKcUTjIjS34GDhcBRrXYznnmk6YBtkCkvC5j2djGTwUE5u9OVMjHcGgGUp6Nj0JvZ8
bUKs0bR02lbc5yfA+ao/OmIzh4LGRDdk7453+CnbD7ynPhua0fmvNBJUYWLHfQsGQjivm/C5J4KC
HYwezgnUSIIyLf1TLEt0Ex1E9jt9wS8nkQ8qa/slfd+g/ibK0fVdwIn09q2EJK2IhhzBXNM4ECyM
x4vXjKWfeuFukV3DdJA4Ppy/nSl0fYXX6PLyZaA31GnVcBILdLLPjzxVul7aB2WkRi6gKjnSKaEb
75BsUXc+UPPh/TsrV/D8T+ebS46vOZFrY5QFbyw7JSqx6Ag8qCAbLXiTcrHFN6U/i/pCwza0KPSe
xbtVbkCDzv1WIzHn5y/x5l8uMVyrBS+LpIwJI+sEX/UZJfECmnK50XmYOVF145aTrMb+T+x5dd9i
sXebcHfRoN1bIT8I4lBogZNzIWw73YpaFhDD8/WPCLQjiKponNbbiCXmr5jdZdzFutznUcvjawet
LVR1wuv90nfTs8XbqDPuy1K1huzJCApktIW6T4V+sknMrSlrVgSHXftB1nSNA6fyfAed9KrWI5xN
chM4VWvDh80iDfL1+G4QfzPBuibXoA3oFMyEN0HWoer6jTQHIFpjoJm9z1eCywuB8lAIavWrA9IP
DbqnPEcR+C+IY7J6We3Ro9iIlArgU9EKrRhwrtn1BPwyR841ZhkBXEFFCsJxMUemI7nWgm9sVA7Q
6YnfTTWUgbCEPtsXGNR1EToBcEPA8HwlNPWd+AffhCxuqiGa3NyBKUZF49gRVI1fNLeJX2Ev+9Md
IMWLf33fNoCSXye1b4Jwxshk4ViBvwa8KDmoIScLSUWHpjDtfWVN25fcMGSUL2tQWOBkbosNBfgO
uW0Cuf4YssDStfOJ3v76jz+65LJE6SACRh9BUzUrpl5EmRi581XnnEzP1G/gxXQcoFzcrm++H/b7
kHGua+PqU4nGcKvb+wrs1BRGLr+8F/VSWVhrieMrrQHSGnuBpyD98OJt7qZH1RX3xswahq8Q02sR
h81blL9VIeV4xuNOQdqB2KlQP943GDTDCHvcMwZRdI9rzhRqS29oVIdq0Xv5fOeYmarsR9Wnya9x
O6GWka7wFv1drM9wpSvF556ZrMDdHDtc7OBUzdxcfhumxrX4af1ml4K5UiVLhLHk4J//0LpNABK1
jQCcR51UXE6YKXomf9nLiRegBf47sT0Aloh3/UoyGLt7vp5C6O4sq3nVo1JkOCHJifxhQJDcWwKH
dzdJ4asSAEOEpXRaEgSPIS/oXqbSbi/68JhVxQsQ5c8c0LmOBm26kGLwC1OAeYoKIzs3vFggeuJV
0BBaB9dUVf2JqnGD+bwnv/JAxBX22gmOaTxC17qT1iAfsagauBjWuLr0F+xW35oVm6wJjh6SITnv
LgapHjbIxMjJ/mQ0NPZAqJwleOTlp8NAAatYcB/Ex2nv75ISR8s2MdQZ77NmJzVW6xdk0MBpvsSP
OyOWANr5zmSY/YCY4SW4xnRK3yOo8u+ooCHAftMOeOOX56RDrw61TedC+zd2GQgiRQN6lAFng32S
XECCE1EVmQ4NShB/1KlIdSP+psJGwsVJjaVWlW5DcVJoN04Z+1N2iVor7ioeshxYcrZWpF2YYLMC
5W6bu4TrD44j0WQvApLD2LTZuCTD5l3YxIumm/tGRt27UCUib+QZMKXfcbN3TT8qP8ZSGv+Azvbt
oqhhIApFMIqQU+PJ9MOkfL5zkr6W1b5CmXDI1UvBfx45hhOlQzMszhu7gOKrQEjMJpWdTkZDo5Fu
+mJkQGGja25LHTsgSbJFOQl/R38gVf2jxCQ5kfiQdXfPHu9Z3lVEgCVLlEloBRshoc41HMzdqxAo
XbjXZLnQDFDi9AwXesyrxZND4zIlFAn6VJLBEG9XTUoXBjF5r3kuLXzPoSUjz+hsr1BZq4rLMRHk
QLKQOxvcJf73snJ3IAATjNB67eJAZBFSNmZw3gSu99p87E2fAUvrQRzPfc+WHIGS+9O8GO+INlWx
J9cL24ho0/HpgIwiyhctVi18AC8ZsCL36gHORY2Jz+NGnC7gdEgEFnwJiX25mASzO3K9DZ6FQSrh
pW2q1gGcxMH9M1MERNTLjOFqQSCk9EWvmzvvDgpUJPaaM7E+duQDj+hBF+q3DC/nZfWd5ZSVJYoP
WOBtJs5ihV4NP0JGEEQT7+4/0WplCACKEzss8HMFE2227njwTgcdFlcOjUgGz/HxSy9Lyp7R3eg1
6iXA0cf+t4FcIlkC8qBS0c5ilatzyNMWe1vPmCpdVje4UZglPDBXXvd9YJwpjdGb9Xz2d7mp4lUh
sa42sj5IPAOfS+XLkdyTzdfmW+bjlUB9kHxMVReQFrbI2urOvUJsbCmT5JEAVlsh7ebx5ppuMeji
+5V0zw70OjSswwTY2GROMAkP5FcU5mrpFYr7M/tUVQ+Mv5m8SSvrSg2Nwc38PebwzerllpLbJgin
MY6paM//XqUG/tlNEjkia0BRg8e8b/eNxS3pNIQGZtT0OCakNRyAA0L6k8TCLKFPIhDKGyiSDD9+
W1M2BIy17htCOeaKRfw27u8SLwZZfQVWndx85M+0o7LMvSKGVmHOMmlTnsnINGLiI1t4u2MNgCPY
ITkLQ9TJYhtjqYdUpMiDscBl4xDGtQkN6Sg8KsRPY04PpIf49JA5I0vK4c9OsNqxnULMO2qr35+C
E+zTaiPdEgGQjzXawgLXI5+gikL2V9om6VPb3lY+PqPPNJIcr2spPbiG13WiiqEdcWqlMY6lJMOo
Ks+a5PCuPi1nPMPr3IYMceQPBH6G1HPcIPhAAtGzaMjjHghUi7PRrQe+dCpauFCIorWFwJovKnJI
NoJ+hpOgE7MySP0f5GemUi3olBb0uH+9epUze43oUan5y1QvOZXCwtPE34B/Wz4b+7znB3EclAD9
rsj/8VIsIMwNVei3tPI3u3Tc+R21MoMFhkOp7SRGCq94WS07FSgMos5mSTjiHXf0N2Axe+SIA7D7
jyWDpxNZpXhxyUiCXsrlfaE1Lv+gJ4XLsVGTmGr7KDp83YQZiTpXIJOAi2yjuXHrWpGLmGzrbbWy
SKwcb2hEGqn7YBsY7pDAYDAFOwWxTszYXLXgE1iMfmdyC1y7IH3UEII0Iab5G93kZrNWkI1qKe+/
V1cyKqBiYFEgd2/+9ax2RbxBWuoJdGTxnih9d8NzclbrpKm7BpHGntpjYc9cUq8M1j3AzSWoeP/Y
J8Cu6r4PKNLVRUArJ/KSz4EC/AQvXkr9fFOr/g9Q1QbIzIg6mv7Wa3rTDd5rd6AS0Jfg4rvNh3Cc
5Zdkvl5KTPWmtH0pk0WCU9yAIn/WEPN+hA2jVfa9RaD7iSD3Y8o8bLWZhYZIVKIqdcIfmpmhnkh5
Z3TNmQSU7swMYKXpPvSiHB1qClEE2qJly0UDIyP4ZABKz6C3q18kL7DXDvPdMpV0dvv6MegDTLnS
U/IlM3RSMeHAWjfo2Eapd+Duex8VMSLTmjvU0dGK7eRz+L62Jr75JG+RTZxWVb4yWl5Ki4HXcCKv
0HepMlB4T2FFHEJ6KUlN70vqeeIGkvLtjwMYvflCzTVrgaq2BuUWxqzzWEC8yalR+GXtVq1TXIDb
RZWSM3wtCtnW6jOUKL+uEvl7MGbsZrI0B8K6AkYzu3hcJOQ/P9GoeEeW+D3X7nQFShh5qA1pWpda
68KJmUBppwLNRSHKzCGo5UaVrAy6FrKENSL8NJ0rUxjImJwCDR+AsUDtgy4Iv1T3RVj30HrcJDGi
TdauE8qtELIeDz9m1WRqGCBcA+tEP2A/1vKcIJtTHP+xdrMHtDjtBXbuOkPuVmktMxo2gM5OGawy
x++UeoY3S9oa9A0Pu7S6m7DYL9HZ8jZH/D54LB/Dlk9KUDglKV1q7OC4Wd27cKC26jhfP9WmrElj
Ysq9r5QuReAgXMHBzk/VdVDkO6HoWySuBZXKzw2xHXdiNIJ3TqswkdSce2TCgie/9A5cOkLMWZAA
wOR1LmZ1haNLvUB48e32XSwY9WFglnOVKUahNnjGe0FSu/7VREYrvm+xjRcYKMZkdFGyN+Oxb/Eh
NAtGPtFLenBDoQ/UCWvQrx7B9SPqqASfoWMAp6iqPhyPfHCczzbWyowgzvhf3o38L3Y7oS7buf+a
5GnSAtAqJK/HtjmuQgWDVH24INFPTlNxjgO4BDOFsuUniEsRGnhMeQjGXKbiMwTX8CD4O6VOyL1/
ASfzI6z5CeHYOGixtW6Mlpz6hMWgwJHAdd/bLv/fYn5C4lHA7Zb3QHl4tXUG5lWZhbyAdtKea/LE
yFi7i4EJHzq57k/QpYI/7kUP6jyZ9zMM57mtProMPK316A+95vNKMVJ8VNDxJ+KJSHbAIMfrIgYw
UHTmyMCf9AGOR/WVh2xuD95vttxtZNJZv4ss4VcOKL+st63uRu6VKGC92atHvyuWzJ2LHb5W1upL
AgSU63eQTtqKx4orSNL8hptVGrfuTn+/xcUxtzIuaFxY2MOq6gBboSZcATPsDhtetycyP5yp8sVP
FdM6uG1SftCJJbyvJzOwVT1kjCvn8To/RfnjBAeqNuXO1G9Fyqg5rUlcDQD4NwHrr2puOzFiVLaU
Xk7oZCq8BCIGYhPHHMzHb0HcBxY7MvWlyupOYhH9hMPraDg8sTuxX1zvA0RJ1oXEHZU1fogZ2tim
RB58w7QYIpGAan4IqkTHCMIUIE0PPic9pQXkc5ZDK0H+D0ryHEql755lOjFOPg9rNqwZqN4ZDw9y
CQZIHlXGhrzteMYVsFZCrMxYpLB/1Eaz6XxktmAvnSt1bI+DvDrMtqWYwoXw1mr+y5efDGlnIXrJ
Z/8FhlW8FQ8qOTUnIlHaEySXrZyBS0E2aSDn1F9GPCbIsb3E06bNzk/HUgEctQcGTJJTrJsgE+p8
wtRhWMfh9JfcmQpb4Xlpl+7cZ+v866Ko3cs/7FbFMQSezIfHNyCKJLMQPZXKQJtwIPSNQmBCFe4K
tV0z/d0vi0wAzqvtfZkJ7H8lD6dcACgbXXpvnjDzJ2Sj4sXkKbZYcp4xo234sy1p5WiqPExZ3nQ9
L/6N8rONhDccn+mniKLFGT6Ucz1RC7GJLfw+2xzpIGKjtuFPRswqUUSB1qK+1g9MIAjGHmHrpZ1P
2ZvQ6p8W8usLhQF2qSY7qul4H0sM+BODuyt9g5gTR+u1o5k/BbkM5ExV0O/cnBt6sbDOtMcUStcf
Btt5Fr7fuux56R/ahv95Anz9nN1fTLArueYWyXPzOK/1DbwUcKbY43wZM5cNigFnt2XUh2wFzwaT
7/sh8yXp8Hjkov3Q4vjeDxEI8Vcrl3h8JaF2tWpxYi/7U6dFXrovdXWaKHUZlgCPIxbBfIc6z/N/
etl9LbX+Mee31Vuwpy5e5MuT8zXbMZfTR3nYB0nsQmisXH4RHinDXxhx9Z42rLCatUuaWHzwixGQ
+om0VGWCIrn5iKT42c0vhKfft9TsXZAXKSbepbK2pAGkxxlHz+q6q79846YXfiOCqQapswLlN39C
QN4PJmMlN/1PBpPo6rc2r2HB8Bp0ikYweWhF4s73Mm8b6cPCAGDKI1vc4yUMe6fQCI7Q1NDdfGcp
iejj4Ia6KEllyFQMOvE9x7096PgSe2KNKNwBAiQTmq3ttvElcwZ6/UwUiOexsOPVc2RM5b7aq6No
ijbzXZkgYsNHjZmsl0snbNjMDQZGnoEBA1PgcDF5pqbllZ+PBZaaGsumXcs1iRrqo79tZ363A2Z8
dxps9V7ABLbHIjIUnb2ejCKIaHL7R2SIRU6tiiTy3/60EjoIasm9cTmoB3rv6lKkPPZ+VLZXrEeb
6Gh6NEhZDb6h0pWFFprepda1+/j8uXb/OSaAmVgCEq1nz4KYmyHCb8tZtSTzb5uqH6q67dJc1GO9
Z6k/fe7Ht2P2fzD/J2lT/W+ponO43QsIZUd9Mh7GGt2QOAfCZuR2SDezrXPU4oUFjDDJAr/VBMVk
EwF7l/rdhoAqVqKSTrm78iHrlaQ6lnhQxfBp1yrxulYCZtrE3AraPRN0ZcprQ30tgaZ3mGR4Vrcn
XUHygc4q4QoN8Sun8LFEDySWTHj2XeGAIh3B3SyCFlHwr5QIqU0uNcb/d4/2kpqInhC2qkvclR97
ajmD7qoW4WUsYG0z+8ThG/YtAJaef+9UEpM9xGSHu762quMFoDkd2+05R0XF3tKwx7eoWJeWTi7G
vAA2NvnKpqopIH1SNuN/3jft2J9GSyo2+oO34MTnjf/RsG/fMngyXAmNmoFJA6PTzrYP/XP2LQsp
RLeulTMktbGy8GJh/dA/cs1xL0+i58XVB1JJpwSUxrUIUeyqCemgTQSOKkqMI19lGlJ3pYDpSwcO
3wfGDdaa1NT0JOtk87vLK74GnSys2TUIcHmCm3z2as21we/PyxyIW7IZ/LU/keI6vT+BqwDsdWf9
AwmwEM1zmK6BvmDPaG7PhZLNkHjI1Spn1UcwzMgf2fEm5tzZrVtvEAzMVkmOnME21Ex9ENN+OX6u
wqjmr4UDI/Y2vMsTWx+EWXIkM0usPqgf4G+Ii5tQAkQBkYn6ifSO0Ci4APT3vt5qR8tnaO1K7OPs
2EPw0ZKhXsZ/RrZvgmOopB7zZCwl2alHuQz+owx5evhvgC4m/kdXugR2uvN6Z2gXVTwjbKj+/Wn5
F4NBPckNHWd+3ql/qS52WiycG3HDgfvhMsaAXN1tbc1ZcYk0YSue54cNm8LU5YVPKGjNmNzDWvsL
yYv9csKgI59OIvmIlQzIP3ExfcTejXwiOVcg47WeZBaI2vrgeBCyURs3psyXsBkwdIBN5P4na3ly
V4ZTk5BxN9MMNEJ3yi1WNUeCR5hv0x69mto04Bg4T2qoo/MjzK0ye4ovvdIlkzklDuKwsHtXlX/Q
ae9lVWISLR0OrCpREdw9EPJWy2LO3bfHtsEXUgWrG33H3ahp0ljNv/k8Dj5IUDauzgVM9VLx0T7X
9Ft6Zdq2D+ePxJOQ5j7LF1O8C4hArvsWBa2YV5todK6d3gTFrudnQOQJNdhWFY2zsamioweM+x1Y
+qFBgR24iEeJgUv2FUorZCgr6bZxS55J6GEMJtiNZmR78L9KcAdNryMjSJVINwvda8jA/rSxtlcr
7NKp6HaISjkcomYej73lp4AuQB/gLfIE3vF0SBGXALDjjNj/EH3E42QowHotvLGTEd8v3YBs2hl1
dDy4jgH8wf2BPuF2tiNangpVZzf2L4sfIn8GGnBqIVWZ2Dk7xAbQSibKmtqI5LHnVXmeecoryoAF
XlmL5egKy75axcgqkMiNXv0vco/axAF/w1TQS8Zelne/A6XpFtDAzQwgx9W8bOYgcdvCjra0Tijd
NTiocstcZSUXVPEQqzRPBkCz1GcuZFjYFVy/JF4fCQYQ4sXZ1m42dRa+Y506ggZrd503oQwzE+jk
bKzzwre+oG0Bxgn42h39LZoSfz4vClzVA5YKwTv92txf1IuyqVwMF4RS5tWUZkeaKopareF3yBGt
FxaDWbp1i56mUj6nmgivwrWrgUDDolsP/HlvYHEV+xrglaagLknxJFWMblMPxGejkzJ5IT8JJWTa
ajPKqxnLekyFAwx59ivv80Rl/wfVhaapHcomWTWuuHvb5C2M7SkdkIuV3fSsf6anv8WkP4zNwtD4
JMuyUYv2KZ9q46NBFY7S8PePdj3+dhyg2enJkgBrMZOpX0ed738cCXsbjkxdrvFaMpsLN+CoqukU
vqKmJcD3Oq+Z6B5IezPOCZ/Cvrp+CZyWu+mdGPn8Gti4iX+Ox/fSRXln1ZgUPSmFCwAGjAtxl1BD
tL9wIYdF7cTkLHCIQyWmURUD4E204IIyg3IpGJhiFqguOb/VG0vPl0oVb0Kjk0ufp95Iotv+ilAq
B4PC9QREb2jNiJblR3irqGdiqX+HCky9OVNMp4CuVVUw8+CRtjIXQhXYaXO+/GKvLCiO1liQARoF
rDvP1vF53+7uoFGbAh9d0yXR1nAfEALB2CQqenwdwIFc8AuYG1cWxhEo7yNDIN0ZXtfvIFNnqyHo
MOfNTAySP3UilsJmlR1ky70z0gOhe7opSj8pqHqL0p8k+i9WhX+u60zSTEGoJgM0b7AldHN4uRZh
aamGZXHCgA36O5kudlk6uzVeT9xHlqw3+6VINEjDLhxrsIRyVHccOm3gXysp1zHelMtG8Wvd7R/J
iKZEyVF+dd1oHAW/avoP6vU0ooTv9eX2eANuvJPVqNbbfS9M1dH/BJfGmLrsOc7V8XFGXdOzXLT1
MAJNqdzjWDB0xfNjlp53v1kQiL7Ij0mPzYHLGi8G1IEOhGIxtlbZKS9RQW6Zx3iC5BmjqQemXdR4
UQf5JRO0bUIKQdnA89vZni2wE+jH+LN4B0JmspxL+/hqoyRY0UKrUHQvg4nYEE5FmITiOrCRF86A
GOLN75New9BILnLLuTFVc35WjRw4ul1yoDV25UCfzv8kvS2OwoIQ1CCRj3yI3PMCtubSljtGk4y8
I9HZHMxRf8wLvGeKz2kSi3VqCZrAtu+7I5gYykDxxUMnWWSW+gI3Ve9k0HCjcOrMPdxFaEFs5ZpY
x0IoTfX8tgDmDHZW4VqBJjKed2aXjo4GKL3bMuqgU8IX8MVFr44MNa1SDJiqBJBD2bAjkzRxERgi
i/+2aNsiI6wy/TYzdwbamQnmN9mTizYE7UUtUmeRWSHP6wmETYCScfUgSaZOKPoqHTvkTQ6cxfQw
xnYpRFgYiIHLcqI7tQmdUOk9iF8yTZltXiwvRqy0u1PvsskzKZay4u4PotdHc+2s5wB+/mp8WdvH
yK0DyoVpHS8LPSmzrJMjhPZU3hLe8/JPwV9uKFlydOhqV99gTxb71wU4ppqn+5/gjRhvEpqez6L7
PeObQhUaaQE2qeK7Id7lHZQnqaKsDoOpccg3wo7bIa0iV6xPD/UE67bNtPNZOAtOZSYHuY+7r8hf
cpzGsEZpGjpWQ0T1BaanBTaVSqECMuDvB63X+a2qM6miFalzAW/v5W6Lh0OTg1MsXKrPtPKRfApa
yIb3SCXW2rqbi2CnSey/wUZhEMPBqJFK+tyBxzrrl026Vk0LG++MlZTZHbiSS9sYxCJN3SkfCEW/
vE2hcHy/m80ZHIgjk+cf9kGo67UA2MVSOlDl1KpnpbE2K4AAlambQK695xsLFejPjRvQnPueVzmr
MZk6NvrbjEsjN5uhfFg9/FlVwYndOh8HtMQltwBEcNnl/p4VOoZnFcSaeDPQRniK9lT/pzf9NGHN
l7NlzJJ3PYbhR4cm5UjBiqahee4gbsuzI+vlXobrniXIEQGQNKObXXBt8Hd1QkzFjOqp8MLS+Bgc
v3tNfNhHz9bdPTpTw8COyHrcU6gGiXc8VYlg5joc/W/IHy51Ctk4OkXHQebFbsoABSTscSZnBEFp
xZvMM5L/scciD46xCF8ex8N09XkAQD/2ldUrhCxzX2/qa7W4b7vS9met/H9hqbwRQ6Cn/ln7qBJn
vLyXFRIpdgRl24rLEYZD65epBUrTY4fw2SXb7Il3HLJE3duF20YrjZCA8k2qTwtmqgWATXllYjCy
mvJXnvvJKZefvtC7aYP7znby1pCn/skd1xoZZeRszI1vjfIk6q9EUF9NWd7wojN0SFnpy+R+WPfn
MiN+SE6bc+keR3sMJTz+yFqYY9ahvycG3WW7WMXWBc2EBbkclLEbI0tWjDPekvA/fAsRhYT44eOa
NxHJCxfLazel3LHLjmZ/cgg4o8waSbTbh85I/5rrnXplspts2zEipTM1ViI7gRWg9RQVCPubI0bv
ku3Wr7FDETwQHVxRsOmJfAwQAoODqensAppC4GvRwdgVr+5zQg+QVlHsY7yc2hFYxCGbsWrmb2kZ
Wa6edIlSnXz7hhgnn/XTI7k5sBeLVQK1ujpCCj15C0raZgju0mmy2p7pxfTjC7uL7ceNXLLVrhYf
GUnYNKXaGoZ9OcmzZRv1wQKYXezKrdsGUsp4HeFvNGiw6aC9cM1YPNVxft0Dud0KmIgEGivvJKF0
4n06OmMDHg1tR32r0mRzqfcQs9MX8JwQbqnw0eu5nJRHfiZmzv2297x/jAlQScMxy1Irgwxnxl4V
aT6jnjfgm/smwH5BRkI1J0APiU8WLu+wSOU9PyQeEhFi/jSRCL6w0CKb0zYFp6J9TfTI+QestwAL
XC89YfrSErdCtdDBD8zFkYrMOpMSdRNNkT1HTy8+6eNHrPA8C891kNECNyRD/cjIIWDa1XsPYHPu
5yPM/uSRfO8EtFUtmqsFA/SEcdA03Nc5ueuqEIQ8me2l3KHC419AflAQZbQSESsLwhr8nvnGfYLK
gC/XC/KY69Br2LtAmNv+6AeN7sWIPuqISmV2BhPay0uW130bkRDlyrBYBDGoX8634JwGOZlZ0hJb
+fsUhJmtW3D/7osQKLTa7jm5fRO3jw8bn9WeadfmMytR4IHI5HPePVLUZ31AFGUSCXDY0l2uWyo+
dmMVWLs8TpRX2vmF11XBEV/MPuViO+Vq7FdbVLHmVapX/00KTETHqfDjiAypSfEWb7XluYqwgz6S
rzFfPmKPyf3e+/SW54c/d20TTbrf6S1sYfrr7waqXu41Vo7QVWg8JJH7NuftNfD1cjxuk1g7OFqM
/XZmCO3QoFQonL9cwLf1LmhUtoRYPRm5fpeJ+fklGRdN2vtlK6qh7lpk0mv/nn8SI94HD7PQNofD
1/Nc+BjYN4DiaCDjMd7DiYO6nHkwbx3j40Dk5E06cFt2V4A/VZYWk2U6h5D4LjEpRUM5tivRteUD
j+bRrh+DBRzB01kAv5gNuwUjCiJibshSsm6UorV9KDHmrFHdg19hrN7hrzBxTy7s3bEXy0vz6JMR
hUb+6yKf8nuVujqyiCVCpto1TldszOp9wfN68fu0zbOVNk0ipqzoN9kR05enMZoE0xRb465MaftN
vay56h5f6bmzGJq1roPIJYF8Ai3HE4lNWx3mtM/xibnAyl12kHPk54AI5eSUA1SwVfrxQIT3NAUH
qjRBGee42fPxbdxU2K5SbVrL3FXLUgHeWayhr97mhFPu6Vjaukt2xHHqCT1ya1Q18JKbJFAQ/dZ/
VEThfqme8cy7hcIZigIwm9mZckC1XfseJ80RCGpfOhkbnc9rJLLeWpngFsEy8Eo1RHZjVsbVCW2N
3yiwZgdb24zf31N4rbIUy0gC1s4fJG2VWpNPtsE9Ya3/CToEqwyomhOY+4558xPXhX8fKlTh/ZMp
eFqzoLjj7jkW/2vMhg3IzEYkr3uOpLMAW1URl28wTNvLEjyuOg5h16DtHk1Fqru9jV+O5W4z3hCC
Bift2TUWMFiF1jrhqtAz0VKn5m1VqGvjYAEj7NB0BEOO5vNsxMkGcOhVLhm5mvdwxXyri4qdr/XF
v1TerFGsDEy8jfTg1ebjAsbEO3GZ5dpW9VyhX3/L525s+ksWSgLDD29yP+EB2OFi+5pJM3nhPi9o
tBqHYogxS/4zCIFKJGuH60bJUx1T2X+nAQpJxpmxDMKbjrbu2RatAn49kaTN656mUaYQtEqT3fai
fpRmhVz4I1/fn4MNMk7ZSYHR2UCJWxSISx6TOmKRv/2qFdCFVwgvlpuutzyGrilsjVsW5SxbmMaV
+ErIlQBdLw94xdtgj0wEY3hUSo8qQ3mYP/4YorBPjCxspc+Wj9GNNRHjqw/2bx/1Qr4bS53Y+BmA
jO36wA4wP1Viker/wUp1Z9TKDqKqsMRrDfVT8rfc27LrNg7ydmnU5TTPCKp6G+GFvvXxb31H67LD
RNoJHdR9Z5/wEa4+kNi8hVKIyWA2lVb6m55MOaeauRJl11Pa58fui6s8s+N3vlZopDHbe2CZDKau
zH3F6s9xwfH1R/KZ/SvCUd049na9KjbuJnEohOx1HPgTHRHTtjqarlOeEXleB9jWk3Z1LVXyNuKC
R79/H+u1+f0VXZc8GcERSg/Wt7j3fOoA77HsveOfLEPrDyGl9b8WNGwY46xY8Pp/ePy4HarBwyCU
0NToTtjBvA/fndmtfSR5SeCHnvAlPbiSXD2T/GXucPoeXSpH5hpXXOizuwEPgEgio/qkT0nAyJA0
pzB9WnF4F1uYp9oGSPHosaIP9MHRrB0dRURiZ9Z1DCn5XCcPQNgX9CFhf0gdx13UmZfM8JvEXzT9
vmVqc3lDzzZI2AMJJlK4lIQKEg6n6AuN+nYkNj2UvXy66nQIukJHQtI5bilDlxocraCkwRCud6vP
uR4hVsPXljqHxRAJD/S0E8yA8SkGQvE24G8g3KCCOarvYwJU7baQCruPPJqDqhADERX3/QIFPRp9
Cph22ce38H0XdG7WyqL8npAbGCoQQvEArnpXflmBPdMHqhSeipZYHQnXESf6cui9ogc3q52omqPq
9LatosVAiZ+TDj+zQBNouy8Awpiw4j1DaMrmOVMhITgP/ZFpKYkiZik5jC8io4uPcdOmu/BTQYpY
ImpIy4cxJldfF0EYOS2gsgr/ovKL1EbXSxi1zL6X1gMPeFWfezkBb6zlZfmAyb4pkmzNzYM6mnBG
4GGnoB6i+ZjezcJqmfU6GOmuve306msbvm4zUXwsCjRnwR8DH7H/GZKylkKulCjbAMclOVws4qoS
5KzgKLDHTeVHrjWdBNLrczdlZUXacBzDEfTupoOkvn0xf6ABC0ir3EMx/VJ0J3SuhD5ZEzQabTKa
udywLUEhrLpqEqLOBiiWVMS7JvX3oY5jYc8I1xSfD1UcoYfrmA1etBYzwFqgTnOhbAfmfRJ+7abL
L0J3RXoT3Q+cJynnLbbhA4tWnfzYM0WOOIA8tKyhWzrmEv0o080XbkcNjkS+NtAeyvYFBE1k25pC
yGWDGVatos/l8QCcGWg+GkmRWAw9/Nmg4Ol9pWM2Dnp3a3gpVxMCveuHPY49FJD6P4Gq4ZwgSnwd
QBWYg3sJofvdDoKRyhfFzJCcTH2aGVOHqVH3iQ/tZAQE0gl3TVCDDHZIqtMZNSiJA/F0fGFTttfH
gWIG9uYiFAQcadovp4xNrdXlAjfU0AB1hBeSYlIF9OwHUWdq5PYlcdC3eNTOzlVeGSTRe+a7TCdL
SQe4AOLRO609xUh/aAtHG2LXJVH4eZQ63hprenEsoqR1KI/CQBC+rKYPU7a85KIBi/ITHbsIH8ak
x4mVD5aQ9FEMrqHcdVKOOlr7VJYXQElVwklIwlSI41t5+UJWIYKztyVAcmPT/zabDftad1ceIrfs
ZSyEryt+xFTus+TzikoDLk3CjiH8m2JOfTiMpfgTYo+VRKldMjFpMCZUA08Jh2N2n2CXryv4QBal
o7EiDR/0iTgGzbZjwdz+mQF6VOYo1zddYVM5lBwGIsaE9q+aX49oJU9WRdKTTZFqYVSz+aUdpVsh
C/DHrJrP+BhvM0Uhj45zPzZToOI6FiEtL5kxtITShW3gWSChoZtSslWZ0L0wQ7GTn3fhEdhStPgz
yeeFLjRwDdd9+Q4I7WC4PiRtqpF8UOJbZX6lHI19LnW2B29mFZg0SGrANFg9UC0O4dDmpsBRZqZi
9IjHI5lkhCfgq+UZpU4QCNsXgUb+iktKPO0/BHphSwqWq0fyn30JNNVsd2dgSXEgFd0ncBDff+ZT
W69IdHURb4op0wYKmVozyPo4JuuLOcR30j/biZl51ttoldVNVVjmEJhw2DRxl4NjwkxxfIoDLcYz
GsoQWrZwrtq6nojomCneGvWzcOClWhDiDMBWPVL3Mvaoc6RfKjBLwZ1bUaUNoBd+YI9JKwnB1BQS
oU50KmZCc+HtXs1vIcKjfhyIFRIyfDZqZkWt5vyHpAhn6IDtfXCFqynds14h3s3Tv+6NwEOQ1MTn
ei3sTfJJKMOYBdq/mQAyjQOdkPG7KrNPmAwfsPYwwRiQdzg/VxYldPbRvrGbavExDs79nhsWOOsf
utAEu12wNhX4AzVAmSiuDSx22g5vjzj2KGyuMyfXww2fDajfEYf/7C6NJmlWdrmVqxIe5+FtUcpg
cx//aNGjfzSl4WN/KHGO61VNG5t1LFRYIgpi5ygnMTqA0UoSjE5SmNAtjnBSEOAtnTX1SFyMQa8B
3C5QWF/fBLIrY8sbuzAduVOWQQBT2OoG/rKW/qIhX6KiAzw3KRlJvjYjzgga321ud501dNIJwRAm
HjSEZTlv6tcup1MTszwRKI7Rdh0LCdhP7cB2DcVF0+0KLXrr5XGcTvxXk9PqL+Grm+7/tyeC1AQz
6zygpuejkIZK1nZAwVDLHHioZUwTSraZPyTZQhtJLdc7S74K+ow0M6jVTcBbRQ/u+aDQ4Y+a1JCn
P32oy1cO73vpboTh0CBaWKnzWWwXxfC4+vPbAFGzA9QnG/IEfB+Itv2WqtIKsGf+AwiH7xws31MR
D52zqzwdjIufYsElmYXHx9r4b7yNBGU06ML8qqvQ/VQqrnktRNT27fGgKw0ZAOE25T6M75JQimBh
7iutd4olzrpu8CQ6RuzpBqPlryYFfk4ObW+pbkbYvV2nI2InhjKb51/2mTq+4Fj2Oa8xXUhpBvtH
6152AgkmJpNKEqAuae9HSznAcI4EOL23zcjCXUrApE3634aKtyR8/oA6zcAlswGVOAzmn4M6PeXs
FeL5b59UaGB6LWt85YyaXbRr1YDZbPqV7zsKsIg36ngRC9Hdn6vB5Dsi1rKMPYKzwqjru1zvbfxj
NzcH+sGJ6swQjLUxWfdJ34OrurAObxLxm6JqFTb8dN0zMAq3D1jlbKrCGRsFfagM5/gwOx8nHlA2
CT/sYg3B/SuvMGSouQCE2U5mexDHirxWuVhJMS5y8kzXd4sBB+yXKG72vzolafsd8pH4aKPEQxT4
ZsQTbdIG8IjwXXw1+7jusTsifPE2nGuwvb8tV9BL+Yh2Vsm+BkSLkMUMuYvhGMX8LdvJS9OsGzrR
ot/2gTlFutWwAqthYuzeLsone3+OMumVyu3gveeXIt7v59apExyqLA7qeXqugpDZTG60NttwpyuQ
AGcsDHYYnYe7apyLmD+oA7LYLgUqvt90jMpwfp6O/LnOnvuEiGYxQ/qseQBHUHTfqP6n62G/vsja
ZV1FtQlL11y6aronZifY+djnf8i/SexGxvrlB/RfxA+Mdvds9lLyyRcH72b/b7PceLNg1MTo5mVq
xJyad0RvBgyH4x1uyR7PFQSSo4+nLVnzpB0zZmLY8WUpyBqTumSvQxacRBYBiTD4LTfF2vpB5U4n
YQ4VlXkEVJAF3pyqk+JHHlMmIPynH99Ujmu0C+ZH0vuFoDZ2g5/7FYeAPd+CwCIdeXS30iwgtp5U
yGZ7KwSj0cjy0PMcZyf8n+sysvZZ9GLS2QmeT/JsovhSjKb+64bcr6GgSYdnLia7IAOUuYIEcvPS
cEVJiziaYr75zTzs/T16XE7Zo9Kq9PrDQITbObhi6o8daZHUQi877htF9zMo3+yMj9v/YTldHCRF
r1tErhMRMRK7pfDPRyMukoB3otMHAmJS9OsaNYwF4M2VqdEUmHhe7Sk/MHX/Zk06IJY9MkyrrF1Q
s3yWKJZDMU4sCvILMjoimK5Ue8K840WliO+OVZXm+HdsqTJUt9EDKcqFNTGvRMnpmIDBPhdnVilK
qw06qtnM0N1299WE/X/RQzoM/oacslYpW3qEXhRiDez79P7nOOjpVOwfYS48RDOJxnDc0+kDpkPb
iadLf3Gg4lLTKcJpSdKLJ50vaPiVbH61fn8tD5C/S64YAt6lHsSplXKgIizV2f59J9oAiwE1eL6w
9OzBZrL1JE2s7fnzK0XlPXM0iyR606WALuD7zRhu+3ceQfcJuSzibrTNLkpwh6lTKBvSZP2uxLXo
QXHsATHGeyemwpf90222MZHVoZ6D9bGh33PjrfLUHILbQPTLlOYNNQY8R+W0LnX9Ahc63EApkzAF
6pETxa0KdiCf9f+KA1j+p9jml6dhJnC9M0njGlBWb/NPl0aTz9E9wBfN5+byQbmjOtiKgIpXMNGg
dvMUFVdCMdDO1vkZG4dc/5W4h/Ch3UvSBaWEcvEoXvoXMmEaNEZrP30kIY3eYxaCF5XLKgUL1kYY
9xySyWkUbNH5etRUHruMCBRIJEsQ0ncvhBH8uNM5ysUApgLNfobQl/e5pbMOWnwXtdFti2hFU1/o
d7W6L+BtH2hMlVidocq6YXc7odwHbys/OUcpcURvPOYKxIknAisNkKugXZZTDXOLv1g45XxaBs0Z
sM9xryvbPY88ECWz9o3LFjdY2EvP04i5YNNmfLNRcchj4d7WJH38cQ0xIwQX3naxX4jfxaDpji/i
GHJ4gfTWlEMpxF6aW0+3zwtV7FaD2bhY5keNeCw+LRTMveRwtkyZkHa2nkKvgw2Pp7ditu46xMfU
+IYP7EUEC+fapQnkfwoh4G3uvs5JF26PESPWCVBqosNtbJ6Q/Ug4Do7b/WYn2wa1egt7BLfcSBKe
TEc5mh73MbXh4VRcPG1U2lh9hTV+F+K7OL+NG+OrZoetdpFXL6P33Q/HvZ7Sm7LP8QvQJtUMulH4
2b4nb3rb1d8QDi3ozS2QS/CQnciwvP2/wL5RTGvY3OvVb3Q8Hoa4vksM5ElQbYFK8Y+1KHCh01pM
I7j3iCpyfHZjAvNkQpnVOoTb4rEq4d04YQakiD5aw8JyukBnKDodqio5Lt6uHRPU5GEpQHvJwD3Q
HewSiExRQNXTzmHsxgrsgHlcbT+cRRe45knMANMW3pTteEOdJ0HNz/zcHEK7fYEbAGdrVWviX11t
hEO/VrmgIB686VelQ3Yys9Am3WHkvKnWnKc4VoUGLxwz8tonpHcguK64QqOvYpTk0vMoOJ8jtRd6
hvZj0p2ZKF2HyYR9s11pYZJDY6e7lZKbG6YdsEWVA+Zi5ZUuNQCs/6aOnOLzzc683wMjYX5wo2fQ
G4rYx7FvwXieElwaKhWgMj8zWMuUgzhmcgd3p9gK6L+sJJUuBnICT1EZ/PlBSmA0skXqL/AVp9PP
uf7+PI522KUDfCuUPMQ5Su4OWSiVzJEAbYRF8yqT8l6n6/QSQT9WBQ04j7IzwcrQw6MW+A0YcXY+
PEEaFroR3auG3PCl8sSIVyZ6yIztkC3YydBindhpgcr0WQpzkE1Zx2vdQEpZTYWpucw4A5MruHv6
HZ2L4Hi7XhBbCWuv0DNlqj4JI20QI07gel/UZ5eTeVzptD7sL4KnwxbX/fkCRGWQKjmv466Bk9Rz
yvnLhSvJSuj3Lg5XUOEsa6Z4kot+J8fO6Rr73XE9siHQyVGLqxtN8Ah+D5HlQIYcJMXe0cfGd+Yj
ELN1aYFgvWsYdhmXCj50I8FILlWgxefYrZRmlZs+MvaGLSjDaOgO4vakShXA/sCULmdJsNhLaj9y
hSvENbbsfBJ3KJZCvcIHTmdrEWJ1qw7msm1RwqYdxzyeeFhVpTnURcp6fAktxNAqFNWBbd/yqTQT
J7d67xuatabJDtssY4Ns3nFoElSGObddYDeLLP8pA+0gPnN+yfaeELAKHa0S+Dwv2oKkVX4dPAoE
aTI03kXYZQX87egkcFHgTpQweGwbK/LFGa3TPKAtoaZ0kB98Y6X7q0D2QwD2NaOXa0iPlXLGwcZB
q0cEVBpuYDTe3AUHigKkOvtCl7O/rPuwLDOWRng0P2ksAC0jCEFtW6JTTElXdPHDMgOKD/QGqK/i
904gHSoKjSNzGA38N/mWoQIp/RaFgWJm4WLxfIiqJVEzBbiAyLsiggSwGEvlKFfcrh2siyVeNSKX
9zmzZZLVuRxNY/QkMwCsYXGkWcZWjRouPxs5WHxB7Y+VAT/efkE6j9Astd0yRhP4IUoDV70FXGop
RUACnA6Ffi8e4azDkAuxTsYK8Nl/6crE62eNnp9N8OHDMFUXxYVj64/ryEZxgtfJrbZlBXLngGMk
xU1KPVIbqNJ+v6q/jAC8hZzY8qLGAi47aTDo73QSPZ6xdyHpkoitiD9ad2LOH32q/SpJKbLOsEBL
iwTHw2X+dNdIxcIHa65fOWiSU4H4pGfVkBxO5IWIu3/SFVLgM/HgdXCWMazwf2GkP26WVQSyXUCP
rnHtLV5bXQW9CpFeeOyvt+UtS3jxYbO+b1hQMhp7X+V8DNXxG7K2YNd4PdyfZ0YcknL02p6mUz58
amePBeG7PDQMzmGqQxXCEoTFN8bbC4Is0yMesdOA3TaM67OXI7RkEH5t8jxMRmsf17emvDtK7gDt
cFB+u1eVg1gMy21yXYQ7Go/4+ed4jxLpK8ELwov3CcHoHJgliM7BP3NzN2EbDmJsAC/FSqug9fuN
BkLeikGqszuRrgmsTvKKFbVL/8729UbhRlZ7s+zaKYLVO03T6k2XuXErKW3jH3Z0Qe38zwPv/Bux
8bQGoxAPMG6ksgBQQ7N4Cg3bro2VvY/9hEfF6fKNNNefBKgWN4ow5DaGM7mDx1UGGlA6dI6+X2St
9RJGwBx5zjgBnNvvvvCs1vfRPjhIWKILFbGIrwHJ3suUIfR06TxP6fNBxe6YFCve7tHApX/41x6m
irXADp5i70haniK1v2aGRQrVSilyFJGUmlNzDSogSgh7uEUbqlK7alMBP1u/qR1wMeZ+DUi1cSkf
Jysa6nXq/qFzYrHUbVMsziPdXIKSRUZB3k/XCIz2ipThBLLgzfU0jp9Tlu0zdHzC5jmpHifVZL6d
qoU8FtX3JFET8JG/a/xK1SNCgAFp3waarycf1ja6WrqOXn7saG5vWUMaPL+SP3lq3b3WixUXtmQz
tnXpIygy1O6jyEvV2k5+of4sUDX8Tz5ZRGabTXWDbE3Lk5tlQBslVM5Z4VRwwkasHhRy8RQTTWAj
wGmLDRt8Eorc3O7DfYh0PIVX/IrYoxUmI0aKkrPXM8OZRqGVBbTrWy1uZy48EPyx1f4+hzlNPxHa
rEfvKfiULPtiR2FxY4TlQj/KUDdWVJFssiAdKwijObadFVGm8IUqpUSz3S+2ckmUjMDub2pVhPLH
v1OY618GMtWWAGN83iPnXE6RnS9Z4IyZJ+XH5oTcwsod2A32Y9ITwBkohCbmb+YDrXwqrMQeEcz8
GJqWB8SuNqW4qmLAJTv7hlrX5D2d055iSaQg9Yi+bPBwPoi5LZmpZDCXjp3tJ4NGBlQ+HbSBeSDJ
asDJ/RXP9Qzay3Ebc/TDmsA+VlsXFmiKuZoHNmn2IjIXc142ykWvvWUtxpvjpHjS65gMDC++kaKe
uT586c+2jelkB8txyPp15XP6A00ErQwnIhfHHo0SoSuxaeQW7pXTc8paV1JHwGMWp7m+FQSj4c8e
3+vkhEvjBz5DhurFjAdwfaDLYAkufLX99Yupcn+qhUVbwW5XrwpLcdKporTVUhGnT7K7NN5gH89f
WTkuBt7to4n4y0PST4MXd0Pj+slAMFs3eEStHtSR/Jjs7XmOo5hlJ4fLKIa/wLvC2DkjqyZcgYXH
I8+IMgkmhPsDVv1EOR11WQaJypcu7yOf4SdJ3iusftA5Dy/aFom3wK5AMugWBk7bqv/TRsDNIPZj
Yk5paUUVur6qNRSbe279AF79qJzzdF6XOknt6yZ735OPW8Uw++50XY7gfJkO1D+OOKlIywRwFhZq
7gzliHjMk43BnC3RnYJw1aEEtf2sEgFTIX/aFVRW+O8sDOTmzy9GxJP6UmF1bcX7a7LB7ytxwY6K
Ede7lXuve5qs3DyzT5KczJuh+V5+NNFUTxxOdQkl0TY/NO+c/99Z3p7msH5aFcSKDQWq5yUr7nt7
Gxzw0pm54WrS5gmdpXBcKqQxVrBHvt9faoGVjzHOaxPufBal+aYUo5A/MNri7dYDIPibFVLQdZ3b
gFhTzMJ828KvrOp1RTqTKDmCkZY5ByxX/pcKkGuQHtzBQIJNgjwZDyFG3C1QpH5QoIujANzWo0Zv
Z4Azlh0HtdRheAyM++iIJokRqsaqoCLCeyADaAKHcbU/T6NwHATUncjgKF5uWQtek536TfFyr5ry
m2z8gu3081d9cqgSs9k8YmpJgChKMK/MrpYuScc5PjWB1sUZXhRIZbziApkFQuB4sJ17BLD5JT69
9ILLzCK3wXqvlXM+/0kUdovvvFqOq++vDifqgjaZBdc5LXRKzOy0yH8ZxcKzaX+8A2MPPFVY3Nbf
ZfLUdfcRzWtq0IGNTRdMH52INOvL1DuPo9hnVIq5yUGnEzHR6nRHzRUdRaAqGjaCdRxDx1z5EmQZ
MAPEofxyyk3Obml93Zc3Gp5cTlUGM9VS/nlmbInlRz56nrv/lhEG5QEbwWOpomGkf8/zvCdrMMA7
NS1Mlgmdps07v3Gp/auYnSThPa6tjH4XrWcjvVvt9/imDAXFTWvjTfzociHSW44Wl5EsuWfVSyKz
AaEUsVMuzT3vnLRaZr1vigTJUQsySy8k1f2d68r4WsL/sdJS5tzwjbxSxvgdxBBBNcOQYgf4T4GI
WYRLtxVa09FOesvaC05BQiLDcie8UzqVCbD6dAZPIpsYuP5Gg1+FyzRaRDEpUJOoGL8y4OzUR2xP
Vq/g3Vo36s5QREjA3WagwYI2lOMAheXWI5MIKDsG2Vr2rZyPnxG/ERsjEBFhBnqM/H1fnnlcTw8v
DsT6hpwkeu+pHDZZ8KjYKPfdt9r8vAGF4+DqwR9QuJHQH5kWemIZKKRIQsmt4ZFh7NKaLJfLAx+O
8LkC6JsU8XkAGOlAvrg4YMX+XDwl7uyJsDfPuKN9EWARSwkHELj4oDrPiswdVWawrtB7HzLCqExD
04k1g/9Lbmj70WFjtqWYchNXXQ1jg9NTUSxbjhdewEo3X6SNvdKOgpoASGKIjsmLDrP65KYFDlMa
qaE3eJ0K5c/IcOMt28q0zWBIyX0vcz+9KhPZNMaOR8UCL0VX0MO5IkylJbypPRpkU4dKX/IiHwD+
E40srIvuIu14xTGeGXETGJDITWjgK6bJdAGl9QvpeX7m43Z5ckIUzMEeG8m9uscOdT/9hV4xeRy8
RmYaB4OMOKAuBLW0elojBT6eu511yjCiV4/Ps8vrP8laSmS/3pzmwrbhnXuaVspV1XvVvxgWIBjP
sWwIHAx3mkDbi1cJoua0Ak5XZdrLjhwGAGrZWZ9cZGtveA6ECNttmwaJZoKhGCmv2Pn+LKWZQxyq
AFK8xoqpEk4csK3SX3f+sp/7BRU20WEhagtFBVZoTJPZXCjmqGkeU0rUysivmweDT/w+SrSuSIlO
p4D62Fe5th6WYouNN2ZJPegn2wKQEoKjQ4jxC3YdrVLM8xisFoLRn9B9FpPiVVtQaN0Y85pt29fz
sgKkj6GHUdyNn+YDwJlSXs+zy1TyGho4SSqdZUHB/jVS+Kw+spmuKC135jmKE89hjdMLI+Ah3Cci
7D4DOWPxPF0jdLQfxIkC4jUKZ/YXU2JT3RQsrQC7kJGuG0VTrd31j3/AdGsjfFiinTAJzNb2+/Lr
KKsEFGeoG59dwIfN1xv8RX9v9WDih/i+rlL8VW7VWZim/MuUUEnfj2fFHz/zqnSsEXZARLlNBGWQ
4jQeKmJa9UA3b+INmuhiy0nRgR5Vk45z8bQQxt4JCrzFy0wuFyKwvKB6z9UsgwLxlWl/1tmsZygo
Gzxk4vIeM3wcIpQM9CcGlpPw7oHw/DxAC6NlKJ1nvU6L/XaU9xgmYPhRzM9sI73w4cgl+J5Jchb5
c83TAie6tE4TAyHjN3zy18CFGS/Ie+NWVA2MmDHlPp/SjilunjbI29c3pOPxNv6j3U6T0mRjJD52
oAfP3iD2wNTDosM9pba9N73huqJOiEYo4Bh7xyJlnBT3plHFzRnev2MCm3YyqTSmr9H5OYAU8uYo
j1No3j/x7YXMzA1gQVxtU3ys9x2vi8KfZn8KdoVpsvYK/vs/0mK+6+E12fx0x4XckFEKYUsufDWS
CG8FpDv0tle3KmlL5KeJOnuQ3pB6GIuCL7Kg359ltD+yiziDwBto26WRfovgXQZv3UXrYKcGrot0
wNqoHZsjWqZlQK7np7ZXJW2lFVPMfyOCrwyOUC59puFPjDFP8z3g4IHHhhKZLFFji2eihRqGIq4+
TlIm298yjg7derPqJKbeH7t9blgEp/7nKz1CDvWDQ4vutVhY5kM0eQRzQcN2ZqmltmJ+BCKfT8Uc
mrj+8p0Ptle1EdWhcf6g1YPCoJ2DGC7ne+V0wrSobeWr4dUsqvy+yIbcRjg/9lk+hMWez36dyVz+
I2Lf+xAy045oGdynJwTmxIU7D+pzn3YZ0adHJ2lbdVUb8MRqIwJqJrW5u6RN2mDZ+h5DY33YfRFU
TvIzF33KzWanUv9NVW6OKuN29MONOElWX+Rp95dfVyF+IhgEMzUFXKekIGM6gAT7fnWIsUusIowL
wtQndD4JuaqHBHOjSDxCmIicfmS0OJgD6yAJYMYmR29jyUfFXibx/IoqswD+zWXivdZjrMi6SNkG
CYi2tbeCRuTkW32FJD6w+VAifFLFRNjcqnSoQnJx/+H53doFhKL0AVqRskrmCz/iPm83BZXEA6a3
33gmPjTLcqEhbxVFVQ2euFk5bT/RB+wgHIucW+SqnBdiQ/1l/WdwNGQSPDoSvAyvc/lbV5I3xuG6
WC4kMHYqzNaZzo8etfMspP7rxLbCe0CVaxi6Wv5k+WFxIyCaNT9CoqNy8bq2LoEZSaljsG7x8TSg
m92pRMDvX3kKrPR+1I+SXKac2R5y98mcwWj0XiWGsvD0Fv8Su1Mfw/Uh7GWpeij3vRN2I99BvL6U
qe9xJk2yFIACOTSVsShA+nSePmxmGBga8i8ce0Nt4Q7DyKClKH6sK/V4QjVqtAwAmYkDMR3KODTL
Fo/ZabxOlAQjIBkXD4evbzrBWbyUUVIxVha8qz87BBaasqYeNCmcPJKL3k3s2nHqVQzDpJjJkjzl
eRJ3umNy9mRaWjc4EIWsKmqMjb3YxVEmGsGvuBizPNUM9l+YS+6xHn71htKJPe7XjEzPKNvOfl63
XXut0/GCQLmk4HN3phOBFQtOf5DK4F5Ed02irw2eSsOgQRaw2vaYZsxkSrmiYPg7Jpv5ADyFIKMY
RbpeAOj+d7VUnRe2O6WzGAe1OZDBPq9Vvidqs3U0URyNFR3y1k+4zIiU5zxJ6KjYjNa+HpIbdhG2
5NwIo7H1rHUXUWjPjct7XeOOvb0DmV3/+8x0B46LrH3f11m/NZAGpGBJnBJOmsHUG1ebcJboIVfM
JGgGxeq9c1ZF8Reid2sq8FXBy+Yaf8PvoX84js4J6E0k1zgFw5YYYFUrcnD28/NpawMx1O7NAKxc
HAM8ZEIJsGSHMlaZF+2Z8rNaXLsMSMsaqSyojEsmCFJLecHs8DPS0q+9qvMsffYItVTYIbG8wP66
PiotdugTw8xzAgH1RbD7rkCs1QMYHqkIqt+VfzF6Cp8ShCDmWdbEooSjjs5iFViSEcDeha39XLvn
jMSJYTa4dxQTCAsAEUgchW5Ihja0bK/3Ndrufmk5hHnfmzjxjkVuo1PGpk60zPNQRjzt+Sjy+3+s
NlPxZIt63GSeaLSopgFdK53NmEtN4Po/Gf6OLDhY58EaNpxUStbQJAE73jLx67NxsQsGV0zBAPa8
+dQFglvrvtsnI+FY5IQ1JgDnw2gtBa0xGfvqspfQt2KNVw7HvW7o4jQL2FhZWLwAq2NdICkTmHLV
IVff2vjST7QD4C8aBWQHxvhVBqTfRwNDM2LeoAsy7l/PEqLa52T2HyqprfuEkXdfq6u8lMALSWyz
bYzbIUJkGGEeRX2RQNSalSiPrdpKKJ2eNcgFhqB7NGDNFIo6ZeVaaomCGLoxwLxd2pT9wI7gAyfn
JwRo/cyk0/gGfrbQMhK5uZ+YptQZQSKjxY6NZEE9AzEa/wEjHwhmVuLsod2goG0Oy6h5Om9rreZJ
2VwV2bRWbi0az68KQdfMyRpU6++CVXICJCtcXs6nHNJ55jMBQjNdhj4SpT31Wm3Yn9Z4ppU3MIZW
XhAICFntV/vokzqoRb/GvknF62CGnY2E2gb22Fg7Jagiu66hryXhHG1cbiMVDGWyGVCCiB0zvl+s
sQZCfiKD+qUVCdIh1wfzp8TfCdldfDqftFA7IAlADdOZROHnj9cFgJ9CDD263JhNTJRske4qP8qk
LNPo2O8F9wsWVCzKSf8xooYf+g9oI/BPDo4+pBH35Pn13p/dkkCgvgOUwllmEk5OiFPD8vC3r3jo
hVF3wwJ1OrmAbQdb9VFUy3vJqGAoanY0227kObkiojNotR+U7TYpbNxF86PeCwtF6eAuYkpPbhJm
L9EeeOV8xBtZ43FaiU7uMvRY4y5t0eZJXAq3D2qtpt6qvtO9wrzYw6ufcrpW+Z1QoLZh2VLx4TW6
pXC1tfzMP/B4EbLaCUwXU4CaW4vyw5BxNv2DQWAANnJFcrZ8KJIZJpZ/kZYUuk2aDo/gtwJXKTIx
WduWWuai5v8H53WopNe6TQ5DexB7xVdymOVs+tLjus4f4P8iCMioePHCX+hfKp1+HIjkM0cM85ul
W2wdylJSbMREpwuKjJNwrOoM1Aqnq5cg6EuZREFdxYrn0fBWB0rCCwxvGgmvOemDH8q2Rx2sAQc/
i2JlqDkjK4L4q2dtorVvfbVCddWOMii5tNmehzp794luCWP4OntZ3alt/tbMRD95AuQCMzA+/kyF
o7BSxPLFHfx6oJMZB/q8V4qVXFTVqq+d++CA9IelTY04tn8Hrb8elSQQ+ZRSxlPdSW/+aLRtNuA+
BtD7YNNIA8Mk1jFbsKP9wge7av32t03XZq/pVpjXYdqy71Zpjd75QSymNwiZUtTTWb/6YFOI9Y9w
SnGbAbm7dopmSwkdyFf+DrNOB2dGBYOAOyfC3Sso0s5LvSTV++J93S1jChYtmPWZR7J0h+UfHfBh
L/NqMRAItQUFiJEWVYQvdfc5O1WitGNDwi6xoTLtVQl5u7Ch8K2Fe7MlyqoQelq6gVmCs+twAitV
tJ8lKYeY6R7jwAcLn5QtzHosCBjIB1rBeVUZljS1ZUkonYLUB/oub89nPEYy3IkF3/X5S6rdsAFf
Y8V/Fr06ZWTd5O7dMVzj/RwbsLJaq0Uh5pH8Vkti1RKfEPy0mqZjLd+viaVxHM7+mbPv2+H9qWsx
Y7sQjC+5ZG4fYFd6P2IZTnewQEp1AxcMwrdTz2+r8zHkhg9ZihFWY5a8fANQH4C6qV11AD3WbMfZ
my7/8BbAfYivB39mW2NUrcv4yvrhQKsDUog5h+wbBtxRtIgBaTKY/Vln/yf6vg7nynF0/3sEhRNX
9p/g6WQGXWyzvEhQ5vTtc2palhx8GS8fuzcMyPhbwNZx3jmDZxsLmnYlui60mAupx2Ws410wYZJz
B7yRT7dTaGawKVEgce9T4Fvd7ztNeRqBqZelN2qWgDW/gVb12AZgL7R8TTtrwQtpN6sk3q8PS6o3
cqDOZvGthr7Vw3MNcgM1/XNJFNLa58st5I0kAcJK50K0DtmIkL08FEU49+h5/LVqP18kW7FAFzLr
2u5F0D/a7EzcX9LkDObHufTZzTUOscKBVoLJH3TrxvGeQCuEqzw5CcsSn1EosCL2WBI8+AO6DGKA
2k7vwewjSlSemk5Zq8vq3XhU24ZQhSEWTWVPSdCkqYK4tMIc21VY0DHXMNdG5MrJNi3LoT94LOlU
GFUw54Gw/g4XACAXBDLGXXxKdcGCWms78wUunTyKu+nR7twu7AmWjSXITRp4mJh5FcEnLaweBJD8
heto2qEE6YVD2LkMpci1eKlXBjKq8UQofBO0tudY4h9WZLz+oWYKQkOJwp5m1mEyJRnAy9McYx00
6ZKoU+Pb3SWwxzrXhkHi6+pfcWK6i9bMjkXKFM95H2WIPNe7shQETSFjK9gz/vSN8/wvGV84fGRh
aBx+fRCnIKK46KnKP9cEN0bi+5TvLasa67wCGk6jp5yQ2QH5DyXE/bEPqpvPIuT8YTcRr2xAKM24
C7UQ/cUUXT9fiYuqo+P5Se4FN6m4bEy1XSzwH+voORsEs7HbcfitnkhiNnS3R8+H2PpDSZ7UPpyT
aIrlsxBOJ9OU5u6goYABneP4eEa1z1NEP3qngOCheoGSVBB/Kze11BEriDJ34+5YqC+Uq3f6twjC
gyoxiAg9j/6dZIOpVqSiW4QiBdX2c/Ed+Np5IVcyFXZZwLoOZuo5vRqPHlU8MTJ6dQ/NhYf1s8Sr
uoTmBQeavwxqqE/Tq82J42mp040fjiWbL4KTi+BTpwXyOhDWsM2wuuUVtuWxWiaswwpqH372gn+s
f8lnGH1bBHS8kmkPM8SZZPS/+HaEEBga+wmLgcwK3fgN8lAQ3SiMGyy3gB5/Dx7D5OegvLGgYbHp
CQxU0sERpJ7cA6YVil3GFuax6BGxhYYzh/8G/7wOyNyCG/OARg9/VmK24b/EMzJKI30cEDDokWOs
d6APMJkeveZ2By/BcUGJNQrCTqZDDDKNrU1+IqaN9rnZgDD/ReNy7kvBW85qV+HVeQzJbRP4ANDr
NhdlmRW/0Ibay/HQTQnMxUv8FMgxzNdfh/D5EpcN/h+6M6dOnwSa+GPlhNI9286Z7AAucIGAWwxl
X9p4+aIpq9X7Zvd57rqkvbUX7mKm9xfuZ6plgiL/NL3mCxRBk7x0f/NQT0vgZSh0hiiNCCRL0Uw+
DOVYSLDrhsQ97yrd8XlQitBk6ynxOvD9yUq3hr1EVq3NFsoiC207z7S9Yf3eITNzGd3wwf0LbmD3
1ESKoNFTpVGIVGgS9wwM6otf00Bl+pGEm2bTUztbS0j/hiSbyVWb82u2wgadUUXxXAniL6ZEtLaG
Srusd4x+O/1KHS6Eca30O+PKI8SMUeGgVWVFNgZs9RH/2vf9doBNCZsLzt8+XB0BDV2nirrMJhGj
tyr0nbKSUGFlPXGqIYT+cJluf3QrUJ/ZdQT43tZwWmA3IxX9xJqIuYx+zmA7vhh5F12BlF+0y2y/
L27P2MKtQAsdF9a9rk8cNktSauVG3Aq6+ywR60hRSrHnUyy45I5SZdWPkhEZiPtvNOmdxFOhQZoX
2qN+jlF89k9TWhRSCoQwmi4o7sH8vEocs69CZ8IPwhTr2Jm5qvsGoFmtKmwqC0Ws0slFLbEvP/BC
ON9g4DcZOjGaKH9UL9HD8OP0PlpO5HaycB+GtVerm4CURAVxmvLmFxEDDiKt5CPF4Hll2ND+mX57
oa2YFU0FmNJjHufTk+pVjhq+wJSIBLRROrY1fI/Pv+8sN90qoaq/RSBX1V6bvdHpupCYBHHvn3ho
0vk43nvDCWUP/ENV35jfnNW+z48KllqPvbZ/lvmDwxMmPPGxNdtQVD1mSzd+8kgt3vsIt8AUjIOB
ApnMrqK6VF7F8o1LWRLmF7zV2YNnKBIBmbjG8pDzSmLqsU5noLryrNtFNNVaTPw7d0kDcnmc9v5u
QHc2QgPLoHuyrPv4ILv0BLeApPdU3/iJfqCqvqRWSEs/IIeiri1alavAKXUDrBHwoX13DZ9a6jB5
HIlqkNcUA9e1q2rPmjkYSIFQAe4MKysLyTbE9V7YlALImZzBWpPM3aP/glW1eN73fG67Gh+nD1cB
xhoq7RYU/v7X5GX/MZV5Wluikptw6BjT5G8lHdOAJoGpMHuecmcXEaWFn9+EVKtyAYfnjpGCR3H2
s68qSNry8LSwvB66X5WjTHkZyjueUv+0N6tnk4J4tI54g97sNSPVnI1Lxk6+/rNeDSI4cLEYA2W4
dMn1VZtNmzPLn0jN6TJX7EWMKyAgDGCTB8b4WgplYBA/TYDG09VEZkqDq5IW88jAdwB105ZVlVnj
q0EJcu8Dq6ZCaQL4i5WLZ4mv/X+6tdsfk8sgw5cXLPJ1cwfWLUJpbZeKtvAAWxPCWNxaP++o73w+
4T7kbn2OcF3JkSIoKJhCUx0PZ4OgqKlBGLdC9u4BbaxnfRtkc8vtttP/P9t39Spd/XzuCpkBB+in
WvJrBnGPhbAnsCKeDbkt9mcT0iVhk47VbHJbXhG65GQG0Z2XjSqHNO3CPLGrhZn1iON/7XLM3Kvo
gz6hxv0KdE3r1xUhBSlCEz7DkLvBoBT1jtNDWkmfgXEn/vfsAlrelTycS6h/uCVqnD7/QHN+uY3I
ySIsP4eg1DGEH2qj7phapc5Rz1tMRxkDMfTHpRo3sKHYRxRtaqH1vokgBt2938HWELf8BZ3r8Cpi
WGFhy88f1jryRs6bULfYN4Ga8mrxrJsHjmwqyhAdrk9+9Lq8Gq9WcDBn28xZSM/s4MC0CWXGPxDZ
1/w2Uw00oxF5+yoVLI+3WB8OM08XCYToCKvm8ANzCRUYNJ0cRcfz2pZZhFlzAuXApK5HftvJMzBr
5/V0R3bD/qP//KuoZba28Zm3Dd1a8D6s+Lvs2HKTJ4BVyfyZbfrYJHwNPYQDPD0bCFGLZZM22s1x
VZvToQQJ6gn0X02ZHTNWzlqo2ADg25FwKXeHR6OCXzwkBk1kXS7D/ZYdZXyfHLob/HXjISL/d2A/
iDCzfuq1YRvDVjyrXKFsxMSjuUCzR8+J9sxha2K8o6Ovag5cPNw9BAbUsI2Y7M7dHMjzYzVk9/jJ
DRWjA/DFgDZoDYtc1KOHhipSzyBkml7j3qq4dDTMl2VWPFG+3s1mHQSm6rWeeJuxMbNTmEf8UEsv
mRyNDfAfbjRFX3f10pTZlNPUikC8Jd40LPh0DB6EJBNE0jcD8Ys3XvqrrxPU6kzx7XPNdwpcw//p
4nfe/ctLPpFDfGLiUVBRQED+BT0WOr0akjiTT8J39+fQhE/sgh3da8g65I3gdpDfrjsmOzNRSyMk
4i/MuaSz0E8WLfmFlfaUsXAQxTNNSbUizNX/tA6NdgYzzw+LzeKMBQYuLPVIfWdrlx7L8tzyQVan
Od8gjf/4QSyP5NRrt9gdOpBvuJmirhlStFMzfe2/E7hHSZ11IFgrgqIc0ovCsj1rE5BtSVup09Hc
Jus7arWUEs/uF99eVNoDWql9JVsQ+wQEc5fN+YJDe1z10SVjBPHxjakG6GdX3GaEGKodsi80oesr
ECB8BQ1OFdxcyMzkdM4PAT9qrfce5xlxyFmGmIVzgNz5MjHNqXKSEaje3HIwualjpZosB7VIha9Y
45/qtZ2hgz0WUtIDw1PwqodtoN92enbBE4gQs3gkKTQYAX4Qkbuv65ITDL3gzyRA5mnJvHdwwvem
TezLLdr09oIwYSZIzylhSgzFC7b6acniwHcLnorDkpx59qm8vHzmAbL9BFQYd4955OwKcUFEH9Lh
1up3Al37XSgjVWNq6t2gcMaCARqpT9O+fLMmFr93Esp1SVEZZUNKsu7/s3Nki9bWUesssk5FYD4P
pE7W+f0aW6/pWa9x9yZuLu2fS9sNXWRXSbOOv5t5HShEdEDxUUR17sMrYpoKC73RPNDf/1+nYxhL
RUvQuF9xdec8KO4H6GuOnlcmwYS4vkR97P3lhEsUvwYLLClUgLYYWW0XUsvS9sWDlHZWJD0R/clZ
Ytg6zrG+8ejNdruJkDeFU3NDIBGh61X963+YOTKB1rwhG1x5pq44+pFKbxbn7FOBz2OhNSsfxYoP
iemDJCQtPhrfU3W/l5Jeu3scdPJtQQ1+/VPm9OvK/HOQIDEVsahVIAJMo3luBqgYpp56/rek1q6Q
qYgtHhy9Jmcbzu3MxifnGo3vpNrEz9VFGmPbog32NK0dyLwMRb+Sh6/HK6hjguAjUXc8VpZ2jhFE
ABdRJCAehlsD0zoiwM64PaAcUxgSNvz/D6nY6wZRO8WgGWPJWRK6E0bWlIp8gQYeQQAdk6EQEvqm
Q0wgq8YhECCfp6ExuizXMqmYjusm4yVktgZPgvXMx5WvPLlxa438X0M+NOIyCRWIwRj57FqeJw3k
ujTxcKMRhCpd/F//lvDWM41+DebHgYh5bBHjf/d48nCozYzDtwa5N6W/eNWrgTDpTp92EeWVZ1ej
DbIP7x/dUcssK7jsFUJ9MhKlr9irW7A1J2qAl/DAW+aqy53O/O/thERGCcUnyYMowWMpw718VkSX
IlWG75PcWCsTllaDUI+BdNSPR1OrRDG1I1VvdVWmSIdjxZTn7opJywvarMCiM3Voq5ecl/Vu12sG
ylnckbJ/OwzpZd0AZHrY6Jq7hNkmaTZYT+Z047I2ofr4Uw1Fi/iMqJh18NId22LcZYMXmYDtEiBw
jv/FcrP1AiLX9Qo62jDk0bxir+hR4tb958LBguw/C1pWqHuzQ/a1YfiMwuhfYllY/Fd90HmCWeJr
8h484XMBU0HgfmNDk2gsFhHckJTiQdWscuo5urvlQuTzlF5BRbpCH9e8m6EdQZbbLtMylO4H3UaC
z5+JnnjWSqQ7MrlE2yhglzYehJ8/dLigFtb7rcL3nfpoz/vriIlMbqKuHHDvOBZHUNjhcom+Exwn
051aqRsqGRz5HeBbXstMzm5LiR7UXx+IuhGCg5lzJti4cUEPWM316vAPVm4fGjDfiagKw0ePbqS2
t7h3j/rVoLGJJdMIp5IC3zq4HTek3TDUq7NNCtmbLmkEkS/cryOc3zJBLPBjLCptW3ye1ttcopkd
H4XjMn1XXJ9yK35Ic6mhtjBNuPGnS1aw9CF0CxinNmTrID06KlnNggv4SLmDm/BWZfTK9rsYFlL6
FJhaoG0VSR7pVIS8W4c51jpSChI6OPqsGFJSkJt1Be5plzq74Wghi9n2JQ6RYpfDcbgONP05ykCF
Mskq9AJn7igUnNxjbP+Jh1/WOLC04WSEj4y4XVqvbPoNjQvKBETFQPlP3R9neaL99hZkMuLxmV9p
soKVAWXvSacqjCdy8630y4zKNNOS5/JQhX9V8A+Tpc28vhQg4QtV0ZXujGV9202rsJYxdPngDFpc
pXV1AuXPAnRQWcVhMN8kiDh1akwAbieTJ/dMnRTKeXJV1ua6cz/iMLpBPgSTx/VN78KVqjufPApR
6pUJ6F2kY0rFllSSlisMPKCAO0A+PzcDtHGZ4xbo9sdeJqqPHxSGU9X+rqnamsZ110e7tzM8510J
YNCLnE20QNOqLxod5uEJGLXdaHgGVF1HC80g+sxeCOhT3W9MlFIELlQh5Qe1zjEaQmAVt/JMm1f3
XIGSJJTQxOJSNcw8sxE3lO+mdicAxEcH+GZPzAsbuNHn/7PMBHudrV85lwIWoF0in40XoYmLUpUR
i47liI9CG1DrZiCfkzlRQpEv9JrAUS/Sq+uV440V17r5XyimwfDcrJdXm9JCcEr4a0G59ywIauxt
DkPdlvh/68k5c6G/sdkeY98eRJJ5wHYEpnUFb9ebU6NAexP3+ykiWJ3SGvVo5Bj+vHzt/grHDmLS
6+qFxvlhevtxOEvzb96oSq/VdZOvhTkAL12QPksWxqQ/7Mx9e72268i4z0MJH3/Rs9/2dPQn3NvH
i8N3ZTvuhcooIHMD5NmFXlJ7l9PEmKSePSL+aiX9Br/EWeEwIDf/P/qR66YvIOsr/FRsF2DQu+2B
PUYAEBgZAzqvqReYsZoFKzxIptk2SwM/nTp8lwcwOleQfQ8QQZWcoS9wXRbgHr44GEe/ml35WeXz
CVs5Skpu85MzFfO9k32dKafO4x5n1dbRAWkMmJvod6x8RPSSPX0EvoiZqwGydLo3ia194HXpe6wf
yjhiFrizluSs1GaSgHjX1Az7K1lhTu26oOGrzkES5h/aC6rus1+iWzl7/eBxgOnIpdpI34HgPuFb
mpwjNf+XsmH0JfP1h2t+KvvU1vu6Wr3KhCqm9Nz8erdtUrnOVOzqYfx3phxtjOuQNjPrenQT6GT/
FcW+IyZYp92fJd+Wznc+5YspQg3Hw/DvgviYEVJyGU2CkSN1V7BOMztbi4nlIS45TuLlyPLWHHSM
dgysdM0F4uMXGy8TC3dCmR1TleoEHaMGthGE5UMLrVMhaPekA51wPRL6jf63V2ZH2mQURxZ7JDua
lbQDHuthZO5ytnbVOZJbeNBK5bMGNFhDkLk+tDepLOFgBICaZ9sTEuZv3s6kr1b1rTLYv8c0S71b
XLyBN4zMu79f8a2wplcfHG2ZeZ5U9rcQi4w9t54lArjLQGzXX0DYy5zGf2h8gbfqUujMUn17gaxy
eXm8/KLMl5JVKvfFZgJ2dC3WNSwaXBmOThoKY8PU1QjB9SzRTkHhyTL0CzOdDgE5ZFvNrAGtJo1H
+W9Rle75pj1+QS6Bnj0m8C4uw8py1kpdDbnO0VJO65onU0UdQCGyy9f87nCloxx7HYbZHZE3cXh6
dc8uoRKlBjBXcBvlQzyluoVGcjc2x2J94mwlv2KlM17k0PH/dcmTrjJk64uobz3+SmLm5Lzfa2pG
mvK6qvkewZ1q8s8gmGJzWp/aL1xZdFQEtih+mwhhpZ3yIhJ3nH1OdMSJVVy76C9V/mgsumrI0SP3
Zgw0Pgmia/SGmiexIBaIprbC72KhrnRGW7aR7G+AEDxgzHz1LwGLSVeut7CE5T7NMnKaPFXX/Elg
Y38vUVMliWh85NEK5fRPgSCasSYf8KHvVSw4sHNYzgL4BQw3NDXH/oTkPf+eOW6/5KTTqj8Zmhpd
ZY7W3mqcDBmd4OkoM3HC5Bc+Ebn9NZLSZhR6hqL8+juf3MY3KmmmI6I4M+8GmWqPa2HCybwPOHKC
oQTDltHMjTHdZr39YTOVwwIQv6e1M0qc2d2wG+oInJNaCfzqTDoE06783Gkiow9g6LLZA7dhUgy7
99cZ/nTuTNuBEo8J3owgi2wd+rbtlMncfmPCqHPEcW2S1+410x9/z5YewrRDtwTGRwMJD8NVJj1i
AgyOh2MPPO/6w8LYlkYV4uxYHBI9Rj83Q5/AOEu32NwpIWbc2NtZlXCZIbgQjYE6ppxoc1zzXYlv
XONuqR6L30FGjZAUjcUYD+aMgrwIx+65BUPQyjMIBujAr+cflxO3YSOgbAi6QL3sruRg6EEE+cZE
DTHcjvqPZWEusBiYUASWMDuXE7EF/1aSgY9VUE3vIHgT3cdvn08GKbCLlFifjbBx5ccSZu+GwYP6
Eb/hvedBoOkzy3wze6yC0ArGSmWxqjQB3xVst4Lxl1annHvxAju35inFBw3Yab2r/DLX+YSMgUYE
6jQX0tzytLgZpfR7wHqWjo7saIpneyesVfUOUIoaWouLhteQ18FtH4eIlYuqMtie51k8IgqaHtrJ
X+8jSKDvcpBhszjp+N+78ygyraw8TSszQAKM2zi3gWNC6Hd82MdDj/rqh1SVYmsqCmexXSrGqs7g
VY1kNEWu7IeIi29I/HbA7RRm6kWUayFcgTvkusZjdNLnixbErkqd7oR+JbJkn/WgyBX9AdUOgXqP
FnabPRsNfBeziGuzdDhMa6dzYOiIC20T0M9NNbDra6TiHXmubfMieJls5eYt8snGXdb4YQPncOZL
WX0kGVad0NRuLfbOLnlYhJtIBQUzjx7QDtC+HewsqWdev68aSiJgoEby88dB7p2UO5pJSL+EgPMv
yKi9ZoJlDNohJr+2ZMr9cUqxxl3+kEZscBNNpcapEwwBrOHzM8koFg6hgVje1FCwap+/ABOMvAfi
4LgVNm5jhxc1gOt8Wx1G2rAF+ffZ48q1JHzIiIduiQx1wf+LowxreHSQXXCoEALAVK83YtL2BE2F
E6sCL50CF7piNO0S8OPghGF7ltBdATYCL/pOSBvj/LsfVwVF0yBJsh/8OTW549b1eqzMC95TtxwZ
moV7ibYLVEJSu2HP6NztbHX7JsGBMZgDH5Pkv+oQCder84xM/h9QNfj9/WuvMT3Pns1+tS4zjWZA
5zX4nf1NbK5GYSpXebR6imW561doLgM59j8NO0SGTJJUzkVDpZdhMNxztjr++mSWVmFfFt1qH45Z
ZVUQ05Jc9r6R/TOktJrngwkW+zW39QCPt1EBfxAk+oNtYP0PlXGBA/obDZ9Nv/X3RRNamqlIl1j4
oN9Ll4NCHBbpWFmO3bd7NMDQ4JzmWj+IRnBW9qMGGpkTqkLhItcUiRApIsvt0Z4Jb5esHcSiEY3a
e4At1JsdQlwO6GezzCeIEvFnCQIEJYZEq3L7UOX6raxZwPUDsUsNJsHGWN/Cosyif9fxL88+1Xma
xwV1OB5v2J6rwsI6dvczEBlruD7ZHsF4A0pvZv6VaIAjRscA8oehHYvFLDEkvC0YqGkSPX0RkYOp
fI0q/vwnZW0+EgUiuwnI0bl0x0SbgxJcOWz7AQwG83wsEFOlPkxRW5gbCAT/BfXyBocUnJutAQ8h
hjpp3WaIBfCmT3Y0qx11D73ly90XZ+CQ1X6XcP7ZIfL0HlTDryThjpIYnUTaQMsQnTUzs8A1MfYw
NRovTYbllPPghuGLxP3AVrbBLVttp9BQUJYSb9pS+ahipNACZQTfomfwcKrbwZvtjaOBRYeTfMF4
Rk49ifCusrdfUppWHUPO0TEQO6aSVb9mfoafxq5r1T9dG2QG5sB1sUFUkcIaEXNiR02hqNMznAh/
eRv6EVERpiMNxGBt2o7WUCW4AqJ3FBIIRWPPusn9M3t/lQF0ND+/gOFYvJUO9KXl5rqOONPNhWad
54SG4ULBb4/LUjGo459MK0mQn2dE64tDdCO/gUT6RwIqQpYm8Mr196tnEiK87bd1myc7lQh4uT6p
hSxOAYS3X1v3nXpONZlb5ni6gLO3KoBrwlb0IZZmNC7uOvKPeoIwpV7pDgTEcNSxYCZZNo8zPFxC
PHxkJL9ocJtZlacipi+5OEFl60MEG5hjPY+HWJa52ohGs/MgZSAVpDRIxMqTVWSpRcmxMHOnZ4lo
Q/uiUWueb3P89b3EL6w+wk9vW0Yhs6GDPkJvhNyXEED/61BIIvOmME5NU2RpFjitR7xJc0KHvB2v
7ZnEhT+MexWREn1gV4UJatRMoqede4eo6NZCweeKnsit+P1GHLvLBBPmrM7y4Os7JIjW/ahU48tY
K8F/Y2lySwtdcOBENE+gjQC+Wg5WxQd1sWhSLgRVOxF9TbV6rQs/Xa783U6J04mIFP99F28dK9Gt
1ig5DGVZ9rHbGNyecNf1Sa8gWLFlFIraBlBua+99mhni66wlpFCKJmByy9aj9KQgCF7kKXdbLo2N
5gcdDv9blzSVutXQZuinNgWADSvpsb/5sEmflysKch+ezAvOaQ6UgtSixT6usKjsotnrCFzCuDKP
3WoZn5XuefZVxmoC3cWxTxwDNI4BnWmVZASp46Vy64I3GJwm1jaroDk95MrWuws3rB+wP329vxiH
xQYqM1+7kGJi8kHuFDIXm+1qfc01737mocw7n+9artI5i7MK4UXES7UweGvzyiyoa0m4i6Q91vKw
lmrTjWSjF0bgFPG7rlA0qPbfnDWqKTcQqxoEA5q6kaXWWR+qv9YEW3CH/LghPt86QuA0tjhawi+z
ab9Plyv+EuyIAvxhMG382gbm+3Y4W+ow3jA6Lljt5qLp0QZHKiXxmhCIaFR5Y/KHht1evkfLH0hy
sMr4o4xBZZkXDct2o94+hTiu23EauqY+ZfYaMqW+cIWHyErXyWqX4lcu/wPPwCNnFdwYFxs/pAVs
pN4VcLAw7ngx9TSeGOLCNCRq2CLvQb8kGmgroxBCc1DO4IrbsKyRUnOFWPvZwLTY0LZCSk1MDssJ
jSyzGd27YTyfdjUlCjvM04J+RD3zeUE1olxpTzHBTnVmbwer0doLLNBmMFC1XhIXLRDsYo4s16Hj
o4B+nMLijGaeBE32dcHUrHHKa/+jgFDVybTuorbyE8o2i8bFkoUfWzxnwhzIjsgZFZDW1zShsty6
RPqrh4KRjRe25XfOSCAA/eCr7kIwWeLNrNAUzmT1yQQbvc4FGZu2R0y5vNGmo4jj9Zu9KGgQOtKa
zB/IwCTAL7B32/y4iZgUbO4hYVR/0UgbmaIDcNStO9ozOr+59/vVd/v/Lt7ESMiIfKLlrobdK6Jt
wOEeES4oObOzEawsQVz2wPNa2aRdAXWt5DBwHAzJSmuXQWg1tdplhx3uyCrjWM3e982VQl5Wb0jJ
6Dz9xAyLm03DsUC0q/qXAmWc7MRvZWVWyuwsk2joMZpXpCI++IERwQmk84F+Y0ZBlC11ijqyomLp
brv3w8XN+RouvRqEtYBec4h1HtORTzxEFrTkUi/HclaXW5TJILXmrDO9VvRgRbj4NHkiXNCyZHL+
13ZsygXa9wltoNDcuv+HNhSxxdBtcWlYeTecH3rTE34b9UMMne8WUapeHU4bRFCXv2fyFuuN9aVG
hGXz/Jk+DYm4R2MnOYfUe4BeJIF3FTywo4BKWKuVo0/L5XRhnIpPKSCVqyJYSrcUdVUqqPVCGp0g
Kkt6gDdtB1Wasvle8NCcfzRKHKaLQhPTksrTx40zdghjNzoo2OaeS7FyBLvPA+Uyp2qwFpDsDN1g
A/h621sZKzlfN20ZnTk8rmxCKLvjxsViFSiywsVaLgaAmvzbDovhGfat3NKo7FtVDHw5vANoCzJj
EIwsEeT/NX7hF0cbaKYDUSY7bqVwGHR1R8sTEJ2TLZ2XpSXkIBaKroGSLdhnnqUBbUvPyKJy7l7t
O44Bd6lTDAVep8Fbji1bXy4MUfZmQGqu6LPSNGJ2CbnQod6vqIgnueMIp9JKW3+mbEZfJ3Futb5R
Upxt+R1EmAhKOpBDMDA18ZqJ62ybiU66x1SJ/a18xPlqy1bTWn8RCxFz/3dSGMg5JGjIia0JbRI3
gCw31aQUagAqdUt8Pws9xGKIAWdTATlKCSATjgYws4iY39t5S0Q6FDR7chCx1axZi3BoBR9bI6Lw
x1h9sSTvMHKANw1IFI9ZQ7Y8X5uHrJU7UrRvDNQFibkljMiJVXph61qnpvcV/BcmLmztoJYZFbsv
xxAOmbNh3CaZ20jNQFzfx0a+RYvL19I7OsjGQgwA9Mm4EPB1QlNWPIRm0zhrsI31/MCrCjcu4NBY
ozOv1aNsN3SJWKYdL7S6NRdO2XMXOiQ/Bt600k1PmGZQOFGN2bNNKdeXUShjsixCTkDQXwX1BW4i
Xk5fXDdGsensHiSSbFsEkkSd/9bE1fomYz/Uojstw7sYh6iuqY3JaoTtrOMBRnyll6otpgbkwTt6
O9lTMYAEiDPhZjJxv5VrAPy9a5U1n5k2DMT9aFxn2sLSoXIb+SowF2cjXuYandQVFD9CD+QPJU8j
jcLy1L5cdcPLs5JNb+2BxwAEmArrnaA3CUDcs63tkh+mbCZdDo96wE11oYgyQnVbMFOg8Diz/Obx
muk5AaRfJDMTSwNGCen4Dj6R773foFR9eVXTETeKfNE6mvbnpZPcWhBhJKrUDvERzJ36j2vrBgYu
hekyaeJWkZQvc3SWVwjZSYMtM2qr5T1UE4y01/GiWG5t0EH7CcggtUIdWJOsqa0T1HbY1pbzGfXL
E4J83fWXQz5Lv0qkOm6imyHNLSffv+99xa7oY8n0r1PkH2i1JQXlQ30sXcGY4tcr4RNsPGHfn9Us
z1T8KLZHKFjmfNxXKqXHjGUu7OTt/tr2+YPvvdsNLeZcoP1VQ5ew4pDC7JDympFT30kqwIN4Awjd
7qchXosB59/shpJUu9qwRAA7NhVN7G3h8EsQXGZFgVs87HoutVjIdeztgqNvbTyZQYjrQIfQ8Bik
X2KTTPPqmzOxI7JRfwSVNgwewuAGmhTdzXE4XZIcVKZQxMeDMYMeT0y4S1XsQIZm5tYcXoSFXlKf
hDmWV4T/EK+sIHGWUE105VT8StmcICMho7ckdXX8rbikX9TCDMrBDjBQZgTGo8Of0w5Rn8ikM90v
DBg9CVTRmM8DdMPm3aSTywYH5LM/UcQpt1+gayfi7yrYqDTYDz1ACXMBDhTebKxOOLE54IJfWqo+
PO1uR4vz3e1K9LZyEvFnWM5IUmvPnGkptvNe9lSGfrJBqoKDKAW1iZqSVTuU/KETL0HxxO2GH/xe
z2ZOyzT1+pcylJSTHu2xaNA25fV9CyQPTofM8xyk9Fnr3vzYrAo/4oKxbrGeftXkGVdh9OS0zIl1
p/Ex59qZAM8qYEjcrI/yzJ0/8Eq6BR6t1Gn9WDinVs8Tv6Ara23js1VK6DZhzwbNFWrNEUPrMyTW
Olrpa61xRc0GUlUZB4GPSSCHtON8vwNEhN7790JMucrL7XQJ4SQEt1tTXXk/h/PKNbinOvX4zWq1
0mgV8/uSbnn44jPun45FEnet44GB3iXmO5qRd2LMSgWXkziXxWZbQLHPD2al+6CLMWq957E1XfVa
uV3FpTYtutEojlPKHUUE57Ggr5KIzbqPGbY0d5pMahRTs5s93VKZyf4BSeaeYYAjoNWk8+Hlb/sP
TAPFdFGxAUv+yBMBG2TSG9/mZEEs5OnC9/qBqNx5rewWZauPEpB919yX0qb5EjVBPDrmr5AWq+zd
tk9QngdRIpugh/+V5m9emq/rXYq/o2GKn6PB7X3Ka5JrKM/hlv/w1D9MRMHB16AzRBD4dO6kHwp5
3ibyxkf8FvdLexmuxHCWLeGJ2cOyDgrMOtlNf3KNYwB4eVWp3BC0aL3exHpifQjEh5bjlFAniHkX
udm08XHNvJhGRxN1w04YDfeWjGqZ5NYA9aDwfGNvKNxrAkjeWiUboudbrbZLOlnAfZPSOj4VIvpx
3zSVj6lSc4jIND9Tvvr5OJBjil9f8/No/UM+wh2OWaIt8sf4X3/0LU/S37xKDfocdpy3rzG1i2D2
K1ljnDNifAh3vMBZlB42afjov9xr/PjOJF6dFYCF2nLNO+oZfsN2Ys8iFi2pGQSj1C1qfrCLw8h6
L7jQiyRn7+Md5uPnl0Sf9Ap1kmHhUhchcvFT42xitEQySZVJW8hgtcw5LJNBixcbONdXQHz2t5aH
dbIkFtvo23GjUAiq361+IbTQY8eLt0ccqy+L/UzIJFsXoq8oQOXkPtRk1JLZ7tqVniwwVRb/ZEdX
mKDcqIL4k9I/+i0TgqGP+zhq1nUe05lxF4ziNa6mkD5PEuUyqY6aJ3LJddVs9rq6t6YDC03/AX9M
tIDxEorb+OTTxMhK/yds0a9U2PSQNaMUzbaD74yLY7bvAap4FLir4VptB1oH3iLTp5It+Q0gvoUZ
oR6z7A5j89HRFODNH/g8WSsrCLADwH+1iW+EaGwol/+JN62/4eEw3CI8EREsbPlZez9wOINKDeCo
mnkseXd94WJQVXBt30roQeDyCbGR2deuQPc5QclVNWWH/Zl9kbhDR6c+SjXK2Kp/QArAqGCfh5y6
G/75pmQXbC/saBBqPUPVDjVfWGHowtWt2L9gk8Yk7JCh70Oxi0QMpZa0gwSUXpKKLypiFfD0nwv+
XnEcSxuNPF4Pta5srso2IyEI6AcZcbpZu8GdEYGaKuOgABEI9ZEvloX+H0b47LjhteXsMkxOllgq
5PFdnJ6ghJSGJ3nDI0epTc6EEIhkI1WqNUMO8sfu0oVBdBiLFmRcteerz+RGA1wxhJPPK5iSOumN
Au9RA4RI3P3ta5MzF6fdUCFl7N61hroIxiitKDsA/w/wiro8Q3jSlvXDbLym6chKJaan7cWjHC7S
mkyoFa5IDt6+El+KMILt9hIMcG4vFZG7wk1oEQBgC4bxqJJIibFhpKXmKaBOCWlIlzzYtDN2MIsO
iuZ0VeYQTwkWmzuQpPgPWOmgSTAhGM69xa0nNKbyk3cfAztYvywkM2QlDOC1NXw7iDzDaQ0xsa3Z
mXIpRtpkuO69K8k4wZJwa9c4bugweLDSBajUcPLv8FC2Zaa/9eYbdav7IPyFYFBDGtYH3ysSmJBf
lU+0L5Vd3bMhG0EDbmCgowavvHPGiSSeZv+HECTsXXAOh0KpTodIf2RXIuttOcnrbyoNSruPYjyy
FR+GC7r+5rkrsBR6ugL+uHU0FtUROn7c73j6RQDP9Q180B+iEcMIOer20+iPr7S8JqPqCwfi5oJt
B6f6XlDY5eh6pJkfHz3bfEHF+nn96RN3/SY/7/AkRTS/3M21IYYskZ1GNS/4qrcI7YhCBIy8Xlts
N1o4dWlXkx33vegrgPNabaEl7v2tjMaQJEeOtAirTRXhJjWMElOy1qxxDgqkWnAsSN8vdaJFybGi
V4ejYrGF59fXKgXU7B39MJjH9RiTk58zv5Rt3yhtIdAN+eJh7721X2ijjbNQ/O6LQMJXkanA9tb2
MRoypZ32IFVzpsFOXR0EgBRykmLrsyDv7OuPTUQThfpnsyNgqUPjtuzdi2+zCtumyscBQzA3w1PB
6rrCGiAkV+udSLvAeADOViJm5KxozYXxgfnCsjCFH6gNx0f5txEPyOpLbh/JKK2zYo0kFLTdaLpy
4nB09Mh/Ld9IBcsAKhZ0xYGV716Y22twbE7vbuGNGwCjx+WsYwXXRJ5eG1lYuR6FPwymJOVwtNfp
hEMUJjYkPXL0AACt2xbaCnviJVKnaxR04P7+5RkAJlWr8IOjnfux8b828szmJpr2dLiTPAplKYFy
N0IpaljUjjIdKMo/Za3QSLJZmMMk9ShWPNr5dppQRCZl+FiupNMWmxRkpJNKs6t/UCMPgaTRd55X
EEF3OSPCMvgVLJzFrk3+EgUbqe5sipMeYx0/Mk2CzXgfjKvFjOYUF55b9XloOthAdVs31YFEPTMT
GaGzotc9fTZ5YKPCbJUg5ByWNWYh+V1tPdFmnXzYus+L66bdR+ljIk+pElvzoYPwjGmU2DQmAhEr
mfKvLgQt+TCWlY4iGaHF27gaR93BTrzVjAxdk2psOL0vCjgYxp3a36dmGsGOTfbCt+JS68+O7EuX
fPG8FWZwn1P37LqCl2G2KAPVZj+Z7I2Wp8smFljI5LYEpL59kGb8pR/vf7B317CUzLd1OhiCwJbs
oatd/8ezxXavrNjpn9QisO1iejAbNuDQNUgjf/Dl1bXEMfvdMSig2l7wjOQnMqUJo9Xvmz1TrPOg
vToO1Qug9PKkb6wxPj14CJJf3ruXMPsz3FHDtUzmm0dHkkVES/bO59yYt/zsNMp6h7CHhGZDqZXX
wkrpckTlatK9tgQ7jIsOF+yOIVeh9mp/AIsSOBDGNehq3mA5Xk5DpBNPJuboehXt924Nj8OhhUWl
tmwmgGWuZ03KMrxff29wzZvvvHAKk8V6eZEwOqVGj4E4hVQcPxSikD6fcf4L7JvUbp7Ob02/oEdN
h+kWlvGlOv6ORnsvIhdHXJAGfN10s20f3jh05iaoO779K42s3BfPMhR9QH/Z0i8o2+UhaUMHrAFh
xRSBRKFsRHDL2xwGJQSMYLg68qmmbcFNHZLYX2I00dW/OH9MjSSZPNX++WeqzmkQq2ezRfPywxN1
gF1zYEji3BCu18zmOWiStjlMLtLAABe8fAeNjqCL6dfOEE9+HhKgBw5WL4yC1IjerAo9BceNvaWd
q6u/3v2zrV5tBlQgcBMuqiLclZLTPvd7RzZsQQS9MIfSvTSP8Sp7FUx5OLiCuSjil8ADVVyq4V2X
YxKGPoB7gTnooLZRe0vEEkoU/VUE8jIURvnDSD8sNZHk6JPCkaf6L/jt3zz3c+VxS4WNRkzaQew8
owufWHVDiHwbQT2kVYocHTSvVd0DD1QvQuhbveWBRH9mDpmj83qskv+O5JkTeQdbLz9ScbnznEd7
FVDoBUv1B0fK7eNtL9iQb+BiYMYnuyTW6dY7EhQwJ7x6WtUqJDmZdl0M+Fi35GhG0FgSb8K4uBKa
KbKKQbKBz0xFttMTnBUkHdCL6kj7ONjWCkH7NLcdk+KB0bvdocf2Lqe6tCYMHthqBd+EcukR7HBM
grX55Pk43vH0l5pdIgmbN0Xrwa2kj6ueHd9FT9/B0abkqdaedU93fqDBbYE/zHNMqCMU6s9uUhFe
4h7lyWq8X30rUYovSQqdyyOdpjQeFSrTnEWlPGlapKiIo7zyrniBIyKi2C7znOgssDDBFP/54/Bm
bSk6ZXhYvgHru+BtUFAuidtATyYXNGam+Urb0Y0tgoKTVyoi6eUURAYlSAmTt2lbuS+Ppr4L3FOY
mxm2fGcZlv9meT4wv6id0+YHsQLCGQMh0TeNV6AUhj/dlb9EwSDX3XYGWfbSGJYeeNP4DnSP56gw
ywMcLuf9sSxU/CRoU3H0dpwAQ7smWdlEv3nc7kbHZuEz3cQvvz9B4XXsNk/6G8uU7Q4zA9zdGu0d
9iymr3kfUlXJg8qBwMFw49G01QgdpxKHO+buQKQVGatxC3TZQ7BOxPnRamtlsRecV3xpKttg/zGe
5QHLDFJo3PSYABezbKcEEe3UT4r2Yx72O9jw+5H+lTmIkg5XlKB9TLhDxb+is/P4oVqNOBHQVDzc
AWojbLvS7jrnOQZokp6s7UEq4q8/QSGTQ4+Rsq9NLbL/+0LdytAHrLDzRy2Okb8TpmdA6MzMqam1
iNvm+bYzmSRG4+MRuQE+zzBSGo2ZzN/8zdAuJyp89UJA561vg8Ntc+A1ztUTazAOglR5dBXVf59o
K8c4pwWai6yZOlWWGq66j5Fdojr4NO9obiN3gIMscW5xYl7U1VsRrNnz4W2mFqBoq4wNmTh3KIxT
GNvSWAlQVzxB2FEBCzhGBLZxcT01QC7ejyPFwfVtQRZny/bM66GGU5iJpqq8TH2IFpd0tys/rAH3
B3/6qG2zRnPqFYhzzZ1sWz6b39Zsns4TVaHzB+vJWo/Bbft4JfIL0U/Vr7Mdmp1hn9Q6z1GzuUde
KInyBJqzXj1V4zkNXmd1MivO52pwQ8PCvD5dhhB97JCm8auxlv4utmq50THK4x4qWTJ3g2WVbF6U
6l05eOOpst0/rFxbzuKGayvR5/mYoD8Qnf0LgvWgdeOh7yOjpSTYw/0W7t5FcPXAjHuchFZc4Z7q
3d5ALL7kqvahes215jr4U7YQvZ3Fh8zB1PeM3my4JsYwfVeXrxo/113LborgKjewoutZSSSM5cMV
FvWekryuDP2wv6sliyobYMXRcKWNqijOp23z+fL8YgCV1f4H+s/kDILtHYhAFKMUunan5/fXOnFB
qC3gU35+hP4c4oI2RMcuvkNQYoCOfn6XLs3STnuq0CP6I9ZYAOJSvc4Va3Tb1OLWGEtY7X9ANcS/
J6S3YBuGN8u0pEqb6JW76RBo0Fc2gQdIMWs2605V/WZvjKSjx47/TA8LRljM0580LTD17wwj45Wt
BQiQOCS2nWsycO6Jx5BPf67jB68ws8JrOSikOLLcxIlVOBqZZynQSwUSy2U6ifwOOBcqRbC4XOLn
PMRXsmuClxrhWIw8vLbDjsFNpRzplQe8N2azfeI9hVQzaN4pPsjwGznhz9zIlzq+0yXoJgL8sC6w
tGwtR/9Oa2GoMF2pi855Q3Lre7frtRJSErBlPTuzwrsmPrNnEvAq1mHQeP7ozWjciumW8xzQioCv
9VELQo3JSdmdfqOipi9iEPkIWohK8c+GFt8rMAbBXUl83MxKyawp6hO483zgn0CH5DE4SGfuGaXt
T7gYqJKBhlWowNVMMWBZJ2UVa9o3VlcQv+Vv+cto6AwKOWXqn+xKPxk4dWQsZMqR+0hhn8s8coPb
F9DTL9lf4RQgka737cy6UZdFTgNpprJM53ZEdMthCkDZvA3GCayijPFwMpS11ON4tJZC3Evwu55q
Vr9nKu25EcU0ra2grEvHLrBc8tOLtft7AYbKGCkhCxbbeHY3bvx39DU4TmCS3U34IhOJiuL+YhYN
vgg9znlw9mPvp4DcfZhl4HUdh/fmK1nOnhkhYgFtWkI0tUFzWsaGprD+3N/ml+z1oxvieECYf+T4
9wueGNeuKr4BLthhUm6VfWiEz8wScgL2rAJG4CSqq8GFmf6v84Up/1DOV5HBxXnMs0FeecMRXlL3
Tm5WMXNaQ9XS1biuXsI44Gz5/jyfQOqXy3gDBnkl2mUwDbTRIIz57OUFYYytiA9BuG6mSa7l0ZXU
mCwnbUR7B8biwfH0LoUFKt1m61nWth2298JjnnlA2C3nzu1kubhxt2UzTmS8RH7Go67f/R4OFACq
eFYLvS05WQJJT/E32hyuHRxSiz/z053JDwru/q4YZZCtN0f8xBrez4Qx2g7P3Yv2r36nbXW0tA6g
mgxtvdrCUi48epcM7oD/vr94ucEBUZate05wMGJ5lpeci6aRa/2EDslZBwABQEXb+DmqQOMaLKeA
MZUmpk6CMGj79BhxsB29tjwR16wZpbH/Da6vbY7j+KVIfC1W1PR+9sDFAUjVKjN13vIHMmVIzKxy
16J1MAZVTitAvlqD6pvwejnlLvhr1z7StHQdwCrTxZtv56F/ljSbA9WpZ3BQYriffKRF+vtuqlBT
BhQ6VvUw0ZKTf5ekZUQ1uyZuAMOoVPm+u5QcWIs5DZaYyggEDa49QYOTxS8lDInw3T8g/tAubGRf
hC2PPvTaRqc+jLFSrJN/ewUx9/IQ4a7h2F0VFSB0uEaj53FGRKXIHgLU+/d0qbeH8MDdJYc1XT7A
CVxJ8cyL9bVMQd8M2t+AtP1wOG9x4UHAlJH4e637ZQ9H0y5oXX/fp0OjQpLWdkd6lQn6TA1cjXsm
m+5xrxyxtaWFQeEsuBgIZipaFL3jWq2XCa640oTr/AcVp+9isTTJsOXoP/E5F7K5+DEkdrqmpF9/
jG+QcmYKq8vTL682rSMdc/VRBZ7BfidCfW1uss/1iDs9LdyYGNtEo3tHE+DjNCJAhx/HOLQAOFxE
MXgyL2StPfHoXcRZRGI+5orLHWhYrReHz0Ko9lqKj3qi5f9SaM6YIS7UJdbaJRuEOMJilFDLXstm
J86KgBAjbS56OaX0htT8FkpeZ36U3B0iLz2Xi2ghvLg64/KaMbqUQgL0Y7oc/MS+pAIrwejhrqZY
SJ1mPqYF5lwQizTEEXPE/ugrgEp5R4XCf+hQQGAhdpIo23Y48/LWs6xlVDFnw+eKeKXd7GErF0cA
sy7I/dvXpfJwYiEHUhIa9inGDrMsTfuAgvGVFscqsh/+Ju8sncYyhDOPVmjfexHTtKf4UDOuSsoY
Yb7u+k+Ds5QtHNUYWEbYZg+oZcQhE96dZfgfsnrHjtI+jXtvrN36IOqdVs9hkMtq0aMm+3GdnYfA
Bf8/cmv/tjq9w4lj6Nh4SnX4IbB2aIgmChD7QzglJ0MwAcqf8hKbayGADsFAT1PebvJWaRB79F3r
N+v72/wbaXfcbq4ghK/OzvXQitWfi/VU/V1tftPGRIHQ++TDQAFbSdtgzsla2G9Z/Wzw1X4DKoy6
HXJBjeQGvnN2P22/kNS2BDRHeNiIBbhEi8/W21ic/1MI9RuyIX+NJrJkjD62rievSqGoNvZqxbpb
rqJLYiQFocJ2XyhzRyfn0J4jWHjKuhPQG0Tcz2ry65h6qjsGf1oqDA/RqyXemYypU4T7QzEsH9RA
UZdiFiOVA3MJHsT9er5DoDA5ZoHi+a5ZJRjGEK1N2aXsu+mnTn4fAZS7LqrCtsoRMsuTytggN74q
ijB+m8a9u3Q+N3Bz1BMxClSL2zJBgqfq68LnoyVp0xolOMaJpD3rthgUNhzJlHNteVyrdiwVEnqS
1ZF/MYdlUoe6H1Y2r736YS14Mi58VcLroM+2RJXvJo/nNoeWy0gIQFHzl9hnGNHhqSWZR3iZYJ9o
3Mg1jmhw4QypBbqknYpAPDpqhBtvaoL7zws8on6jb1M42kAQ6l49Mx6vinTENr+c2iB1TUzAf8K5
T9SHnXaNDK0Okty61LEmncCOES70dZLISzdZs9hMdCINBTDTBbDd6IRArUsTc8JLmiaQZPJL0s+U
13IaAUZ9m5pPeDO5wwysecfkAb9/V/YyELPMBXQXaxl1HoOqj33U+bj6NFaXc2D3sV72riJhdNxs
/2gh3kgV//Jf3v/nELvPtxrOulDrf50EmrarEzr4AIiJxtiMRpHeUM+40ihSDO/BtEu5x2Zd05Ae
Msf9ft7uSOcyJodsOERLZ9IuNWfWl3X5BKyWNI8AjANp6WaX+RHRflXNlTob1l0seMdAGL2H3Yjj
+hS5qY3Co8sqR0XNS3WdFc+yrVU8IpyUAN2akvDflkFnGnJQPv4qg6fyPDaCquFU8J7Z5/phcTGX
cG8d/ImCqZAeiOr8toizjudHWWi2nZM1TCmD2C0zITrb6Xmu5ys50G63dBG4XGzVJyHjIteLZ8Cp
pLghte+swaP8xY8VM+DCzJttYzMMPg1gEYJdbBEsaAByNKGj6y7kDWsymSqHBUmebTWMuCM7jsEK
cEpLq/pbdyN7jTNT6xsT+BOU/z+HzBZOPOWdyrKotSJZlaxv1qAFY2AQtdxNwrNyz0/a/DQaO2yj
pquvkKUhAkOfDESTCETXjV1uxjJ34LLNLdpRU/bA8hRvxFWsuptO4J7m8OXkFJt/zYFXOaD8klPC
h4VdVnhGuamxyc1YHPPvUjffr/E1ENSpBb46Htvj6V8bWJYsTfcI1HgPpBav2r6c8hHc/58v80gO
9o0Slr/y0s8R2curjSwJqEaOiin9+8W3gCDLmwsSmFVJVpGix/GOxGZa78k2yW1IzW/R/8zSJ15W
a+aSXKybPS+DmeOhSNqXXcuJjOurGV+5642G4imf5GN9EVf/Wuc+QbBK+1+rMvWbxWC5Yc2YGKf6
WHC1RZis71l7bDZYoMzgX7GPADgVNKTUGgj45W1KcWqpmA4rRRXsGpwlW1S9mSN6QGlKe5RIOWr/
SjjtHcoJFCXu4f0qvrZesJB1DRUFFuw+XQ/jqqzkeVehJTy8V27b6QWLo8/TnaBBlRR1U2KVR9DC
3iL4w7s42P8rYbuITw4s5lg3QsPYyJfSInwcHxRNV3u4qAmvirWwrfoYdR3IvECV/VygTPNRVrbu
P+XrOsYIfcve3VGHD5Oppucfp1phMbMyIPocVPFAcdY3EKWvx5zVjwBqKBHGQOYEO11z80DigTyS
0htaX9dOw09Lfp2DM3+uhum4WInjToiUtEcrLRtFTYz5FbYXwvnGKNuGaKgybMd29/aeCpEiuGu9
iCna3Fb2NPaMV4Wn9q3dXy4Dq/nj9IArHCZwluNvdjWGWKpP3Dc735qEJdifNbgUj056TB8K7VhI
wMlSGeCn4WQXBw4Nm/bx+LbsRtIKaB/ZUW/uqM/0wxx6KOuOZjR8Fh925NGXMS3DqH4nGh5dDFOG
TSsPyWfwv9Jn5mLwHcERx+BWjuklVaovyqLy7uSfPiT6lVp/OhfcxGmUYZPKUBx23hyg8Lzc45RM
P7ONoEaYeGG2E0hac/2jfexR9vSzJrkHI30N81uPXmwVydUZZJi3GwxLvqzo317V1UDRNP6G2ZH4
/wFXGmJB2sTH1OcZJsjPHTYkP9ZYPMG7GKD7Pt2agdPtZa0DvJMWuWk+Ru75SrFtxHhcl3gwITpJ
SSL4VF3qzIBI6RA3jtHBgfvh4HRIhwOqanFTnh3W0VZJQ3h8AiYwvGafVGlnkql9RCvcBsqecHye
TkzeiLpnD+uVfvheQAzfXwymLCDr4aiXiequdYXkEewj0QzUzjthf3mx4INiw8ZmVeNnmyOZTd7y
Gyb1lnxmy2d3zAuumgcYhuxo/G6aSgGhTvW740sXARo/7kis9Gv1tQA/eUpqqPOcg71MjNwu01AE
rshMhaaYKu9IUmSNHHn+ABDB+IUu0z1tPGB3RHO0vnlzcWOi03DWVPKcC9uuat5ILSaKEZVhWdT7
pFMqAipSGDjMKX1Dyb2kw5cx4Pqbpv1EUEgeOp07LhJFqg6ZxOUgF77Dn+sn/g7XI0JNDqTR0xFM
+Ql9Am0625hLzOLnIDZHqVkCNguuLPFj/ytpuqQ2I6ezONKGbxw5QjMQ7U9C9GWtlw+5+RuFA9bS
osdWK/ZhWOotFWQo8kgSHfFgzirrsw/OVLZowWsQIO4dbmMY57e3RsY452ZBnN4lsjrM+ZZp/mDq
7L7/sTz/M6dyZGHvkUFn96uH0sxkub6g9HBh9Ua8NKEw6/ahK8oW1bXgiMQzE29undK+qyXSwdRq
kk1hAt75Pjgb8Tx/jncIrv4cWpx+IP15vw8UC6g16qv6T7X6bi8RPo+f068HryLxfB5UQN5rDsbS
cgF9TK9VSIYVb4QLBe1ftKB1YABj3KIwaFsynMMnW+BahjXu9eloruyS1iU8W9y/omWoXdLd09XV
pqXJEOZnlgsWvdvO/uMS54FkscVhf2PIxc1WAigRnmDTJUluLMR/Sc1d/o89UIMqvpbEaNstA9jJ
szwkBTN5V3nJIIdO11aY8l019Aa66mM5bHXIuNO8RMtroSbSusxy06CeLrWFu+2k3PK5H1SHo/s3
eQ5iEeIONcYcmC9dAqVQp2+aKWQcazE1Lz/kVAjr+Qem1h3W3Q6twDv3LbdTMOT9RNllKYSKwHv+
AkLpabjBtkMvM5StUdNMKMLCmRNtUFr/ycayiuBNauWxLxNJuH8fharRRCRX56k+7qI8JjIEkXB5
CmUTkJ9k3InHGKa9SyTAWV//pZtPOkzdVG4iSME7a5a3hJW2Ifc4sn548nYep2nhwKd9zPc0RaOk
bttFtUGCVvjqtCDdR/GPngGxMvEWOuJcA7QSyikeqQ8fRiRxj6pfJ/EpWvO6fKoogFqa98H3/PhX
68s2LtiQz3APV/D1JaOsEsxEFW1CI0e295MxysgirMo0w32vPMkKQQTlZC0EeiITjSvBVswwoker
8+PPWdB4ortft1eICWSRnyhft9fCbdIE/NM2vjaJ2aYDleyZ3vISGch8AM+jC0bZB+pVdMImsYkT
zujwO4gKCelmjvG2tRsg9PCv9pTQsznKcDvwIUSDo5un5rzPVvw8vZUxnP4t3pkByI5skESW6x7d
/qArc4W1u/T5zO9T2UXNe4Kh+D99a0XkkZ+R8R7O/8sEN0vNTEsVSt4gFhvKvFHGccP7DRjU52zi
iI7gkjM6qKK1ol3TpJADYaW9hzq0fLlek7fuO5uf+unEJ1gGKacJnEuDCn8daxxi8JWsrle2hZac
jNE3AEd1SYlEh9AkQ4KfTrlju2U34k3slwhJhoGZeOU2ahnNyFL66iyf0eOvNjLuHiZhPo47VrhJ
7KpZWVW79bbC7NMYbptxNv2Rnx+gP2HoS68qB0TMhiYtZrU+fOODsWhH4Cq+H2Dm8hsPHBaZ9+dC
jFWXLlVyoTgCALRNAn48aJLw/6vOe/jYJXGmvNF25z8iKh/4tQ4LUwkX7jdx1Envj3rrcm6/2nHe
t8vEAZIKjZSi0GPPPQm4u4OJmvJ1DlxMcNyneSRCMYUGz+rlFG8DedaULEa16ASXbsAtBcoHUqld
7SJ03lJDGK2C0MuC+wHIQOmgjSj6e0jsoqAEZKVrd0CNHJ5byIC6CWpVbgKcRTp222/9Mrzmfo70
XDMbfT6kCOSKzZ88h6fv3MUDXc8ySAUjIrt0xJSbm0TtsdoejRnpd1Nrl1yRFR7qWnxh3C8Vm3Y1
Q4IFUuQbUtfJSl8hkTIhS6bI+upPqx3S6CKa3FB9fRUj/Phrw9yP9uQ4cggbACyTnfsVfijvoxP9
xqfwOjWwDBidUnDMy84jF5ZjxjnI8rl+wwqgyyiiQ/oXT/04oso65LJkjRALdAuuHi1Pf1KaHqay
W1zPRNAGZc01CFKqFGvSsWTcfCrsU5ociQV3yfOpCI66urzYWsOytIhVgR+sP9QNSNxUpMTNwlC0
QtFbCCpayMyieomor6FIKVsHYmXzXmqd9lQwleSeEFTNKajL0KCohWXM2q64y6oBVcrOU2Ftqx4R
MQ7Jw3RRPFwX82FZl3b1dZ/hncQ1FLLww0HC7a4Xm28xTLhM23N5HiY3FuBRweNpFjxX009fjZZv
Q8e4voFreUhYBeFPT+iKkWVokKAJT4qn+WwwsYrG6Er4qPV6xwylMXTVpkApgrATsThgxVjDSBTC
HM+HwfdECHgopeQOleY1/rIv8f+naxGbaZ76S5FPrzgdi16WpEsGc/+QvQ0ERP5/Vk3RC1nBjY4w
JMfOa2nc+nJBxx7W4U16cd1gbVxg/fhfNUq61fvULI6jpwNNhnRCY04LS9k7OiV+DjYHdc2f47+e
SHMZkkIHovtCGnzr6eRvFS2edowTXTYuK2b4jSIzqlELynd+k6H4AyHUGZ2789jGmxU9I5/0Ocu2
2PZbsqag7F2EPx9DOEJUFrqeQyCwW5RkT7BFIvSMU6kkW/fsbvjMUFwjTsWG7mOEu+7PHi5a0IAz
moP3hn9AzNBXZE5MDYv/XU8wThDNqYheJ8L5EzQ8aDzU6UkCShaiBIvsr0Lbh+sA4/PqwtbSWZVe
Dd/jmA6bN3an0kGRW3KyIaGowFvXHiPRUvPa66qB0Ofok55lBZMgIoyedwBUTMa7zJ+Sc9QxlLCI
Ojkq2gYIfMgEejhBeTcnEky7lLFblmmsFQ22uujo2Jvrg/3gZptPtnLhJfRXwmA8G41FOXWjBXLo
e0xCoxgHAN0ATaM/nPq+TofAblvdusegjV3982WDKTCTgFSbfJwX2bqrH3XgyBfxI7UsjU/g7Hmt
QzvliaH70V7lBggm5VH4vL3BnbgtgWu+weWkvPbDRqTKvW8ukJwEP0Pee33H+INaxcH28+gAPRM9
XsAsU2n/hThaMpwcpArP6HUjlKFYJfWkFASLlWCyhssltKjnJCI/MCGrIcNk8ZgZSW6v6ZrjIFsR
jyAqYE83/Q4UfzUpkTNIB/96Q88eA3C/8A/mAEUkM73wntIbj6pQhzggaedMW+EL756TfhWR06c9
9zkE0hDGa1FPhL99Y9RvDsf8O5lRnJj7jsoBnUTncLWHcQlh1VQuc9AKD1HlpX6BtpakWcEQOZMI
oxNt3Yp69xo/DC9mggg8VGxQZpGB1L+c7Vk7BEH3p/8dOrss52DdomjIihlZXZWn65WB1S642Uqz
pjIWMkVEDMNqe351Gi+OhrtW+VdKVYNMAXhAjC61cJ47H3LdT996z+J6y/qRvFc/nEe3TdM/+K50
SLMZ8Mk5ew9MvE1HgWzpvweRW33k3FQUJH7Dym8HHv+FuEIsKcLRJN/S4ZJZDwD/vtuYkHSklJqi
3jK3G2hLT29pcMK2bbpP2HDPrxBz4hDvqmEna51iWUzaoYzvxrjSdTL4YrfgGC1/VpwkHz5DFPLL
qL8dFFU+fUJIJ7ngcU3YhNA2ixmJ7ygBKgq2JH4lLHF5Y9U0/ToAq4NJeuokC1BunNJbzxaRHAiD
l5hnIQzdh4ywynYo5f7xT8yh8aoMibpWDPKfjp+et5Tlsd29Cxlz6hvtOhotwDsT66Xf+fUJ/EAW
38CLjSacZ227mCp/v66Hq1QJpM35yMOz/KiBImd6xV0SWcEgvIpJvcF7nOlj/uMyyGmNNKPfplcE
XVH7MjKnr57lFpXPOLnHPDd/UcmYR9ZIzn4N6dNSeS4xHEWdDxF1Z55eFZ5ZL8jn1whRrIn95Gq3
t9wrqIoHhwj97N7VCFstQxkaJ2kPnPFqk/cqKWZHLt51dwTs5mFpZWFioMWdTPb2cQOSGlTqpfir
mRdzyElqNjeU6e/XWzrIzDiQR/dHM77pTk/tXvALSqzRs63ly7K7UrVEssr1CUlNO3z/8hVYdGRZ
vgmJsPPNJeTXjEtPSg65nN00PLaDinvzPr4xUWF5rEdf25gsmC5kDVjXGAqGrOULoEDQ/eJLsPM6
iUJG4/0B3zZCO++vOs/npsATXCUeAdDdY6HaVm3WUb5fs1uBQp23zPwW5dvnd3tyCGJNekSLAIhL
hfL4oaZzSxUXeYNPHg2raLi9L8X3eKMdlPylUr04DTsFsRN9lKFOsrr1lBRbxi0/7HXYeEXHeToS
Wv+AiB8k8Sb3ycciZkLJ8u/uYjiPjtsi9e/gV3aWj+zNteud6sNV1Sut0PF3t0a0Oo/nGJi5F7Je
9QtXXgyjVRC7DU/iEUrKQmpZIVdLoUFfwkM+powZQoZC1KLXJUOXonVXOWzR/0j8BYel6U+tJJ3i
MruNrH46QZHOCVcufH8Iwk4+1io1Q3tPLRQnrHBC5pEls2kNrAOKC/tfA35gvDpazLrQ3MKD8sNF
IihydPVKVmPP/UFQIJDfyuUs/wHhazXiT8j5k+AZx3D06YUTpt0MxxRmJu/yMI12SnUJnkGk9fOH
d/Qr7DfVls9MUirsIHn6Q4HOqXiiG/zMiAtKJ6lr6JudKoYOtmytPmPGnI2eyID1an5+7A7IJ7yZ
EEm5DooNZ2FcGEGXWKqM9RsvKQEb74GPFYfDt73GNWsmbz4/elNkmYs4+9459lEQVirDlpjnUO0f
nkcNgdlCWZ+EEJsN4CoB+7C3GF5FRxu5/9uRsD1zq4z8C5Imu+Id+OdqKEozwcAZQ+mz1ebPLCbR
jLv4Btcw5ySUMn4EdbamT2h8sqievBPWPGl9nFKJR3QMWMDCaWmn77TnamXbplpSQIc5ViJjt/H+
44/uyyRKZEhLtBkgwf+DpKjabxW3+fEX70eh8EhySdKbmf7S3muoureuK5/CGqJuEN//i/d28Vdl
0MU/poBOft7ixWZCoUyIlXyyfgNGDSpRL5pMHrfSMAUkO9mVhcVx5PY1kkBh9ysehG1saoPsAcfT
ESVBZCd0owxyTHX3+RmlcRUXR94T8/aqLr6f1H2iL3jloOwLkaITqXxa952rVu++039fy3N7BTso
YEaRK8AehYrJI0mhcNRnKVs2B5dk1Xzac7TGduXhe4ReVGPHxkwrnYZdyonIw7YcwzoQrfk79Az8
LDHWqOQfrQW1rTi0axca/Y77+kWTANH1nOTW1rgxYuqQGgGY2RiOz/HiF9p7G8LFeS+FngWbQ1/e
4pudR6x48tKctGBXlRtbtyJSq5A2bhZ9g9RGP3YuxPUgwUaL6xFWlyq8KVRHC0Xk9gXac76Vd3+J
C2M6MDnanyIpML3YyJpS9Lf8QtNDPTq1E1h/P+E+Pi5098LBs0A2xvNd+MkdeRmgkMPC9yEHhwR5
dlNf30QXvdAXR7nsdD1gAM9v0uFfEkxfyyEEevIBIDWavajSgnxys39FiGOOr/gYhva3QeMXkuE0
BFPCBIT7g2pEz87H/kzW1zMWaAuZT3ImD/1wanLTxBfUT4DSIKzVdXoyZDv4F25p8kmpfmb1x2Ee
ClSz7RofqtBrapkDVC1UXJopACpIderllbL525KstgKQrh+yIuPf9TYuYZ7cea7yLT1C2xX4q61+
gZh8sTWeXO/wrBzM49O2D5kc4/rscSSBybwQeIdUnL26ROF9VwOUOYt7f+e6ckQyB7iwgIrnvrQU
i+oIh9Vn5WlBrQf3zCQSSi1XtqUEREExKY4p1tBYs9Qi3R6t2bL37sUXIGn4t/vkMngqqzw13UQG
NlZgPimYEX5STPB5QOrlppmHPY6Lc4D0lHKjqCynH+gBOemJNzr+rLq0IF7RxnyXhMaYQOSw8Pa+
yPf26ckdocMQQ8g2mKnu+4pZZn0uW0yoQ9p1xeaW9m9oA6u4m9k0oTtslco9XgUMQWKSVcwK59G3
dOzSZ2iVHFLxKKA7Mo/H3xljri0CIyiZNH/k8Hoc1RIWojUoBkeJYmDh/ZJhywSC0GGKtBK6Pee/
wWC6DKN8sUx/Ljze5WlLHXLF/ZAkLizn0nLvvvjRrBJUX/EyI+EvecEOHsclzrt85Kgt+N01/7pp
WRHYpA4503JV1LuEAcQ46pXNkpZV3oBTSkTEIciRMnKcJCoF20SYPHklQaDjA5reqrVtywTyYXIM
skogoEffKnK3sreerD/XkQIYBaL6J83xbyko6ZjXM7Z8DJeBn0I5834MCZUGpB5fWenXxc4iMl6m
7V59HETmEWg70z/xND4q43p9y/u3JV0+sckh79fmVQfYp8BYHajvKAzTlfk5LgmJgO40Vs9OwoSJ
rRbZaDYeKx0mTHAH843plE168d1Mb8XT49WQllZKpyTvfmOq+34HmCTEnfwpBW2Bn3enXpXUoP8Z
csSeyH1Rv5qMvM0pc35s7+/oYKeyl38MY5xNeyikFGHJ8sc57viOihxIeMORWjTHtjFkXZoQy8cX
3oGuTVIbQNmEPhBjCxKqc7wN/NJDAoYMI8ZzfeBGjkNP95jL77f1feTBkambFFAND9DjA+PKKQtX
ejDcrUG34EFSi2YlNA6CXKhpM8H2CCaWqRQrYt8i1diQeO6e1sKELDj2sj/sH1unWc0et/Fyrp21
RCON57i4Klr+fdBs6iIMOWsEW4ZidPHM2sJw8rtqdF80Bf6qKBYUpdemY/8Iv1qRlXjt6pckKtpE
meVvZqVZPm7UbMKCb/eZmny1Ws+89OQb0B23aK8Ew828+KjwgTlh9FOvupSe7cjeIJRypaRuc4LP
jnuGPgvPE/z2DI3kJsS3ZxnhobyE5AdEsHlbgBkLJJaNT9JqhEAxDeZdZSg2wLJ4QRUU5e+jAz+n
KHECDcdXQonW8Gw1I6go3k/kXOt0090VF6TsrFyGDlDP25nIHI5OSZN8InTUly9N7rffi1ukkNTw
MeCiPEz1/rXBvanlh2p6D51tI3xs6qlzVCTWG4BnsXUHXvMrt5U+i3Onyw+ntMTyZ4aEn1hLnKQX
XEkZfV8wC/Chw9a9eNQnoxM64+ejO7nLcI7zT0umJMxpLc3jnJY2YYC5L+NaLX0EOCRdEIeZYVK/
D0XPOzqUegSVBWwPQpQF0whiVasEvs3dolO7m3NB13qvKp5NfpSnOA7BRAP3lnaw/6Piiak9iVy1
3nKuo570Kqr4GZuFWiqBzHP9dnv/DIUC7QWUMzWhTtl4EvypMmKkO0A5rBT5dRUbstnVopGb4YUP
Db9ByASLQi/KyDU49+UvczH1DETc/MSr3qTnn5r8QfRiUVT9dhH998S9V5KH7U89Z9xOtwHLmuf6
HbK6/28VtOHVBrW2uJZKnw1JGWPQE8FLk/4KtbYsu5KnHR5e2XgOHWPm0C5dVwe8AvEPl4M2qlnA
AFBfxKI2nBt2LWVSh5IhuSpyyWRDOSmli2PO+547sFt5ZJzzhqOHLst2sIHghlZbDg0bAaBPaCbT
HFwvrUuNSb41so7A2OWDDt3hah49EZCu55u1tYTt7VXrosHLEOoQlFTbSTGDzGMxo/RnEK87/+AS
bF2K/4r7Lmg7wB3dteDJP1E2TUdJsEABGwJ2xDDxyPJrc/gnfpMmuUHa16F816H1c4q41cfEdrhQ
KTsjEy09PRxy9mL59rP1lMnXwXHVyQN03Gm9XVtVeSEMHFGL5WkQf7DwKpLmebVYFMq46mEZwAgC
ea7fBeJJVFlSGsoMx9+s1jVTUiDkVh9SMFmlulas37rx15GFhohXVjBdajmeBLfqcXddoxl17Tts
Zc9yUbHDSiKjFt8OD29kcq0VZJOAbYCyQuCruyVVap9sq/NRlaN7uJFJPD+LYuih8IuLkziUpbdi
QQe5+Prl7+a8SecaMpNr4brWkcNcutHX/c2hgTaSoxy+cvOb1ovZbnjp+4x+iIbGTrRqO0+o13E3
ybiTa3IzY024orKwScwdzwFtmFQRRdjQW0ckm9446VC9mIupAk7pX+DDyHakm3nCRNEr2iPAQ0fl
a409jakivLCrEJmXBpf8C9dFVM+6yj7Fc3fqdpeqJWiIGIy9UYsB/v7e5MS6l9/mMYEq9GgzbDI2
JmqI/oYG/20Ye57qUCI//PA0ostSzkVmjwKyyr4OfI7DuGsXa3nkdFn3midfbUV2VX4gElCjB0sc
gNqOm/qMWS6DDFcxj2QdZ3fcmPmy5urt00uzqKITgp76WVrNejH+gsReyjR0/W0/Tm7CobjkoWhV
lKQok9UVNYjGsyj4tmJt3mphBYiiDwOXOW3isI+UUTVu/nmSwUJId4aSZqRsLbI7Wl5m1flDxC5Q
kwBGlmB1qrRFl2Q5cN2RWY+6TPfp0buqDthEN5E2rKC3Wv4HGEV6ueKp+pwdgpvfTT/9O1qg2e4+
mkl40Cl784aMoy+F7OKwr5py7a9+in8Y6rNBf8PUja6NwYFJXCrC92ka3FMse4T7JIqY2lg2d936
4GdnS6d3IaUX+ejftSo5degg1XNbEjO2CO9ASp/LjKLvrGVvDZVajofqhMzuqHMOf/HFoHgYpzAk
+xX0P01vIS9yrgP6Ogcu+LTBmK7UrMh3uyWDR61vVRClleb7awvFMFHH1iTX+srPbF76ZDuxVhX3
eV6W26CjuFiPsnnNVOPZhrqef4dZfCebC+TAOdtU31jpiJgAa+0y5DMOgOMxRYxicCINK8E7v8J7
qR5l4raH+VL8JCyB0jIcnr/1VWcmyV7oueIh2Uj7UBXZwpsHTUqtAucRhix23EdQbqB8E0Y8f6xq
wVbpItWJZYl1z/oEKDGzok/P7HaE2xd5LaX2B2UPeFbs4d7kSwYYyI4tSfh2hFcmlHR8/bmLGj/7
HPE4NjP3jj0w9ntzbnTTqpp5G3EAZSFQ8042Qx/fzs2Y5McrA6RugvCxYoX95DprcqkpklzH9ETJ
VudtjJZno8V+mZlnNfKClQ8mOrPumPw43r7PUkdIqONj/EZOlfK2nBtjBnymj2Ibd9nGrirafl8U
ZhGENJRQiQ6LO6iXd/PztgM5zbzBlZsSCKuDZPU+px0f3NUENbshTTOJ19rNSkxIuTGKY126bTj3
zOdYra5ONiIYZDn6h7ZtiHtGkEPNPiooAM0Am5oXGQvDX7WykIW0tYAmq+bmO2uX20fWiqQL5EaR
IHKP3mz6yoDOgWB+28rbdW8STZ3JEWclWhluxbIVPcn5je0iwvGy82oep+xQsGopmzaYxzjNsfW5
vqMD+Z90Go9gUOGiWcSxnoqLUJq8Gb7a9hTNDdvOqW2MIHXCQGOnTdxoehFpjkF6JsyA1R5IlLHb
hQC2JrcxO+rkKUq4EG2AKmpiy48N9I22AmYy2ZoSw+cnzSgwixyGSUOGNXToSd2JvYM/wDnNhM/L
NCxYahy+i0Ds82BliCO4vPn/6AjRzLKk2HOsqkpij0xDOvz1asqFRYxOeIaL9uEhrTskbKt2Klq7
N0HSDe7Vme46pMEXS++lWxlpOZ2Ew1gCBU59T5N16y/gU43DS3Nt07z/K+SPJ0RIMiKQaTxTzmw9
DbCU3111DyfU9HWnbqOIf4n39IzRC+ud4FKh+FGKqYxH08Q1ZuYyOfS/s/aqSgo32YhK1ryW2OSZ
3LHXo9czrAS1wQFdf9jh+R+zM/NMJJurgy7G1U3gnRDPT32xDbsxU2NZiuhQthcwT/qSa1AJaLKI
TAixn+KmLa0Wk6Vw/oVuzBry7FiYBdKh6M2B1sinOBbi+5c96jOfctrL4JqO8s4h3ADMgwQoyWvP
XHIShYfymR+TB6qmgKpAP4BZiS8Ix/xTnd5niKciw6wXbtKmns20iK435f9/6y1s6JjZ3sOuK9KD
inmiwHz9nROAgGtWsRQGQaVyw9te22USjPJAI//q/G25NRXps7ljBRwe6QQYgMn1M1/RXUIALc2T
7JzC4XYdjbx59otw9x7eVBSWGdj1lmAopCPeOEU7nl+FJVOpP74y9GEqUG35oKCIR1FjM6KTrHq0
VJ/xIkfU9NTag+r8cw9yz6KEFrpwpIP6iT2uqOWXtSrAHHhaNcYzI1CZI30yYwU9ik8JvI7bm/Ev
Apo0ZAdnC4vRYSCfYFOyuYjOQnzqa65Gfn0+jWq+JhEdJBKWk+iD+KK7VToaZlo17kFn/tKOXY/L
GwzyIYy12Rn0YkLFz/z5/ciS474jSP4+ndbNrMq+g6DYOwyuYqMhs0klNvUmgeNFUVC4xDSJlcO5
YUHWYQzg4cjsLcPXwxBGPn4YndGreYDwFPWTzcpauz6d6t42lcjnuHZH/1tGyrAmYwvWOjK2qxa0
9W2iwXRLQB4M/QCN9czhLuJepp7c9s6nmyOHYCwwxmurx7fBm5OjpM/ycME0Znrfa/91hdnxzr+5
zjI6GlmtsXIFNOf7T6YSGpi/1GSWst91UqP5pNMqMX45Xa3wY6YhPnSSiG0njokPlKtoUVDrDvA7
nO9pJq4UVZufc52UZWNB9ko/c0kVu7WEvjEWznRZ6j4EGWa7mIVuUIqP9xm5huIftOpEh1TLQaSh
+SVNUbtAZF0Hmu/FS/4/LLH1kwOrAcfieR3P9vspF1poQpSiMTBPWx0Rpg1wJeyBrjhCcQ+xz1It
Iyx4GSlBOlkxYDFzRRYxnVuUfXz9MnHg+0R/0HLRKNquM0mDU9N0g3RLdiN4PiR/A5BSTKONKSBQ
SEFn7nSlxKtGpj2k2/ysELoIts2THLhjMYbYKu4D0yB1k+nLkAgtI9Nt9DUTn9+bXSt+ywMElZb2
jaDr4g2VHa9LVZviFGgIbiAFRkOhtSSiTndejzhvtbTgyZxhwti7WLS8JpsRVKvzq/5P3jXYcfgF
9P2T6i+qQoCSME57H7GLj/+Wzmn/YS71r5KGbzMut5NRNI7MGYHkDwDTtJ/hlNNYjnjBDaumOtiN
1doqX6uNczKZ4lUvYqTaLt9IOV6I3b0sBlLxR2ZNN7BOxLs5L62Vcb9pCei0S8UfOVZWxDwOmb1D
TGP6HkiHq+nZMhMKBXuxofuIjiFcGSlv71zYi/dK28JrgPnjbOmB9iRLSkIH20KE2vaSBSSe1uty
28K7KdnFu7qkXkhgCK68MZ/mYmVmB6F5iRbQtdA6ZHVKoTebrAiY3fbr9hcnjTYGt8uGEfFoeHK6
39lEtHgTWgG1SaZZOoME+BVhiwBRVTI8c51Js832soVJJgSSlE4aE1AS8xKBu4xhOMiX+gJovwX4
3alDT7FG0mDgYEomLrODxBMj1m7wpwO9IdTEzy7mnuQCpWr+Le5RZZF3z22Q39XiKxt9PZVGPl4y
z2Hn+MluLfolw+Ot2hAEHJjlNJ8Y7lvy+nsmIek7fLQJe6lRxZfbhFYOMQ/GVuKSQ7Z8KPuletOw
JUY5/gLxhAZ4IYqQYnTgBQ4GjDD8JEkir8I/UVoSrwJ4Ina1oAh4GTqu77z+G4op+rnOijdI8doX
tXaa5jGYIrtp4tMNj/gX8H+RLtePP9i8RxZIwgSEbOY5yJ3HEOrx7hF1ndTxRUJXdjVdI21Nsazg
3UnMzOTjbaOSC6+RjWxxld8tPOBEYCOePvZ2A2Sqawv6ukh3lP2clVZCzn8DTc3828R3PuiabPp/
d6UoG27cnq6+zf3CNVFPrSVN0fJYr8/KDWtUQd+JDNwYWhuw+CxeNjSCqMXQunnCt7sYIMdQAGko
3DwM1axQ6UFJ2gC6ozGPDQeVlmzqgQn3uwA09rxXxf48ilXwn6w54kAgcAP4Qaj0NnFPCj0JKrZP
g56t8GLzU2TKPxsLY4C94kbp2NR2KO8yLuPo0oWfOs6bOXlJqAOPue1Qrqyx5TjhbvIGKS1SEot/
JegCv2sEy4Hx+Y4ZfQOnDNFHoh+rPn2C+X+fTSiJeiXJUBSIRP55j8+t+xwBkekbihp1hpaMcNpN
0N3pZ/vRTvs/VzXlSGZa2emgps8EsW1eiL/0KbYD2G3TpnW04pYoCgu99I8n46ONYE4yrD3O9goN
3s4SUyDchS1ebaBKdS8f2+19Bq5SsNBX3ngvPJ4XKKVWJZpW2pyHpUWI6NeSlWXOME/jNzAjrOrj
m8UUenZZYOeGUWdylFnbHioieh09K2YnxjyOJGDJSEtfJhWlmtT6kuwVI9zffAqs/whde2FtnH1q
GYGMEKa7ucXxfZwdK62eAGivYw4nesOm4nL2O63RIqd3Tih8l9VRMSqEwBfPv/oLftC39niWWrva
S5QeVpYouc1BhdwKsjDpfqloReGq9lLfBt8qjgggysMULBncHIhR5M9MsMvJRVn7TbBPWoIAq0lc
rBkcSJ8L5bw3FdBacXpNtOku4TMQvrb4tOKcuWPe7whUTT4ahO0rpTrmeI/rbYmpOkVZ/BXIaSLv
sE9wKX9Z0PvSi4pJ5K1US3O85shZYQyG5IqXq/4RekM8dCvvfJglO1RUdET2l1nxFjUtpFdd1Zbm
hKpv1/1FHV8DOSVNzT+v4oPFz7stn8CSHEm4eT2wrrTiLuI5UU1sB0k2rZqmGrceN1XPlK9vruE9
HqjMRIr2DlqD4AL6ZAyo9cNmYcwRjuBQ3dZJkv9T4rdQmwi2PkdPbR8aFt9Vza7+G57nx9bWKmFB
C48TVRMxmk4fsSlbol7BrH0xU7FV7VQrTiyxfA0A3fqI23QXqvQJkCzXWl1zsr73lvjWL8+L6wXW
6aaqjKTkUipTDb9I1OUbJR4jnfdfe+qeBaD6R58+VrVKhZIGEe0Tv0SibEgyYeHlVVvU9Vdhn3p4
ytrV89pM5BgbWlinlkk72DwkaAs++OHZ4nVBhiRdk6DXylBShdcxPUv9NhtdtZFnMIRm6XJ7rh6e
z6H6CSU5pXhGCWK0CAXMISHjXgeXgMDuW5UewYgEg6WGJLfnx44zE3xui2yjEV7dJmD2R/W6S3OD
OvHzCplEbr8he0Biijcf1nf0+e60xfBBf+FLBzNAvFs5NQqjGxzLsxcSpTxtajY/rDIgUWvUO1B2
+KUTh0brnnRsFdDOXlP9uZydD7SbB2r+7oxJC4pf6K4dpuFt6wQh82KO79inTojFsEK28Kao4wHa
1dnOb2xCQ7/mhJxelW8v1S2IcA+mgbdGVztO/kHY3WfukSkFb7Lns/B9kdpcUQFgIKEZ88/48x5Y
usSQ4kqi/77W0NJimjXCl2+E7fQ2v1jFN8FWWoO+dGD2VPR4FwtdF44L8PHH99ARvsPxdCEZS7X+
Q0wqJUfXFCkxCAnhEOfCUJl841nbC9C+qEkZllsdWAD9ieBqTZrTNxSLTaiS/GxyGAwbxk5clL33
WXLXiJeCmXhXeguprlAPskV+DU/LGm5apfxx5I+FTEF/rxZIKrzxoPCHoNz4A2KLxxUT37tq6Him
0LYmj4VkbK1O2FmfMKH8DdIa6IoyG87+bDVBjFP2r42mw7+AHGNJV8s2cghvJewR3RMHZ6FCmUfY
jIpB5nsqnvXlcNOgdbbsNl11VXZJpwpzn808/4gtgK3JmpSs0+uO/maT0hfFYYoBshUUYoWLb5T6
2yDCMs9NKijbbq8w9c0khbg/UIZ11VIApzLM5usdGTw7x0+vlNL2zXRP8sztQyfsUcwUZ9nkyRHw
6vfnFO7wzkUdiJjDEx4rvh+0mldkWwK5CUwRiNOz4u1iujJpCHwW808/aXZXlZ2vXCLofpSnBLPL
65SHJhrfZN8AkzMYFsESkLzjVCRj5VErpr1qRT+FquZM+Nf1XxWFqZDGtDAETOaBTlPzbkfS6sDs
4QXIDr1MPcFDSd37lly9xhl2BJjICPVWu7tLLEjRMIUIx6O2m4HrZ+rugf0hwe1kR/ju457dMUbW
Uk7797EZILvMy+TlCTFr0cEpa6NR3inz8yTRWigpWVLfZbeZS9GujofcyBeD0NnwWnoyxjpgS0GN
tgZS2pTl06M805Me5nP2O3vSuxAVoT1otvlL7dGp7uQr0+T0WMgHkAPf+sCGcjvOVmaUHTaGSjLi
y06RXoF70o/VEAtl711LRCfmcSS3BlnnTBAgW4Sb+9BuGijOUEI8yVpzcaO0TYj4Ymuxu0ujDKLK
fa4lFjs+0Z8g9gETySihB+ot98WaZ/IwRSDHPVVYuIn/muuTTyEa6xzvyfxUaMpocgOTg/8lh1DA
cNYnbpmCCA4qgmMRl/3f/cDSev4MjPJzMiSBjwO+2weVvki1ILwrAumTLGdOeHG3qeRlBsmNQH2c
zDKVP/6WEU9upeovfgkPi31mj+sNdL04ISD8lTFXw0FJgJ7CyphVyxfG+E5ClWhm81H+L65ZhgLN
FJd6dh0yKFfbCXbNJ7/LxZOuRedgjsPRo1kWq7fK3jtuBf4pcrb5lELwt8L8/wsQMvbLZ5ox7Gjr
ZgHSsOd3ythP0q7+3cvJatkEqNTXwiaNjeJSXUwQK5MuL/9XzJE2JTATBmnbT4Eh/ZqavA2JvbUU
MSdtXcntHO4hGyuAAF4hPcjXsEk/NsIgSIXOv1PPMjwV58nXxg+LpHhnJF2A+Y39A5ACcBFUfGyW
Pz7PzN0E0PqBFGw2cND5JOGgzyHVZxVeBaQigB3scJ7kWRrd3rKxkGs2M2MnXJbKC9DKiG+qdBGU
HGOnVBsWlDAZGXvRMmEhXDriGPZm0/XkgL4cxh+VU9irBNX9fqdOD2DhY16RlO+/Elz9VjNQ2Uu7
qw51eJuf5x+QXSRGkqdNsjeRvtHh3qhGjgUBTXiguncPIdpmh0KIWWSO1y/SMD0hsv9jWztG2EjZ
tP4AHTEgMZbgKZtuHvaTec2qPK9+JYruIUjgtdC7xiI4jD+shQb00lgpRRKRTgxtMxvw1hJoIzjM
cauN4JtDr38hLT8tmW+05afmYs9EvfjpyLX4d/i6SCNSWwh7UPpfQr03OLOicspsF3OWq0ktTVX/
v2pMcNxvcwgd3D/ZyXZCO0WKzL8zQ7qFGSIHQyNYZ/3VAnC+MzsvwNZy8Vz/A2CmT57Lc1J8t6j4
/fFblopgKRHdWaIZRosoIlrVlV1N5M9DhiLxL6otla+Gc2GZXyskYKjSbI/3Granqxnq4VxrPW+c
DUdAkrOnzRrHTGOr/lIfQ8pouOd2rDBtXcXnjA41Cmzc95YUR9D1o70FD5RZ4giiBN7IjbbkbVrN
f7WcP8cdl9xrpkyt8zSZTnsVCq9oiNL46Bn016QfZFP2jTefu8piztNA9+GGKv0GMMY3zTbA+r8T
Cnwb+P2pgdYE7ca9In553404vRhf5WCnXSA4K5fNMKbIWpZCB+meNu7CWub71+Rm0z7NyuMLT4Wx
VxQllKw8iVpA4hVFaJ1KUxFz7vV9retmD8hFiDJK6Fnpi8JdFCzcfiksxXxkVB1Np/DDqXVUbfBF
/j0wx/udux1XieomwEfb9iyrh3AbU2mg9zInwThsPNWo2gIoOvleA3eJFledXIy+/DBIA9ikAvsQ
5qK1PMRA/m10d3I85uSenINUiwiyyCbFlSqLSqHTUhgcxIcOMLLrxWcu46wBkhS++QDW7kn6J3do
l9jcpLItlGwv7pWMMIIKAfhn7cqZJ/JMyi9gVjk4GUQoP5VUt4cEluDbHtjikRtneuOxWlALu480
S8+TEGBZadS53xjboPncZbDe7jFNF1pzJV/Z/eerAM3+qMwu0ahGQ2NS+JJRfmxz90vxSAkMGDpF
pqiYnkZZ//VqB+C+8MLPh20SMcY+gy0f+ihb5tq8IAMzDnJMuvkmKrujOkFrN3ph/kx8CA0xZfRZ
s11kNFP7RPpQCZlTRK4q1W7IKTHUljgcrKQpuRUtbYsbElRMU07UibjmBUDX9aTU07qwirVj0+4n
hl1CKXwD+Pb4nJ3CPSAJIMKVdXnIQKe/DRaBezugVc6iaHyZqzHFDnZQ2F/7FBT53Ug8uAXGZisG
l6+5Vx9cFSocRTovagJbXidhrRQywgz8N6ZDjPuLhWsXxEgTYal9DvP1NTGR9swDqY37MkRJM8u7
oq9a7BGGfKWeqj1+3tadomWjh+3eJyuE+93wcsIn/otXjzqXfyMpdoKOiPW3x2wXXboD22i4LvtW
4MYwbAPATTVpeFNGIIQctlr8hPTIlVl8FzgTi0qgl8JRfK4p6icTksOYOd5SDhadlNaw+UOeUYr7
s9+C9lx7Xrii3Ig/q8YXWz0wyTssJtDeIrAvGyv2Q4A+bet0+GGd9SWSBDmWpBAc515OuSZOZ1fX
P1oFkoxsn3IYbZwxc7AW2xdzSGFd5l7GDu4rTUG8XGTtkOXUurJ4jPuiydLqmpDIjSp0gaJ5i/lC
TSbUkOEz+nOmakpiVuCUvIjitZhBy6FQRwZDP4RFF6XTEcmuix+jfgPRI5xTMIEULbMB8CT54RTC
xgR1Ualbbp9+Ybxy9qtJanRB1vr/U3UBmW5t5EonqbwI2AP5+uAq1CPklbI5yBeQRKJeAq5ZM4cK
MJUFSPeLK4GGTadyquEdN7sYLzDMY4JeMr4UL27orWy2R3LQCKqj6IOR6txUw8MvjUqUSENOZKIv
7vXsRJMm8ncuV+1uahxO693QSO2FLIZFOiX4zAtN0hkf3ggMoAbenK8V40A403gTo7jLmXmkzQ3O
3SfVEWyxgBvOokP8QF98zVmbQZn8hAyGe4wh/HiL5QG2YadAfIHQrI8ej/Wy12M9rAViRYgCxf4t
+EftaaqKIfp5ZCcRTcTiym4yNoE8bISyDrUFmkyE12X2NuhO1qNvgLzEXYHc9xMzi/JCWf4waV1C
KrhEFnqInplK67L4zEgefnywDjPTNGxDYZpPEvwkj1LFMMgzNkdKiv9F7DHlSguVZH6R7XEuwLao
f9ggB2zTlO52vraDGUYDhfolApZcjMR4vwxDY/DICu19V+lc0ud71cX7X6eR7au1tcv6zhI4fnmi
UjWMkA2+OWeK9zMHM6CLkEUlhjq5GlevKU4/csSqV/FJZK73JWH5uA/vJL5aPJ80Y9UiBZCv/EuT
O3PWEdk1u9qAEiD1mouGZOg8QXBDkW/vKuMMF4RQqTlIwq9ol9PMZTZspjwV7u2UY1QoMBnw0E7A
UlcUvCigBCwLe7WRbmoYTBfs8biprvArD7eIyJ5mWkiEw3LuZYlVQT9uxyZU3Y2bSF8hqjkVT34f
bq4m1nBwp1nv14VLP+CnZWetZ0SXVfIMP9kvjqDY9ksVt2rxQZPtR5T4GY4QUkrPiITQOWS3wQCN
y9fBcji9hhCCYh0a6sY//wBxu/YJtHpuPzzowqo+SG8b36FnZ9R6O0igSkABdZjZv8mn83Ips0Wy
RWkb7lfRkWmpGUsj68dG9sfz72Iqxb2nQzt3JafsbCgRNs4gUZtnOjNjzIFY2uRtTRo5VbNaRWNT
qityh8mO13DS+us1tQFfCkhsXOanhsCQEi/5Kcss0p8GZsSPLxljOUtEj8mz56YD6Jwf89A1pGmY
hNsckPM3rlNmpYrMHKLNfBtcEmIqEDrWY7b72Jv80SELjEc+uuSB8XrLMn5wbUgpADxcoizf200B
nWwpYtfRXxr1sEGok+pmpoYiLPy2E/e39pXdymPh8oderbJzL3RDMppMBbv7uk9emtcQE2lzn8Fv
8NHdQLWIOaNi4OoYIYYPKqw91Bo7MpGw1+c+CtzunLrm6EMdfuh4uYWKNWirUkQz3eXXChHonP0d
T5wq4qz3pBPxjNGBPEbBsPH2pV0AX2myOEkhjaIRW6mgtQ3XobZEeqPbrKq2e+ANCSILU36Usqiu
1wFVUxp92xuoQyHOlkmCBXnvSXFr+3KN8jsvLS5IcXKVBERftd8fP5RMqc3nAb7+5WQRAQLyoFgr
rQiu9p/WS2xImEvi5Uo9XBjm8PbJX/AJJgVuu5RC5410XmTiODho8M/nxEGuXD5cg8Am7aMDH1Fv
UsuW9TPubm6NTDVjA1TeYHNawCcIpK8xH2tC3eD+m92CxdbESTS7qDFNvVRwS74R0JQ9MOyQXbkH
k6LulMmxJpys0w7G4SoV+AUxUG/Y6e7x3940PcWMqqEu4WB564aoqy1kCPeiBOHwZpJWraonp1rl
Swg8t850/+/iC05gCfLOPIl4ZSDztxeaxMv+VGK5ly+HGrXM5Kuls6OJWNZWK2vOgPje1wUuXiFL
dDAOcEF+x50OWmMsdBYiZjwjYbw3FVY5Zdty3cU3dtuG4eCi/19LhoO4SJUyXKT94vDCBps1gWP5
XLFp2xQFDcPTk6DBYvJvuGXmwUfahz5MkzvX9SDXHrcHixoPWMiw9gjPsEbpXNfutPMUg5VP1B2B
KLAJU20FlpW1buo5q9iouDIxaKWFXqkZuiZQEiy75h0Y9A11QPdO3+O4NDmf5IwbIDohhTX98xkH
OzqDj3wOrDZQoY1miLvxzJ7a3XV8d4DHpuFJJWhluNbyF+E0cb1qt7r7gygYN/1KFo+wEZsdaw30
QOredrzI6OlZ2mn6HipGWX59wvvPcG9/LDXRChvdPran6oLCrA0LEltWSqkZUgaDl3SAvrcRLJF1
6D2s6C9RVVW793NnBIjImyr4I/AUQMCFd9KGrx+NVO/2+w6rxXvHerRe6yh3RUk7AvHjITBvCIWI
k9f1bVaCeKCMOrsyqpRWzJSTqZ1u2NDit+EPdqxuvEJIOCIkKOHjDUVlxh9z7PUdWkO3C45uLi/C
kcNj2E73t2EDm885p+R38drY5XgPZXWNgH+HiGxslAby2t6l5vDY8Pk3oO2aWi967X5JiEFHNI8U
3HME56Aw5388A3RBXmW85HEUM3VP9Vv0vSPhXViCAzIqlMwIGTrrPKKd9xpfRqw4LUTe9HZmC1+l
x8+M5qwksBEaAq8AepYxTtKSYqYuU1f52qo3OnWD8hxNmtMVwbn7azf9b2UQI66hQW6y40gSBPXJ
Q9cXElHGCh67gbUTYvpZtn1Tt7+PYp659EP79hp+sbPwVM6PTKyBlsxk10ZPm6Xehgitc5LH33H0
/rwRsnrymI1XypoFcfrHy2pQvclyFcqZ0ZrIFaT6ngUo4sxM7hEDEGNGCW4FtKTqGQoDAJ3s8dEU
IiKV10eHJeeaHAUMumyg3ywbugZMDA0Eo/quwu32noFZS/QAy6zDNcPncch6k37T96FnPbeHhkrt
Fjxw2j+yP8A6SVH5yONBQcelUrVVN6bssv+LHuKXY0HuKyjy7x7eVAn9ZYml6FMrU5rSXmm9+Cem
ddNFeOdT5jMYfVmqirn5YQ9zE4FGvSGEEsvx+etOoibJgV/SPPnLw3WEg7aHR0JcbYZ68gyQ0HRo
f7qbUuRYyIvzjGk0vD1VuzxKumXIOOD4pm1J/GGQlMtca8FpwY9cLMw3JNgOtwpZKWAWgf1vaRm2
0DD0s7ON2pxoYk6B7l0rszq3o4D1tHDlGSEcNg3fzylnPX/0pCGgy0ck/DsumPiIxv10JSdceZfp
pDw9BCB3OAeUKW4LyIV3t6da+wdlaroH04D+aBNxU3B+0L9Z9TrRNKCFg/zYveMoewWR7/I9vLLY
W+A0EdIl2Ftzy3E/rl3SARYq9g3PXPTCQmHlnlTHVBU4JmOUyjTJA2UMbjOdUvnxBHCJkN638w9k
meOCN7ZcoyBZ6R7j/iLYVbDKsBIdeGmVdQoSM3nuEJCq/1lMppR9AgGu6tIGm/Ni1TR4ENWAkGYP
RBAPaP6yzLIP3/pAXD3eWNhXphreZZ8kq2orpjfLeScDpkuB9iDdOktCT42LhWVU9NIKvqhvz+W2
tFpUIoms5mEesXQmeRId5m4DBjEXf2jm/4Hlqp3zdo0wXLYmf7oFXCHAuJ51NmSXvHlq9BOiYMWS
/aHM23uXssjniz4JmZB77J+xkxJhIKNLGxC6Mbn8StQYAEwebYXodl8k07t2GmqcRnGZxzqoH0d9
Gd8+4W5tIEI41aqU3G9ulhOKYB0OLEkmhJhhjPgIwEDazXg9SGKn9ApZ+8CXq9SLKAdEMOtFUy5I
B63lEqBJZwGEFcgBggi7uOVCxaZ67u15i6iOMqsllC+KZjQU0rmUsnfcSk91Ol0hf+Uk4iP4e3aD
r2aub1CYspXT3jtTWnDtR6hJMJz2YAhqo3Bg5Rw0KsLEGYbYwHRhMlKol0B72/jvww5GQNpYvaDS
99nD/R0prkvIKs9D5FESbSU/uAGTgJBDXxp5OSNAEZmT9rlXBP515VCY7wj07tpOGRPw5v6OwQ3t
EzUO/LzKtHk7f3BEoUZpNv9LnCRzoabRsHIhBxljJBSTJkICnCR6W8D0GBkX08grA0QxCT9B79mO
11p7ukMJEOHas/OCb8kIjAudFY6Umxjo263OMUIcfVRmAPYv6m4PXoGzWx+pCQgEfayYFLJNQoEX
B7a3muvc2U1yN1iawlozSKGDG3r4mMGkHeBKgFL+ILRPFniGy5Jz1j14YbTkq6R1UchJkEHWzD9/
BYBC3eH0Ao4GUum59ykW6zWRTJHdJBhqpZBrkbuNs2mfaN7jrUeIVtj1IIXcStLlKPQaBBTgGw54
VzPGMmpJFC0wCo2QiAntP9ihDLDHseSnsrYVQjenvIB6k6HHN2qvu3SKHwI5NO46BCG1Wc/4JqHw
HtrrPWRe7eNhlduhY3vbM30Fd51NvGicdrvhCUgt3/3cT8dtRbFz677xVL7eoDIrilDVg1Qjc38o
oW2TneztGUJ826WyhYrqgWv8iJT7/TQKqXCVMdHEcvN9ldAWPT9n7JoCm4QhXdcx7S//vjkUJaA6
+2KxTZeMYpqfW7uGpaVjVyR/8TOC+Dg+XB8Wao+B4zQqcedl2Q+8CM42RCmKuny30e52pB6WCDx7
6LExpegSz6A5wbJxxV/T7pRPcyYfEz5YDdYlYi9xHemfkB6fB+MT6et+UQq1Kiv9YLyOUZOvBLQ1
RIuGFxcjYE2kRRIni5sUi0bE0TaBYDMCN4fdpungiiQwFoPR8xyKC7hepuH1FCznA1v/0HPzN30y
mzxKc1ORx0FJ5szJnNOorkWjc2hT5bb3ZTr6DtGYorzdj4H9KxiyybTWRBtFnasuk2zaQ4D+sFh3
mSwIDVVuVLbul4xkxu+ZTRmqB0YfljuFukp4R4RZD+1Mhaxu/ogKDc2+krckmMJeLlHj/dtFtEc6
IX6OY6F3Vq4zxpAp9bQ0lMx7jn0sgNdIHQqotDzlsqcihmFIhUKajNA4m4AsCEusl+biy+OnO1xx
Z4BPvdeOxHTOCy6/1+ZcfSAugevi8H1dmA7RftrYgijgPJoea6QMjJRon/mdiS2l/ySVuvCzPEki
C8miqS8C3yRbUS+PCabE2vrBbzDmCpYOGEpYXXVQihBAd0w8ti1eJ+JYdTiVSbqDVxKSFHQUzzaP
hJmK77mqTUKGrN3YCLnx3A421qA61PUyoTSm2HVUqPtVzF5R1djPGpTnGJNpuYVpOTBF1hv5U2hl
qIKyKmYl+VrNxPZsaq4He5J6ZZjNDHG6RbryHuv+McVXgxd4XlLzbvOmekvOb/K6ImZ0PsE+15HX
3U3DHvHWdwNNlvwnxhQ6W/BIkHzpuiL6Qb0vo+xUCLnW+XGI6Y0dFOIxtNnUZVtcutnhRGuQ+pYy
1QuU/7XEdI4N2eP+ERUPkIeD8un+XIcebW7xEY5gH6SlVwVnSVM8gN/FUZTut75VNOlr7xfwK3bQ
6qFGJssyuo1v4o5g0PAnittAwZ5xswqYaRMFHvrm/d5jpAhbGmglmWX2DzCaOWubod089W6oVR/X
iodUfHCPUFhZpyBa9U/gaq2dsJZeqkGtYlhbFFqPBEkM7YOgMlvM7km/1R/uNwI1J0LaSeypJFC5
cQv+GW+WmWv3pwOggVSNCNEOM3xQuC9WQhFWxsIsFQ7L0zIFhV/HFKLTmT6ckG5mRxPHPPeeefUB
20RHnakmHes8cnIXasEBepKSSE92EQnX0AYvwC1b8cakbK1qPhHSLflDdhXXEFUe1bTkgQnrGjWQ
kVMjBccGxbsEhsfZf3jKLZpqWST9CxVbL6LC4p6tqZakhFguMpa1GO1O3DyzudQLlkoBlFfRXB0m
l7MKGVRKw6q2L1Omwi3HbyAoitahBVLqzUsQikYOB1JENOtz1wxlP4FiU5m9+v9poCrtJFFjGoLY
bVakDVUNKvddLa8GnQEswIaqFXwjq2kNAUEHD3NEONXowzF59fM6JOXzRenjWbk59b8ypi3FmZ55
faHeWUAQfy2HCD2axoDcwYB28R3/GalforVwbvx0quf/OerEiumKRM8Zgk6JSBL2xjTQdSjuZyvP
F6rDnWI1jtRyWA+INlOjTbOHwatWYNuIvzJ8SZ/+uJTB8MuY4lobj6G3uElIzFrx8ost4CA349YD
LP/vxDmXJ7n8IuBO48auJ4JjM097D4dtFK1C++mk90fAXuKHxQMBRacuh+3FVS2BKoD5W2btsUcR
2qho05Wb075ya670ALbZ9TfUBjdfChzOQQsNYiDyiiOeg+gOjSEXuUUFusWY2VpdNjGCN+4T05JS
uL16TEvZG7sIgOQkfGfbuHLLDNNpjY+uvpW1F/olwDIpO2L4irU/c6FoB8IRGy/WMWgtVqfU8kXl
stMOsAFvaN7sA2sARN+qDNBWnbfEPJfosRRKuwUl0GCYqr5rAXfVC5xdLOq5tGhsQLKu9nP76D/p
fJmqmOmyI34crt0TbaOJyJC22RwhfAxQQJc48GMr7OLfxZsi1WEzw7DBMIEIXEZxXlW9XNPgqKIk
gljGGiKZ35vseGxS1xw4Ode3FvAOWPK/q7mSlVwCtDTVVfofLOBx2fN+vjVXl1UzRtx2K3j+1D4o
BmPishdDoh1iQbs9UAatcPlfrJ4B8Q2g7i/bvtRoz9jpEkKG1lzglG+mBYdbHNJTwzU+y6bC305s
BwO25pSWmItJmCIokaLvSosgJag2/+6z16oKx+aLTJp2iJ3K20d5vj9y2Qmo+Kw/VvlGSWr+BCIa
N1Rl/Di2s+Vtdt7+yAbsbncjN9DpFqA/cuucHH42CWHc1QU5tH6OsdArS0Oa5r4f11O4zZQL9vTD
TpAHWeTULfJcZlc8PkitXrhSBqBO0nQf/ugTJBGSlN3LR1oFb8ht4aXMnn26i2Jm/mcWa05zpLm/
l5po2KwdASyhQ43nDqxKcnHP/ZAz/9XzBADUiHqs22tkkK6OimQs2mhdZk1no1DwI2rcndPKRTa5
YKZXHbE+h5iA0340SH1SOkr04gKXysP/na50B+TgB2jymRM9Sg3biZzvzenLRaq8VfMC1jPry1d9
YT3jTJO04J4yKX0FFztlEYPeZypmjTsmuQ8cnGCilAR1Js5XLdlgg0VrbLHpR6KYrZq6nGts+6zW
ja/q8/tEzqOxBz24p+xs7A3YSrhfw2JSvCsd3DCOzuhBpkyrH2a+wqo+hT+oiArKK3/s+kbqjhK5
7htsEgdUa+XsV/cWWmJIZGEHbIMHnrjQs/qVDbHVC40Ay+fRNzsuUx8MvgTyoDXGq5ge1+9BtClK
hvaVIM3nK4SrBbOAVyuMSLBF3KUiKbVpRd1DdBPlEeGay7O/xDRwfk1iIMDYrK/xAm8CNqiMKwdK
J2a2ivjiw9s3DPyBhhCTTyN1Sw9mfMU57BpNXv85bl1pnPyHFDIMA2QuOMqvynx6wGpoePts1mrR
0k1CidsXzPL+5dfDk7pYSVZKoGv+fndwoiYqqrCzmYeBLZOcm0Wu1Bkq8sul8TT5pMcfPE7uvxuE
37LwT03jGpuWbsNB6nHe6ozbpMp2EpNQSzghfh8MrC8zYD0KbsPUELkG6WENyM/Dn9mNWTTW1SXn
gDAtQ5B1M0n7gwZIvjbep6acJXOUMg7qxl20pLpsQPwqDhfhPE0cJChLcEVGOKUvGpIp/CzBO+uE
odiOjs1/+Ol8IQEVJOURVuYIRb5eQxjdIOXRiiXiSu7rzgTWMoCh6t1Gu5+pYkE1oYT8IrWifQAK
UHFe5kUYgdNOFhxDdIzNVHSYA6r8BxHYkjNx8WW5us2Sgd9YRmH4ts7elrFnsHVTcixEYpF9D+Vq
OU25mC6ngYQccXN+R7/u9t8LH5W5Ed1e7AgGLSO0e9IMyrfoD3qsRoFWD4tmD0FH39pXw9sd24QS
0qqYh/NABTDjAA4dFPBc5y9EUnsP6RYRk7PsAShbyrwWmS94M3nmArnJUxWXdNXrhedyye1GC21w
7cDh1b8OY9rJDREjxkyp8jIHvyJxFuosWxC8ESjsBnTK8ThJHZ9Tj9km3i9CiQZvmiwI5n2J/5IL
Q12zuAc8PbNebOK21wKs44DRZH9nTkIgZrFWMbMOYIql1AQ6BM0mfcBCNlsX9kxflwvs22ND6aQ9
P4Sa081oEUcdXfGUN+YqrWeNGF7ap1DrvfF1Y7RTVt0+msSGGd6i2hegQvf9DTYuT9apfiaJWthT
oCRgiJd/qTuOl6O9pD4YmCeMuTRAqVaHnzyqzJvmBvfJrAbAYa99C4G5MH51mpGnw4Oq4YCBv9Nt
YRskx4+DpfayqUvX6Vk/VkdlYzUqPDNSFGbtxDxwZihkHC/o/0+415fP7p9EkhNqpiUJ/mh/raI0
ApHUBXFHoAG2+j+pLDoTztLjNdQKE06x1TZpuRld6mp5HVKATDdkAoaZFDVKClb5PTv3dJycVrJW
8vuUzenmGFym7j/lL+tFk+0rCNAHIoorkbKShppNksi687qgNBq01UNtULI8X0DmF9/SkZMbFIpU
/bhGb+W9a1pPfzco+/DxOcxcChZIE+wMjiUlVgWJrg5SWWwTO2wpmtoFlduTgtctkNIvG2BNE3jg
e0iNAg6ipY50OVTgoB+j8Yr3oZ5GVqACmbjPf62uO+OjIXYHYMcF5v6+jsNIpf4bVwyFFgX+MAmy
ozig4BWIETCfQqrSxkBzVOmxQErQRrhz1SXn0K/9+tDdOTpNL71wGNqvFKr0d8QMzjARuLoYC4vJ
pgQ/jJMac+9sy+qWrA8nvGBunIDdaqYV59BExbMCSsU6TnM2JLnOi5zhCErLTrPK8Nk02S13PfxK
K6VXurVOvzyJflrOXdXdLnUEOd12aqqsu/sByVTFA8ofTESkKzL8lweWIxAiTJPbTna+Sjd/tGr0
jMC4IHQn/yqHD+XBQvwGjaYSXpga8RwnLflCQs/HBsGwj3CNaeD/edOmKVhEX9gcmO4T3uJ5v2jr
LvWbcfVDrOynPlHKGdkhVxmiVEnVbSCtFuP0H2Ilc/HL18PcuxqD2vsrHxlnMl5Bzvd7axQy9Dv7
aHthRFzp53elhE2uDqcV1sqhr/xmlB2iaoS6Y313GWKMEN6kINUsRfaK/N9IokVQbck2hEHYAroU
005LszrgBvCh2qZWO3GkVjLb8ax9BbDaTm3Jj0pekVLmNgaGqEJIpTzJkP+pzIeSKY8gQHhQlu/9
E9wUUviE8N7vVDZzl4ZYX3AHwY27G8qig5IKv+QT+fvhAWbTnyDWy1sDEzzeEUenVxsBZFlylDcz
9W4ku1Di6jwmGF92eFSrJb1/6PAjI2jG+4ZN/fcu01epCk4/BU5+mI4m/QleNnI8jq2ss49etaWZ
wgbZvbspglJ89tijnjFgmae1RAMO5EbcpZdp+ggYSP7SENi+EsKayTD9wsuFMc169m7CsYxFqh8p
lrEsIXgkebNCnXVdGyIQEYzj+evBNemM+Fyz0O2h5RwOF7CA3SoiIDG2z+iijoRnWz/h3yUkvq9t
YO6NUEJpcGascrQQEFtFfD9Jav5Ir5SVZDmYNzhZg1LO1YC57HHirIP5PffeojsR8KpEtBGTjzSe
BUTL+wy0gjfT4vHzLy8zdxgaC4/ScVBxpq6l3iljnIPpa2Pbm69Rf2bMkis5EVjFZhKdODNY09e8
Bg35/wOUKkTWizYG34hEIILr92sy6q7baDedPG9KfzF2Fz6bA8rKA1JOnlZTycS+DDaOUz7sa72H
PU9o2o4QNyijkzpu2UheNQhN9d2WLYXqvQGda9pSwK2ufHNNEZbnaHQkN4Ae1noZHgDyPlaGgIw6
svszCzq7aH/JDQIIWEkij8qCqB80tXAk53BRS0O/1lt1nIJUpukqP3Fb/M0N0AVrkhrn3QIshnIM
/TE7293bNnGLkiUYz/vq1pxGEibDik1qR1zX15bR2fR/n/Clt/prLz8LmKkBlO2OsZc6C4PV/DCb
II0Mz7+RXAVMgg/qOzpxdIuuGaU7e3mO9kj13gR0WhEuAejFcPY+ACeSniVd0KIIFpGxwQoGlvN4
PQZZjubYHOGZsgO8B6pI7d6UWo35znaJV0KwGm+njolU2AC8Uh09GBLvZFA3vZl4Hrvy3J7QTPct
CwDOWHthQB5OR3dMN/7nzoo5mIWxyiBFvR++pNtZtR0FbcLG8QVGbpA0Ko0NFFKRjAPu1mOvbGpb
VqGgPLiTgoH9mD3LguBZMFzs1ZkxlgOkMhPssIYxJGIAFyp0TFkF/jN/THVCnqO+glSjdAozvFZ9
13O1d9CXpdtEZY+AkMJQXigAE5JleTrXK6NvemBbDq1eHe9G7txn6Al2zrvhdctGGM8d/Wy+sGA9
/8gcyFGKJvwEEi8m0unDquXs9hllzx4zwvQcJda0hNgGAoKk4rCHJnQYAXazC9lXnW3pcIuUCpkN
Pja0O1HCeLw+OYmD1DXBxMB2ehaUKk8UcrYEz7DNRShzr76Wi7I8jqJEetwxEN8fGNo0hGm0mT/N
bgJq5O36jNws7eM77P9Waqpmm9NYsFy7txgb7VnV8ObtYw+wHNUsxy8zDvktdv0NyXvZAQ6Iy5YL
hlCOCver7prIfL/hfpJbJ2GR1RzulTbDAD1xAAemFGNEWKENTkH9Ncln6p0Tb2o0rTR7ZDwWH0yd
jo22MRUN8D4M1XQiRDXKBXuwulJRMhPPokHVxS0YR3MOl3MbrJxEopKqow0X85+XmE71MMv87cIl
zCCrlKGSmZshOXAOvs+EEGW99/loY9hC39CTVQWKWbbHEezQwrQwSU/NZ3MSDFXIJHMVbcPlvmrO
RLfepanxleVi84TH547ErjbLvFUvrYUq9TBe5KzbtA74Fnibyu313qg35p8OxeECSWPtpRq8svM0
kEFBi/YSx/CWUFT9cNL2HxvFij17BftSrZx+0CG+nPZlPlthHvYlt7ADzQAHStbK9UsWzICeY+aW
0JkJKi8LrF9n7SNpMDplygpZo7xu5V3Z2AaKtDRkvf9LGH+XmxDblxmvHQFIA03SCqKhQPBGxLpg
IEMqOGAgtOmtfOoTfwEWXrZ3zPmSOiO3Xufj1I6EpZnUEiAkFujgLalZRI4XcTD32TWPJZ6uP0N4
tohZezaBIKsYTiQr8PgCBa39bK5JyCazH8J3j0EOTrhFy3mWq3GNWWux2DeGWZLScnTgKN8FkC8f
LTc3B0/JLuX++iszmbmZX8IkxrzS+c/hlAbIP5eifhml+MERFoeOfUem/x4jlbtKMiYv9te2md8B
15xapXpHkrRbRvRe1mM5M3+wLSRKTHU7GNUfCIBdKq35rA/NKv8Jrv9bepBbTo5J1kUA0ndZruWa
1z7SAJ6cvjJqwfweutm28yrf4duhOBfoM55QnowvzAqiRfogS/0mGMD76n2DX2ycT/75qHAAcPX5
PcfUXJcQDWuOVhxFZfMx2v20+gUDLO/eOKV5ORmux2alVLWxWvDkogDfvWaz1Njaw3FJBet0tOpY
Qm7uZvhL1024ya0NMYSpdOLdMz2nMynAIaObNvRHIbBu3kFTgBjDHwp3RY628nSZzKfeuejCg2T8
TCAYBU54jWLYiuwd3hLFxRPoHCFkNbdIzNQ8bc8Nkk2iD+nk675H7qLLsHXedzwKMj5l73mkIew/
vBpc7/SNmktYaFGfuvQHPGpG5fqTMzHjyJvYbKbwPnmBknS+8uP/9XSb08wlLMFCjQWO/WQIJHlf
KVsfzGlmK1JisZpR97a3hlwRR8em0j1dy3ztUY1A0NgxO8zdCV1Co8LFE3tyTd3R7nMUvkVHZbki
/saVhZw4NLM2vHd0QuXehFxwf8yTWzc3U6slaTuAUWjgd43zca7cAHzU+8bxBBMEs/W7uEmkfFJy
maKseNOSRwLBMBHRLp9H79vqPncUOXvn1ecI+mF+Y/iC/Oigps1jOPUg+5Ku387+UjHxUB0trcXJ
r4WRzQM4FHPyDicgotNa3MH0fZL8lRq4hTZ9LKtxqXUNVbmJ3LBkY37jMu2YYiH3NYfs+o+RJbJD
BkaY8/O2SGdbwN2BUkLM4htCr97eLj1LktNxcz0bvOGb6+gJce8XQ1gwDnb26UdC/5F286hqYRgS
FMO+Pz/7RaUv14l0iMvWwlG4WqYHndODbsGn+ug8vvDs4eJApJLcU9Kr1ZUBU3lH0UVoTd5yMae6
t37lP1mczLvBa8Og1LYjkuvTaS+UWZl5C90MqYMPhz5D6S3Owbx/9ZRMdyuYc0Qymv/WSga40/AC
quqDlOAzIUSRqJ1/pt1D9Qxngww6utQE6/IrQ9BaO+XPjQM4T2jdhQUBEjW5kY7MomZqRA5Z4ShX
j3VbOQOczwMnSwLqPOIUsxsqR+BlnCw4UHZxa6HKyp1I3aayOAU/xqab+iNR6wkJLgIP7zGKICyn
COhRFAgb7xCMZPVUlyDp1bVyDiOiSOJRC5mrPlbjUSpIZ4kRZtdkiH2BuD3U5NKEIFGTnBG8yeX2
g6Pbfl+cJk1Bc0Px+WQ7vxWnaMfDfp+mTU0Lrs7UBKsmbRI+QxcxFqinknODExwWqhEUFX49cnwB
L9UZRE5PAxjYW0MYKLGA5KfOAYoCjYEqutQ4JvI64QFQT2hdjPB5vOow15RaipAsABw7dZux6rpX
UCfBJBC2V1NSEPgT4RzCRvB1WOhkqNoe8l7Vxo1W6pn1XDMYrWD1RW0CZlabz3+7N8rISY1oX7zP
YEmYK627EQsqv8yDjX0IixOQlgnfg8C6QyRAIPdO+sMBrnTiapFA0zvPkMh1yZ9N8AKwJiHSab2x
GKyJhH3dWGCCszLDS8MzIB2wIbphf3zHHHrAjb1dCwkKS/6mF1s7O0xqEouRznNkYgGrjEcwjaO4
mHiQ6TBWtl2juwHf5vlVlfE6mjeiY3zucuyD/7eC4xGcDWVMqOfhey8c6m97W828+tdPEyzpYTDi
BehcUGpnpqcFoBMVOJISFW7cOtHq2Xopm0p9Rths5uPwvRDfOSAI1aaSVqX5q3e6Kvu7CPYe3PrX
Y5O0mtMk7jjJPnx953Is+Hc29FtQ8t8Sb5v4LVfkO/6i85KzFgCm4H4t6hOHDUE7DKtiuemGocVM
TdL3+DhCFPrEU+8yGnGJhSsO7pBOP7Vw5FGX0GSYYKDvPt0iFD6w4a3dPTel5AaUh8ygbZhE3Zcj
DmQRZBER4GD3pd7/5NtolFddGbcBfhRwWYNYbNcQW3UZc6EXS+5CLO1KJzBoeoYP3uSyO1fXsEe8
o+XqtMm4keMTH+tgZ5QVXJQwEQ1BY1ZpVIGkk0gwZrEG3Rfkv/uv2RSQ/nF6VPA4WuaJcFjhk3jU
hVeFErM7XMa2oEbgBorpHmdZMFXMeJKzUqcJz6tpnZryIqIE1WlUdeXCP6/WhgIX+nrvqSMMWoCJ
/eZw8h4o5x15AdrnAZ/WJpwYi87v/4cXkdiUMV5uC2bcWPjjJjYT8OBGxH5wtAU8r00d0Er7/TUp
i/3GQ9zGKqGBjaQwL9ry8Oi6Q7yAw83bdwynYjwF1GE3LORknL/CN1/yUxwUE+5QOUMIxpNicywz
viCUJYMQq9AICohUT8jUjfT+WOzVqAMYeg0EDsUE5ghGbzc+eN2zWgN3fznxp42qnuuPkbtmxlio
+SJwPEFyK8NjUrLn9nTCORfQcK2FF7sI3+qEDeyNrPXRTeIkCq6rHKZmmmaTg3s2Wskh7ng3p/Sq
4opvTgVkvYhB0htBT9vgkAX/hHhDq1zswPwUtdXW3/rQaPSW+vYFqaaZl8OypAudSmgX5zn8cqJQ
XG5D7VZ1TCcrEKkAhUOMvARkAWY9peIoa+KDfJ77raZoKxsO1m7ECLarvgH7h9+DjYoXPEH/IAzu
+jEM0Q+3qSpGUvUXIaV9LFEGLoWccDcS6beYMRESqASwfUUbD+V/ambTfOCnJTllwsq/hRkxJ/tG
6hXJRJIMQ7SDmLI+4QIueFAWohJSS/R0qE97ns+caIEVy6VNc9429AHvQ8rHNdGl6Aa46mUYJoF2
GBhVEZ2j/UDIbkVZensA+hOHkeBTrfjriMggo7RXQpX7+opdxztaMRdXCMKxuvCo+dYUUplTLVTT
2IdfScd+BB5l85CdMhWmuhiESzB9EhS4gyPhAjOi/1OxJMp7mU89dYU6Ebh1TLcaP2Hs5Az4M77J
lRtC+g7dB0p1gsGcC1qH1ZXRBM33otVpWEWNoP9nJ6q/ydLEaHO0mGP4J7bfUSZoTXQQKBqDO+bH
WHpzOi/2WzHznbXjp6StYuNp5fVNiFknrhzWYbzCzBHgUOphJqMKUa72Wv5tXsCzMTQW9zkEIo6I
UAN+1KeZAU8F673TuzXTV/LQl2IlqFUUF4KD4kf7FVSgftaLogPqJKmSDE6VsosVEdwspuQJEKXR
QQ5h8CD0wY0NG5qx+qZhKOA1SEUteiJTbsqyDY/UaCHRzgyvFpJqKRfLEQLca3557csX+pG52JuE
XpcgI/KYOalsz1l+nfrTWgamjm5wWSpXFn3cgOCIGcJzOEnlKiXW/AiGUjFDsOGSI7XEbCdmZ/+5
GiNVmOQg4u9Qw2AiRpiJWqSLS5UkHHUpI478el6A0Y/X+VJJN4LkAF73vdOIQ0cFONDVJ5mD82cl
Su3INdxGzu3FMK/G06D38zYQSu04Cm4XDRpVRinq+yzZJCiBozZs4ZC6H0o+AAtTAWWI7TJN/QQM
aSIMRvzmC395jrIGMzCLjtgktNU78TBVb2U4UtGoSCcyDl5r3QGKxYKSVbj3fGoJkYrwkut2jm8T
rw3l2qgh0kAJHheZmGoFWbVffq7d1lMO92T5kRXfKbj40M0yHZj30agKcSctaFRS438d87QLZC57
p0YwQPj1xcLUIGoy5FrtTtczpeZm3nVyB1/+PLKtnbaeqfMxirae96dccIKS0uOoqTVjcB51wvMR
MKDCXSuUQoCQgztkyC19fqta5NZe4cBi1eiuInlpzfSe3auVi9wrwdSu9t5Z9wuByqgsnu0yNMZv
z5VsbqrYwg6LPq5rEmrX8SjkqlXw400dtq5KXn9hszJhgOAHQPnmnzNuzC4gAkK3PfLj8IawLaCt
myy8I7NMNfrcujxrGcdpx9Zvb+wuwb+L+V+VvqJDHp8BJTsEO9NyrsXn6zG/xrjLBmTrlyp8KPix
dOIIZqL1kVSUliqz52It/G1TZvcwa4lrGJTyLgNVGxmNUAf+4gc0valO9pYI6wek551391xjeMqN
HLvtAZ5+dwkgmy6hclWjprkwkXbA5GwzfGVLtCq98WroxxSYt8gjOqQ+Ey2KmKaWvuF1l7N811lr
/jb1e8LzEsOv5ukbmZP5zy+ntV961sZtNIZicG+L9g/tP1YMHljv2fIvHdKQNL8vKkYqFgga02GG
HR6ZMURxh/gGDY8YVr19WKaLTBXysq40mSr75K3CxFdnmtrzcvfWknhB33WcOTuDMC2N/m1JgbEi
1PPQ4EtXuXVfImdJx53yfrh6tADtEQpkhIMhqPsUdt/OWo/mqrvKoyhtdZoVeCSKF+naVkBqWUtU
kOYb0FlSHxx313VahUhnCAX0dWtFAJARAQ0tyFfqSg/0XtCz5I4f/p7yuWYpRne9A9e4c6fj0pib
6S1J4dINTxogI355LhUselyQ3WlsQiTJ7ZhLsTOMcS2360Hv4sc0RIJyUZgXXbQp2Qo8ighDcj5/
664ZomUos3/MQ/eBmyzRWJrHTj70GPbhMGW1AfTcfPeEbbaDFDvxnp2GNx6AtstW24QbVawOer9d
U5nl/WIdlwTj2gXho5Z6RtibnCs6hTKvifFzElAnLItIY6CZYt2HEu+w99l8Uuqa6JyAk8hUWcZP
dDSHl9ptnMBbOJ3czAkFdvxkoH32kqFmYw+N7nuEozbGRk/SJfyaxvGnJg4gUHZnwvuUIBta1hIV
T4uxJjgmyLz5z3a7i2h09sFtgjRbyzsaf8pny7cWasovkmjGS2qH/uK1k3NwM3pJKVFYMY9oLTva
XUVWwxYZyAPIo+ew+juhj6oeoRNChkXMmaMNpijghnNIbnlEJNDH46+I6ncsLmLAJVmfCk6GbAwf
Ek5eL+XV4PU7WzcfLMWGgViWwW5UNsCL/M0jWRgn4FJK0ECIXTLl1moRLft/7pkk1XcNmHF491yw
hj5QX1aeadiwvDNZ28voyS6beavfhlBeQg9V+xpRrUIRHc5Y+U59nHGKMRkERVrgRFmds1ssTv5u
dKIzjjUtRRvYnoQNN1XO9+Y8xOLQRF3hIfOqzanC2m3treJl0S27GTANfXVaK+vMwlL3MIqejTA7
lj6MfFcAaeg1s71ZjUNGRIPKoJN1zv4YuETJZa6jyny8ZH0+ucOqSioYLZHslfGLHAVk9jL70lss
miX1g61erzTpaJZlQynUPShpE63NuacdgXpeQJaLdaEGkaqhkbRTqLlbVpi3zXweb/pcRANmxdW4
WjiLzsEi/fD0bH+ZRFPN3pBAzjOwISONmX7b4RxxHiHpyEGaf4v9lUXeH1gA+RtC5WulVhDIkFl+
FMvwsrEqKHY3chkZeamKM4VyQnRBFtEedsY1ruo455gWbB+/4ae9epWB3LdtnlMr9Rjd8/2HQ6gH
uBuT3TpwJQTQtlUBXlkS/hd6vNIjcxioaq9wJOritMAGSnTnBhaENqc3MDtuies2WU3vCH+H3TwX
p4MAAvcOO1ZycaB5xbALYxIqFqMF3G3XyMpipcH/h/6REPVYlJ89pBNFpteosy3Y1xWv+5V7jYDK
VOZwoSP7aPR/BAqxn5yh8CkJOe3IMeQgdzDHwhAohR4oHZn1QbVcmdzfAbaT+y4FQFz0thAlOVw1
C0ReloF2nmqg7jX9msQTO3v8rVt9UzjDEbohkKSOxplxtSRDOLWaFlb7973k+NwRC1QAYf68y5MU
L2wbprYr/ET+aATc7i4tn6ZjWeu4I7KIClrjCn71p/61STi41Q8WLyyMBEVji12NOq3to/k8gSjn
vTv5R4L/MT6E7X9MLIjC3oq7EcgruWmEmBx+/A3VYDcLKid4hUYHCDXlhmUhtrMCist+ppGwH13e
veZseC86gL47YlXA+S2oFX/zlQ6GefdGxA2tWh7yZSldwxTeZSWe4ZvqgX8tVGagF3bpmfXuvrlU
aAB8tpeNrBZxliwzwKGsW+hiV8yWyb1uHWLQpyQ0WKSJ0oHF7tiNqQmXaNip6N/NJ5WbXhRitHAr
6Z7nuSK/f3oWTCOoN+fsIsTMcIFClwgNA4tY3uN5fF7WV8W/xK/xBXEi5P/Ir828cLoT3c2rWQnf
RdV8NeoDvQIVp/gar1gIQYSL8L4h0yW2HctbDt8xhZqadAnz1I3vmjW4HfX2yTE0tcJY3Qm1TnnZ
mvre8Xv8MJ7K35NirPvxMuk+P2TamE/EMW0JXcFAk1hHF+LrsYaSQ8AeBY+uyJadC6IJbFm4S0s7
A3CD4zDdR2NnUTtediqXZ61HfTCBDUNwABU8NLxmXlTuvB7g2sKzchLqtSCy2fh7VtK9EUkT96e0
UDnKOWgh32kCjKWkvyoNHeUVA6MmJK8uRQ5NJyDxmjvx5xfwy4s8370+CtVS8A4XkhTcbjsnspW5
U1tyuRuFjYVmdz/aCYXt/HTDkQ20tDzJAs/wZVMuULeMLsm1orNv9HNnbVUsQZSRN/ZCR8B/MsH8
c0joUkiwmiYDyOPXdwsEc+54VCPz1+jIcTcb+e5JmKX9MVMu0Jab0ypptK+mZruG4CpTRZA1yPlY
v3P5Of1+KrhJVgZwTAJhpwpQ+gLw2qiRNaAMC0a+i1A4LnY8ubTyOeC7JlG7HM+5QOZY9D93yVub
u7oQgmGjPc2SXL7hE9yWZQAvGxb8GzPEwyapJTBpyFBZmOUSijsWDKyqbsMeVVqQKcanujvVxAvv
djQTPoRWu5rBKX4Bu/07n7uWmUtGYLAwFFysc9eWFA55LG4eo/XZZCFWwWV0rF9LsIAfhR48IVoo
SRyAzRux+Z8vG4yEuY2SKsh8EuA92sDSm3x7X778i0E+yETUk/zPkO9TxsGDFslW3Q0X9NeNRojN
hdgz1RSZz6yzRA3g2zDSFDZY8ZrRA2W1DxjISlVINsqpoAA53ehgCo1AV31R2P27kzkf7znwRuJK
w6fd74fW5gCvxqolyXdmmb8vBT5cwMTmyWfStKQ1c3atOquWIsnQWfQTLt6VGrhk+IrA40jPl3wo
qE3hDxM5pkkOOa5vzNvDBcavZD+1C2mwOtAIgKTp7yYMN25nDriQGDXQo81wb40JC9ml3FVGnf4/
/gHB5B9eLdDpfL43URmc7iaA2BfPukVQI1lV4dZkXfClAn0gsTgzUEUCzeBIyW01ZYpppnuIiRHU
RyYVOG3Mi8D7ydjmdmXOewKHbQur2+GtVhWgRpmyI6V2uUz9/s9UPxZiwGQmoCPsZZvgGVpQCIW1
wbvFYoWl1BBhlE9zEPSxhhsnzJG4AlKlwyGU3CLDGMDvyNnXO9b+AuUiZEmrpZmYww+7MOuZmGjM
ok8pPQNAgW1W7nTAc4wxonrrsRWRXLaj3XbAh8wwFsNkpseJF4gEx0BeTgilC9tD+O4LG4aFgAty
62fTEdro9oPsMUQ+7/1Pjlhz1VD2A0tQcztaOZIB2JN3U2gRbJ6jadON6chWKV8t7//NT4qoyy2T
vH8LAWwBmER2aEudjvI+cqcdnv7llocJ3RYjqG6khlY2Bcvgeb8z/V0cxWBYikvflqIQj4XiYvfT
nrCmlwkDGVM8AC7aiXY9yga/ge85jUsY8s5yeqUuCvhW3m8L7WBXOCLKd5gggVf7/QwM5ffInyXb
kFdnPhbo1792Ih6jFXSz60UXadjhJtrDtR0UvZZH0SGQl+nKciKB+WZ3I7LYoCSLxLXqM2eWoQ2q
9rcFIBdSkyDPrVzfQYx68T9XoY6Fkm7ct1J0cUEFUl2uuXaEYQeEw6WkxJccHLX40feIEKpBsTXD
D0Pc143yhkqGuHS5zrQ1A4RVN4WcnEEOSb76mi9iEHb/oXcXsYopbvEHrHRy3HTDqEITqc8koJ92
eGtIVYdUt7/zznsY1P6oH9Q26oiQ3/kctqOn9x/FBDOYeeSiRbW/YVKiVYYM4F0ufRJGMSmZDAfV
q0iwQHK2dcOlrErYZ8ZPzcFKikKLCS9pI2+bJY6yNOcSRpaXJyNsRZJoYT5GGkLW2V67+oCwiEWO
Q2PCKn7QxEC+zecLHLjE/v7W/Pvtu++x3OEqMP8vAPDygefcdOMRVMrUIaUJFxF4q2JNdZB2ZVYl
4sDSBsrUxebqptPbtTbBvcL9bFoiWnH93sdBVXc8hmEJ12E1/wnk1KNCX+/Y+NYAh0mLHBGrRkIy
NPGppSmXUJP8BSBuyXl+xXlT4ggfTTGDKB9I5t7MMT9ebFUaGeMEpx1MvpS1RuN4GRdpolhA3nZP
oZqwuN9I7pOd4uMU0quLgOHi+MAsyWNJJrzJVX7YGfbZmRJOnwhfGu82Dl6JvmMwrEYnt5p5dT1m
lt8i7GRmSJu0wVD9nW6xa1LD7CyIimm+PbHjH7AGSNMWtBGFQ3cW2Btz8M5713ypyk+lB2AzqG85
mNamFerIqa6gaysHEgCtQpC+qQOEt3Nh+1UWr7v5MKphJy2mVYoVYjKJK5q0GtPRVOvisGpmrH45
Dm1QMUsGqUJa3lTDt3ghlMtoBDeKw7Ep/LI1wGymUgbg8h6pRoZgWfXmF3CowY3AWXnC/6gL1lmk
A/nw9I3uUR8sCLuH4xEiL7FZnmDGY/PAvucrlEH/6JUxSp6eNkZvvn9NwImH+EcaNNvBT46uuSrl
OAwAH4+qsHxT4WzjalrMwK3XAvtiOaXMlX84Qn7GysZxDxQXFVkAznM94C9hojTmg2So31MpKsVZ
dmx/F3wPXR48G8aksMG4xMk+PLKiV0VU7nn7CruDTEEYNDArTJBUovxMXczAJnpX8bKm2yGGIGhx
k8UW9Y5IzlLtS94FiXW7YdMmxOp+/cdnlIoRsti7Ng3tsw7OJ+1Ugwak5hGiZYCKIwVMeE92GNwv
tlS/NKO+dz5TeDLZUL5GOpOxOJ5ZKkUEBkhWQ/Ni1Y2XmnQ1PZWWQDjGVqR+gLo1ktVzF3qL5avV
oy5F+WllieORSalVhfyvhjTLLFbQ9HuxRIU7YMJfM7yknfQKjCsmmhCXqcEIgCqlo2q+LnqbLCJL
G9JSafhk2M1bHg/hTriFZIeYMM6OU1dF1JacuDL52q+KF0sA5Crnnsg0trx1gEhvJmhKvZvb+Fpe
+W0PNtoLvtpfm0fpYRf2/zHqQT2BahWWHJkdlJZFlNkkQJcTJ0A5t+VwZDgZUd24UiAkIChMX5Q9
DaeyAV5VXBO+s88Eu4Bye4y5JBC/lFAbpRJ/mQeR2PnFH+nYUMV2bShgjpieVLsRL+AODcS53kco
XBWbYDJaPxH1Vc0TCzuYlTLin04p0VIYNn5ZEx/sB8zv2mgPTCD1R4atNLSZY4Z9uLwPC5M/81Wu
7FOwLqmyTa0qfLwifobPpLqNHsT3dIB1RFe3yrNtcBUxP05AyZs8ek1AUZvuIEIY2dD5gTj5r7zK
Vr8d9vWDGVy8irD5XNjA1OWzccFRom+2OzuUe2xIcEHICEy7aRC1sJy7VLXsPI+f63WuoQkY6VZd
qmw6fFn6VNSFbyAgMEznmtYFfrbTsP4zFY0y3EtcXb4ByT/xmJuX4NoPXuN1KvLzfacZcpJ5NXft
QqwGlGcuVaLgccMA+OCOtaHUcgZKNbxL0DWCsUnSGeX8V18YA/JilQlhgaYMsGzSpxH6AMBPr6jb
kgIJkTG/GQ6fXr/ytbIPV+05jKwnDP2e4WATx/Ynj58Rk0BZTv2DBSJIHRrrE7yDy/q/Wo73G4vH
zLtsOaSZYcNwq/VNPaEwXry+87SfmH8Ms+crkuKHX+vB4tDLZd+SC1T4qQnyvwZJz9uKiiZGO+Ho
7+XtNWCpppsCv8FE6PnbJY0LDBes/xWGCsCYQWsizTEahJdaGFW7zqJhV7rUm5fCkl7APplzIw8W
2maHJQAyBqvZNjMd9RLZoLQKTRyU0hETP8RG4GIZ9w+LeZx6OHLK15DSv77VxOW/3JpJiqrduh/N
hBslly7e0vxOTJCuKN/12hE7WX9ZIIuJuDBLux/1vU7rlObmDr5XjXB4X/C00Swx8y3FFqs2UR2n
wDh6QlcSFpa+xzSPz61KGzg/DxpKpmZShqezwe2Ha9Fi/61L/7AyQYGMJHLlsfx1esYt5GNlv/gs
FoVfOSVL7MsyCDXlf3eOrT0Smr4ystxJu3w8+khlV6KPUxe+YzqtZlfEdXgnnddLtIJHYkZxxY7G
+8kTmOSpvd6UHC1n4+RXOkA09rvC+lczQc2SsQ7HVp4yFw26KtruoZWPRHcXvrFoWJGrM3R89gPl
2nHib1rG2PubQh2YNNSCaj3dHpv2N2IjG8MBLROVf+itK6pcyCcAmNWwtI8TjsN5A24BoZjtDPeS
dkLiAtQ3aV+povbWNE207P8AAehsDajlf2rAXD3D5V5A0Ymyn9q3iKpraF5Pr+xSRY9ivND8lhaT
SbN6Zp8SS4PwP6UddRvwlrrOjypnhw36Ewq4LmWts7C/6uGyU3DMat+kvYTajNylivu89WimyIQQ
NYLGjBVi9QCvAq3Y9i/TFg9UqA/kId/MvhOhRvNGUEuUUTMbOgqB30RLMjpWBdVMZyNax7bubE7U
POdhXrS0pKr7T+1rTlssjjaEVcq10cZpHF6bgjCIISEeh/8FyyhrXcMkOyHNdJj4u/ug35CT2qsl
lOKMqQH0VeX+rId/dCqsor0Vc6A8DvEdIbpUJXlZVpnEUGBX4zCH4XN9Km3gaaposAGzpZLDN50a
K5vG3iYhWSDx3g8gQfAYko8nmtCI9qQchzrJXBPx+XtoU7PIXWUJf8gOegTVYeDDg3XJwzyAW3sH
GLvVsSHJ8YF7J3c9qa2Z2kKMdOLezMwvF+u9g//sjPlTIzd3IpKegvac4TAfe3ZHdtDu8Bvbt8Bo
I15WJzkYya69xNX9ZFWu21XWl6Tc8ZUH6vzpT8h3C8ngnPCdR6gy0tsrMhxsxiqW0eJMRgxsC3Ox
3P3o4OSJq8Z2t1X20Xg+9uNLXa5RncXRyFw6O7A5Yfr3agz0e3DM6zvFQO6V/tpLJ21dy/jcshuR
fd3b5nP6EsoXyYg4POKidcx56Up+S85+8vGhwSdwidtHfvHdXUj2UhXsE48FBsqY8e4Mi3c1Tteh
+D7mqkY+QlFxNZ84JOK6lCxBlFAQxMN0pgzFGsa8ta2pNbSILIsxAhNu9UsEy3g/NXhVl4rD0OSn
jM90pXgfi/ZC/jAFvYSS11kw4BlXIpVQ5jBVGNPmsAcw8qAJsJeVx/0lbsI8Lc5HfQvQOCsb2SbN
99ofvDnV7wJoR9DaNvVoq6w0GXrMVanYbzs2b8yXL3+V0tz7EYLWPbO9OYvcgKPznEQW/TMrd6qR
ude6igq4/PCsUHC/gFWDfHXcAOYGK0k6m5FBdK56BKScL57ijFnd3yJsDxaQZOH1gX9ip0QCiGl1
ayiV8aMjgekNzPu4qgTGv7iqvJQlJX8HHtXjdjjTuFpgFnpeWqy4jPrkMjB2L1VXLIBhKQ9t7Axg
E6zXlLDXq3ZDCpf+W0gDWsLimg5DMNiDEpMWLNzaYFTUgGgFmpOayZNa/cStAZjuNV9DKld2IeQ4
GMAI4paF4rp8sLjbccPL89OjkoAmU4gKXAKV0Nb+j+xNOFcCE8Tm8ewA6NxjTOfn8XImIJX8HmmM
m5V0niecms3IFWRBBsROYg8WyX9IX/T7k6+l9reDULyU3CgBIPTDe0UQD4sdAE/ZL5hgld/V4WDE
gtQrH+7AGzjqlbWrr7VQNREhir5PTsuBO+iPw0NFG7E4QDcvnogXBIb2gF0A00aq08Z94c4GQRmL
oM2ALIZ0kwe3IqSUBfvco8IO50xXsZbhxYn8ygWsLs595pY8iP8pPUhMEv50xjKyvekcnqF5jN5J
W0603UsPbpVY5lV2v4mlD6IByAFOIV6iq8a4Uldf+tAPEpaDmSjdSI7wU2je4itUVwDH46KPMCMs
R+CS+e308hxdGbcp1aZDHm+Cg0ZTS8pit0Qhw55dLYg3OpqdIoVMu6saXTkfinAugTR2AQARaK80
WdE9E/FytioJkvWsqPWlu7wTSYnF5mdXbk4BuOr1BAFV3xANWWao8YGOzcb26yDj0ikFQ5QR0Im2
P7Q6OW2qQonGXfbiR3AltnG2iH5SN6QvJspTgXoC88TWQjKdnpXUtuEmlcUjgt15/gG4n92hxIVb
6NZE6dNUB01jjktZAoOpx+n6EBtYOUuxZJVufpmV2XQSzki0EPflzz7q695I8NVW+xx6y8HCfXXz
vVnBVSk3uVnyVaWZG5UhgPRfPg+KtMZDba4YqJkV0ugCxE+080rfYBUOQ0k5h7xUdSJKKky8CZuE
XHbA1plIxyXMyx2QY5YUyATCvPcO1ihlDd7G8GxoiBi57etoVHm1H7aLtucqhWSu5Pz3zYmWkxKv
LVWUgF1FZbrK47QHomlRGchKjUkQ8yVCzOS79enhbg16MEQyne/2U8KkooHoVx76c10UtWyoYxW+
AMeUvJbt/3uwdDvn0OTH1xjLZ2fKcuzbtVAVqdYBRKgz9RkplxoOgIj2BxJgHcCdM8hVjaFY3qUe
GmHjzmYJRfHE1feRS3OMuZmoECPVba4r0K6L94k6M8VArgDSwwIKwmO1QIxd5KQDcQXWAX5rAdsa
L4GuYyw59+Fsb5VUmKYfR2YHzrSYjik3eRZGhyYSFNJDtpGCgZVSromWZpNgt25A0lYM8lkZ179f
JaZJpezg/1gM4a9Peth+Eg6j11WFOfLi1UeQuNj93Fk50OJxISYmQN4kQrd6uiPCkvQooMmRS+pI
8Uk4P3LYuFlUoHGC1VbeN+tQ2+k9jRsvteVkamqyQO/L0V+mEhcnBh7fDYLm1m8VVCwwEtMiTIOW
8AZgmx0EVLTCz4x6BX4DM15IvJMugQJa5sIDwV67cNQCOUpjGsPpnAY40YYOyUl74elkiejO7hV3
FWfdpU8CL9vdK7ToN0aUpIvnxIapJS1LLZMRWEgLkJgCbcLG3ODU/bc7k6FVoGYu4j7FFglcwxSA
46VfO3iV2I9yQuxGfDbKnTV1Fok6kniX+xcWaRY+sFaCkzq9EhM87KM6Gmf+Zx+w2W8CzRQ6kDW4
RokSP5ETtA/5hpFrlHKzTlB6g47jBqf22rc1EpupPKIzZsaoVaMwLTGZp1eSKFbMO2BHJUY5FbLQ
myvGaoZUTVbosVvwb16blpoihTyYtzG49ZpIJZeBiZ5HEQIoAfzN+lREWq+RTFca3KOC0RNeBPT0
ddE+fy+gUC0iCiNQ+ChjirOdPYWFDwGjCXr2Jqu32FQ8Q3/zbETcU7msGk4xSOlYYq07r3PalbM6
mtxezJVKhEOyzl4ohVAzIdNLFZUIqjqzvWU7AIzAmnwn8VXNto3IAK7PkW0xasKwFCF9yE1JPVIv
00gtTpN8J2fjvmwkwGp0SnMZG9XLJ1c2lUY3Kd/7yTtjO+InTouu84FL1XWSsUWOrZP8uxh+DYLP
BlcQgO1lUcSEfF8tfG37ARKWHNZP8fJvZT45+ZnVWMrp2l2YaVf8H4/T95jmUeeSG50hgV/ApDkG
BJhp/otmdNJSIDnTKQnYk6PcIx9jAou+Mpp7BwMdt7gjTxww8HpKbFwDiE33XfqLXLnmi/mr8dWL
wRWdjVbQxkLkw4V8f2O/ws46oOtIFR+XWIVa9D9wvXV64ghQAMY92Y8fYW5FpHIAomoUBW71gkqh
HXqMQSMSi3CUpD1LkCc14gVwSyRfl7JCmKZGq9oQB+Kioga9oxj0Q4HJoGLtbX1ABItmayFQURbh
4hlXRaJXpzMsd1vgphYpFxX9vcSWlZOeUFhvKyPwxG8ldunjgxmQhv9HgnxXRhzdubM6dVdVbI57
DepZoZnRfX83LkacR5ynf3nO7iKwnV94i6tHKDGWbzhBekCPlwEI+8Ga+I4NUSEHTrhwk0ZTsIKF
cgUedhBjYrKNn7dbaKY5Fv02dAVt+6CMtPJnjKI4GJpSQDKW5BjCFEb+CFGCNMiXfiAs1IOyxtXj
G6oXO9rJr+xnijYlwYYAa7XpLRGPYE3g7V/cHZOZ2GqEcrORQA1lsK1bhY+BVyNPUJQDfuqj06en
76BRKV19YjXJ0eIHEJYVKoACEFERkGRjJZnbCP9HQrkEqOu/EYZPCxDkWW5po290Ivy0Drcv2cGA
K/AFhVr82Sg4XvnuIcFrajDpQWFsaGd/JHTC9C+QzwJdxxdoDbwwaKTTepSmNeVWTHadQJUjW3h6
q5NY+XWzBwu61UBQYnN2Svyi/7WN3e4DHgpUk6+cew7pilNO43/W3O50rsTg7FPTRj+q9qaxCkX3
CH3nlcoEe6fT9OQftnGpy7lAFbZLetdmk2fnTKOM6YcKXvnR8OfB1+CNyl3yhlP3ov5wSdDUyV/Y
biPh5dL1N8kuJmjgH//EmLKGI5g2mEvkfrUTprua8G1t3SFASabqWJFf56hieaGxU0SMHD+SL1bL
FRqGtP5Yix8kHj63OEIw919uMR0gQDahPnOZF4Nhjkiyo9ZEFCDuyPWUEaLggb2Mm5ATRmpX5B1S
kevTMSO9Yn3VaQWPxpsx167GidifukjxIwEebI6HLfmVxMzsC5T+ylXOHgH4lbXN7q9BBtf0dnyD
1vfTPfFcxC9YXeK+YSSjsMUy4DMdV/M/Ksqr3pofAsmlvQD9vuw6x4tKytCB5v7R3S2isDrpKG9t
i4/4PF+VSD/ieQ4hPL78RTsgcFv1VkhRqpP3Fd7zCyK050L58WXBrx10Jhf+MvRDZk9sAoQjHjnM
JIiOFgOdsE6RENp9sGOg3yJYZDYNjbQP9ndCI1qPz6mBgZtHsjEr0nQxynq6vPunoBK4AIfgtOYr
/tCSk2RH6Xa5BkI9XK1Tr9vHUZ4hizlHbKu/o+V6YB2dLfPHKnSEW5Ukeg97Hh4sVo/6nG58QOwf
geciEH32BiRm6RGYe6gWVlsWtdpPChJ6WifIzzn2yhZS7Of1pR/2NW0cY30tOY83kjrTeQGdvZHe
vlK6ZvVEkteXn/wkPNoj6F6WrhgiJmLr8LRkQf+7ugihM0vosTLRQAqvxb0i8TEtYM3dL3Y4iwTn
3dJoicvMw91vwr18+aY3orZ1OuDSOE/vqPG9RODpvN04Ojml8aiwsqjvF5VzbLEX1y3MvUWy1bFr
J4fviRgD6YQGsjAuCKdM5orndvUCXnrkggoOpAGjgaRu6U81zegV+vXn9D5qYiJbO7ruCOHkZ3OV
W+r6uiD0hof+NKidPpqMybq+dvODsbP/T5iA0rdZqeq1v1bLZc1IchTvDLoPkqPwbiEoOlPG3TEf
BnwyrUETw6PBMfvh1YFQwUUDoXimq8jmyBVkeEiYQm6GfVK2VLhsw+3hR+pbVDNyh4pbEBRzTJMU
nwgsTW7H3eiuM0xAaSOFj6BoP05g61J1d8kJCI2yBzgnBqnXDw8ZdV0Spa3g7nGGOYq0naO4LdJ9
1YcvnXv39nPtnIm3qAubAjnzUDWGQcSjFZEsJtg4AJVsOcbHuOi9KHY2DKY1DaiDx7c6AFq5yDoC
L3dP8JZ5GvWSX1vJ5yqvDo1HPvPqsaSSBNWWmRZ9wDdllWRayQ4DZkH7/P3m09f2gAJSmZ9fAfPJ
W4Glo8YpCjFj8agrvYTplzxWNZNXIMk0LSLQUoS9sW0x+nnnal0Ttv4YGsrquEmanuBI2WJ5CauQ
fgrxTVyMZJvMczZan8ipqZJd5jPmKvFXy5x4D0re+E36LFUEJuNajgCUI9At+9tOVX1fb6GvxLmE
HdnopWUEk8W59jJ+9FEDBy31R+PPOyKNqkRHtpWw0SHtPSKlFHL5ldOkvb8YZG7BPB0Cj9Q3BZ5L
MbTiCfSTBaCuqEtMRhkLctvtcpI0oefEWOPPN3SaUuYjQaSA34GXDC+XxnFOHHnq1yZ6W3uk2pqI
S5x6I8KMuz5P0vw+qnNjfy9qra0R9VdtGR9OfmcM2eN8CoZ0Qz5mDcyA36Dz6xPMcRovKIeBjSs2
se6ZlLZxxsXsTYgaaoLWc89IhCJI+W8D2jbMBMDuLvDXqAxckoHR/IBRGjCX5j0KsOetudUiC3VK
f6dzNtmgyn8+lS01xH/IvVfopMWzGcz6wduwiMIdjolQ/n41PmcwuJAi1dehn5aqbJYa1kg9dH/4
pK1YwsVDq81c56/cEKg7boCIBrtc5jl7EA49znystxnAL0uWVPQQl9HKBEdccDV33HA2aR9btr5W
vROkmJmF/hS2RIpWVqgx5OpJw8MghyzSv38k4pWKqoGH3I4gzV1ORAVMZzNEB1U0xSfy9IwiW7Ha
J5XzDiS4KrTP2HS2OEEkKMLsiXo2bDzZSd4QYHBRkgLsKmDvYBd46/JrC6WvcZF+m3sgNqU43CC4
7wSBAELh0JUO5zQGKsnyRGPNOurXbBgLmVjksUXKcWcSvnDBz2d0XTYLVUVjwtY3yK8R+UTlNKTi
0y592GmxPElUwxsOb+N+KTp/chOS6/886cGgQFQoX6DM/srG0POVtNA8Bj+URSUxUcU6XVdvwL99
RaJoNKyecx00b+wmddg47jaYSNtJPslJoVqOqSFowsvNRBenCFg4YE7On03ieeTdFLUskik45WL2
CzKUM6z0HblNIKAU8RxoH5iZGLhM8knUhFIfLXtCY0CaCif2KAdnzExlfxQ8n8I+yPJs/J9W2CkE
yd9Hyl6JD6q7Fb6n/EzSc+yo6/GGA1DWbmBoLkoCW8kMTLTE83/S+lt0DCmpcphobE2lnKO/LxO+
oRpcnKU+8mNjtgt+6U7UdHOFV62SN5kPaLwnUjViwB/yxeV0HhFXpeSu4ASA5TEOCAWS+UE9gHl/
8HA2uU3hKhWtgLS+46RazZ7X+SzesJ7mJIl+xNk1rT+8ifJNNaLMk4BpGb1WXvUBwYtyxhyx7/DX
4G5fuVPYo5Pr4jz4xohfv0m6kQsdV0mYiHwlqvWZ8oRnnSuK96WKKDxU/mbG2AiZMhuvJGDWdevg
Ly1CwxfSoC1g0QA/wxYXOoWA3/C0B3vFuLoUK2BX7mcM3d7kbJ7tinLGcVN9ksLifUyZd/8qm0cm
PcxNootHyeu2cPaCIhVHi3wXLDVM0BrpR4NQlFC4UDVbvDsTSNSaf93olOaQCn2jsI8ExUOacs79
sadquEZvwhDvwZ/50lWE74JQ5L8cYYBspeNZQhuHyMc0KcGuO+my6n2WrqAtRY19UMv3NQO8sACc
hpkLw04aptI9WiTkgAaM10/TkfnQyX5tvUEBH2uMOt6K95O9eNznALZAL57xjhk/T1BlhHIkaJN7
k55pr9e0e3fSF7CazVpJz3hjavPQt1M6BL4Zm1Ji23h1USgrKr2UJ2hFlKY5x7HlINcbb/18vMvU
1+2vw/1a/2HL1Z+/WGr9urii11ogpfZFRhyqYrZT8ErXEuX2YcrW/SA45LzeUF4PgwA+2xCefscW
V9YdidpCnNioEXanCQC1087Q3Ui8y+GvPHzfpOVdTch2s7QplPbpKUSHVPr2nxyt/u7rqIMF7Ttj
bP+snFzA+g5iiF5rndHkQYqwEl6o9MdfLF1/JmEHvIl5T18Ex+WXxXgjYpZ061hkHq+j2uMi3SVz
3vSqHA2vbLOWRtGjPSCL/Gw4vqaKYUn5Ml2m8/33UXy3+rHLtdd/pOHlwT+hedpoE8cRMFyZHkCs
uAuVbjLZkcHxqxUIKZJnzFYtex4EuhQlQacxd/1YxdlBZVlXeFwo+hJzKIE7VkbnhivxohqOymQL
KNRaxrNcwFDYT4xk2Ha7gBBOe8yIFhIl/NejUKLDQd7tkLhylsPV3EUPx7oE8H/T9BJxy4n4yryM
8efJVhI2GjFm4/KadtEnkBqYDqrhaTir4BiXbmF+NKPkV3UDQOZ9L3fSu/+J2BMhRiFzMEdJxtee
olSw1/qiBuLFVOGIO4F3pZZz5cnnGkHLtOTWw7qRqLRvAyxfu72ObPDqZk+OqYFtt1Pdjj8O3f3R
HiIPtksa8dawt+yMRA0aJL3/UZs5SQNncjlDlxBERqNiNNgKP4s9mYL2/bxEQNjWUUccmgvdtf7c
01WoVI0zye8GJ1kZEhnERePFaWWfC4FatIOczdgkhRNGVusIbcjsMrOHIi5uZoq9GdZUBSSoCv04
tGxzNu43twaVWF2uFb1ORyACFZCQ3ThRaniN9kd8yNOsms07TawedoBai24ugutLmGvzIkSdvaic
LgohhzaL7D6kU0+M217RHuqO72ePog5i5Qb/YnsyqCpI84c441Mw08Ol7REC1GwKu4IrSJp3FiEw
w2T3ksnCvnYj8n6+/14P3xAXeAhfX8xaeuIOOSOwKnzinPRN97llmy4ppTixmTfq1qydgVXgwQms
svnUsf+Y1rzYUPuhryfdFeTITKjl0H5xOpZAy0ORdcJVqmomtJTSSO8RXb1CKQb+1j459pJbpwCy
TV25BLiyhVa2wykDa5TNpGxkNJcueZM2GuKo42fYXA6F4KiDcItqAhhKyzZCKVslvdlqGTrDIOHr
lZpyNSRtiyTet+m/jYofSfB3UiB1GfPTuMW0wIBDhbuQiDYQUl9jGPRQghKJOhe5L9Qn6Qt85lrx
7I1l23hYO7QPROjNEILgVSJlToski7R2sDSCZonzn3jaoPsrWO8XBqEl1bIL6b0u6yt5XgMGBwh+
7IGs7VzADuIYtBP8fs1vVhjrEzzYtEf+Yl6o2MFdIBASOgzk3uRadQ6qmOqaVuaeCzKvuUrKyNgf
EVtqJcuDDyFNlG2h4a4hDgIaazSfENYVrslkGq8rvOhBLvIWFlUsW6AfUW7QUSRntQy/XR67kt5J
mP6nYWEadKz+MvUW9n7tfUHhIMkxUThixu0wG/tHnJJh27y4PWmP9lDK8SpmLBixki6jukj5mXrS
IkLAiAVJ59JNc4tK6f074+19S/UEeEgQiPHNGCKrM9xBNEss/cplS9QpRvKOBKOzF1S8eJABpCCx
AhpzaUWnAhWBKhM/nOQXP00G0z1T9Y41uj0oKKK084+Gc1Iq4m+uxqhpiLso3izfGqVRUYkFwgwf
VjMOIVisM6jM7Ng0UUKH2bQ0WRdJurrIcKcqWeIjAz7Xdh9PqcNeqAqMlbfVgQ7GTB8rMgjByZfu
/UlDP0HZhcmf2iTsWkclthTfWn9SyWkpimrXc8OacarHkXrQ7AaeFY1AJKtwYqpNNVrTXqHi7Z9C
+5QovxSGBPlqRRcg8tkizYSnfVyM24dJ7i+93ueW6sPs4ufwYFiq+HoRwnsx8HWYnXE5uq/KdReU
6YSpTsbeL0KtlZ7AWT0ilZi3UDTzlEVTZE5w8JwQxM1niMAd6HDluwcIRlJ9C8eADFg1B+gPvira
fMQDwV+WTkmq4rgCwUzlbZDonlKBlpwt7j45HWoed2PU159AX9QqK8uC9vY2joMJmHy2jaeMcmyg
8RqyW0Rtvq8BEovCjMG2P/Snf+RUMmRvs6S+wZZAUz6ViSOvt7dN/PsfhKH2ihueOxCaRPSwhI+P
94/xArDS6FabZwS3H3WDPM1pWHcQFGLwSfK9zmF9WFiMZAp4keGelQWiNepfRrNNU+u1uorZlBtg
MfGr+mYNCxt2qKJAsAnS2NEOmImpaBd8SpOZ/arOYfa70vstsL6rLZSXqwuD6sxhBJmv8vXVW2SN
/35DTHdsjG1ZOqJf3h9whOs2mEXQ6hOJ/fY7815wZYmN/vc2re6PvqF+4SyFe1T+ZkH0GNFYR74u
iGr61fzxWIumUucYT1e4A7a1yLC0ylqZ4Z19gBBUK+o+WRCBA/QQp1Te81kjPEz5av0DGL4clcd1
SPr+5jwmf6vXoUibwTasoiy7cIZvMJIeWX7J75LfcDT3NxJbaPMF/huv+/4i+LOysqQTRW8hR6on
j4koz0PEtITF+hRv0fwWJ1Qo32Or9a+rQ+jsyFvVYmz214m8zU827k4Oa392CYPwpTsouNTiQ8r9
GgVWapvE7pMarjUO0oBp+VtqyyCYxG4XB8n/HMMOyNfyfIb7slHDeUp0j9F33PSIUpzpkjSQ1/+2
aUr7Qr+PLk/i2dAk4wvbpgezfAE8wMCZa8cGfrUWtyDPdTttQ5z4Mf54BLsLcedxwkg0C/o+Wb30
MKiW9nm1nGcpdwF8w/3bJTkRv+msVXJan4vr1P9yLr7XMvWQ1w32S1471cR6zaBz7FUGz/wFtxvW
1m5v43mF4+f/SXgsgLh8ltu5/jum++a9KqhmQvV0OWjw4z5YMgAvrxbmzkG/WNFzotDKMMc2bwPr
52bIdRAetbWbBGmv5FvOh7R+SPt3tG1KUOPRF9Es9QqGImvbv4YErtNKnpcps8R50NulmQIU0ojF
LJQmVs9rkXCnzOHpZBMFVbJOjDu0h9MxKhxSSdF1dOxTFayAopM2gkL+l5KU+kzBYPsVVyQje0H4
hTo3Z0mWX1XDprNZydUfC17CZ6TPskQPrs1fuDJvmwpB19q8Rd90bQnBOMbUFq7sc9yBHi3UftfO
GGrf8vPIQG8M25YVzL2HbobKEGZdKGd2v2Flgoc+XjXracvXOFiGteTPvf8B7fYw/lLw+1xnqoCX
4EmSfooSqgz6Pe3YgcunOWNWct2Slp2+4jS5XqpW1ADBTSBOeTZPaiKCJaKOb+N6iqxywchco970
UKYlz5HApbUyGbhOSQjNDLLYIBi5M3fhEc+w5fvpRIKfyTa5/HB4lZiZXUekEWk/tYC0i3L1V0p+
NF+oC+udJswsIHmcF87MW/WpkJ3EJP8MlPrBDZlnJ0aEs7ib5BwQPxql5nbh2YEsICYcJ2CfsFqU
y0beTYAkkkHbPgF30dfax9DOYaOgNp6HGOnyG4OXRVUSDvaMbpryhyxuYNLHPa/8tQ7F6rEpFdLj
qC3usb33DEypL2BXuF/bSLR6uRS6ITMg4tbSO7ucS/+6vTueHB34CGMKIppAogAsnJmi+91RITMg
yxELcpGIbcDa9ixbQ5yzbEq7JB/SWmGXDAdWSNR0Wa+BZ5JaOK6M73qEnJaeQS65p+Kkd3ClB0rt
sXI0XXXDz8zPjt6TriTvp0eUUPRg6UQiIxTD6cBtjllf2eg8xHf2lTKC+0HHEZHtkizcSN78PKBX
4f8RV0iOZIcb40obKJvAuH98zzAn7J7LKArHy7rT4dVmUPE3FFvVcEO/GnhqBi5xGIGK87wvcIgB
evQzKZaiaeUjuTgNP3YVqAl94fqhFX6t0Kf4l5OtIu9CUaNu5T7TavsJ9tlrxrvy8ndkQhwSzsj/
VQL0TVuQZtyf981HHoKDEijkGhri067DxkqWPbT0+fkgYWIWfhRQ6MWGfcgrdXm3WudwN1Ik6+rg
cnBFCgc5haRhgFHAr9oyL77Dcfx+ETc5hHHJPB8S2/WEnNhr1ojgGE/mvu0rwZQ0TKqKDlvh0I2i
7vEKRS1Q2ceKv5pkiU4JDwS1T8UvRIYz5alY7McWrD17G5dz4t1VDz4yWssPDDWjXhFHKRSuA194
5JuBo3BingV65TRqcuJKgqzY48iUxgf096OIKd8EN+fD7buxx5SusLvEdhC1J4D5WAesK0yr7tsp
D7Kt4nV0fDbfCzD6g40RWzx3dZRzfmcAhcLh6Gki9kI3L37Xh6NlpNQboe3DvpAxuiSgLI6Gnycf
xeoahnjEcoJKdcf1Nb0qYTN4fnG9NNH72W4bLvbHqH3jVlSY2+iY3YsYNouGJqmymRlxR63rfWoB
+E1r+kDliuhSt56EdOjS1n7vXmwNpTXiPfT+ozHBSYHlYE5kxAsMD9V+STyvEbOl3fj2JrN1NU4y
ohFkZo8wsMakXfoasd/mXxeb6Ldb1Gy7o06Xlp9QBwrcbj4oYzt6Pl/DiYoDMwvwr/dYYVj5PhXI
3e00M1ibWt7JZElWdjm/XjYPz21kuAf9N56elgjGd0cevfWqdng4l5QdT0IhYFbfsjmLHRb7XNzL
5lnV7zSZY5+lMjL5yP09gYcHlr4rmtW4K7u6Dp+hKvrmA7rzy5KF1rEmcok2XPmZPnLk5v5rptUp
Bq4gw68Swv4ZbH7Tb8JStwoT6K4SeoVC0/H75m/uNBaTP5NaaMa3YJAZCih2pxR7St5RftDeBoYt
kC0OwHcPol5NtFHyITcp5MIox9A/HMDPJuVGy1Ew4Nmmy+Fgn3yUG63uao+lgNtoBWeAFkAQz5FY
qsap5dUiCcJunDbkaR3AQzBypQz99panJZteU71bRlZbHC2ZfTvWm5WTwzX2oJn/sJBPUXiJxv0I
ECxGqBVo2cvydhzcx7HyxIMolJ2S9FXtsNe5G+GaE7XmcIYPReVuGxJf5PFfiayAt7Ic5u3C7lch
+F1CoPH3BQHv3s8GGoDM6WNg1vXk4E/Vnn9OlNi4xqmST3Ksnt8hrosBQHvE4KL/V0opQkgFtqZM
uFXq6icQaVrFVaGnuWdR8JlSlYcRgLiAM3zv4twgvtB2X0m8o+CzHFTDcuyvZnYwQZptqnZXqBq+
tffiWAwCUNXuBd6P4G0qtKwrIAOXIdYBhPDsKFUgL6wY9bDESFiD8k4o4EoISIJkWpvYCga3hAn5
+LrLtpDxAom6j2/9oMVX6R/qXerkpv7Z1gl+wHHKLlbr6khSIJLElR/NoO9L9ph9Ig9OXtWmCP0c
XmB5loXUYf6uVBas8qu2yDN9KuNAVLIzGus7YfWiusWKKrTvgWlNzJom7xFCH+pqdq1GopHOtRWu
xUBDB5oegt2CLYmcb/2NxFuYKmz68lEFlws/WozmZ/kzZd4dkdvBn/x5fqzvfy4earSezyhI+g2S
+jzVhFL4KJQZLCptrbNyoXRqdH1Pl7u4Y0yaOzhpccEXxd39ObVLr1NypTTYnoYGdlUi39kNojpx
5q1MpTOiowlFjbblY41Rj4YUhwwoCWUdnVjT6raPBKjRrZysod0ayXGwL2IlAyCEz/LiIooeFht2
O54/kPZWWp/iDtQnQl3/DFx8u6QObnEeOTxnc9/JDy+EfvW19qrVOLRm58kc4wY8a8wHwZZo2Jbk
OTCVoe2fZRPmjF78mJkldNuLfVut+Rlp668GA70VEy7iLzWtZGzjNWHbqSjtXPhL8E96991ArVce
hhThuUJ+tPVz3yl7mkpzr3shx0ZDe2tY/joAFthPOgf8B/zAmlKV+3hw1ofC38qg68XxD3BANqPe
pvrkd4LmugLcpUuLHjpof8Td78UUJvG+62AgFrSaNTiuMxegT+EwtnoPzaMNJ87wHx8BOj0m/314
uApKc5jRAWOBCkcwPsCJ2yPQTUnRvdT+mYWzThKTe257G3P1IYgJ25nKZoq+RY0ghuGuSRv8II7v
cxAMkA7et5IHjXfm/zsqJ8VQmzhRcRGWd8R6/TFzHLQSlS5HTxUd8OovmkWt7mU67tZlfj885my7
0TIBgWnudkRc2MhwlN9+f7HV1EPJ9Dnhoyc62Z+ONPAGXMh8Aev9/OyftKxyk389mNM7u8V80Muf
Ec7Tr/H6Mf4XGUa80C+q4KPOz2g4PDi8jAuym9oMdVy7YhkJKWl8GMM6Z3Z/HFfzUG1GmaZq4sXz
QDQiEEohruSs8QjNIjbjjQoTfvRQqmwuFNiAuQ+qX7Db5/GRHZ7dr9jTYob00xWzqD9Gh+cmol4q
lCQDU4xwlT31MPt7sky+5EJ14Mqp7QgRYbc3h/5B6ISLO9MJgaBYZM6GBtDLc0xR107304PSzxo5
Aw6u3xp9gAulYllo7G8VsUPLjro1mgum6IsB5OBxN8wdO4My0/cTOQONyu2znBn7n3Ba9nDxpSvc
XULbc5sYFBd7ZwI+5yLBqsyfzerfLqycNx8c9HE6UpLJET3el5psHg+BFSnG9uQPKryQPtWAcDnR
QjHFy8/LguUJsk6vW2WBUL/nTje67irkMTpXpqkeNAOU0XPps9nda+mpbFFd9FNiB2AwK2EAfrfl
jcC/EhkhV2P1EMTD6v0cN20NUXgnM0oHzEs71f3Rg87DvY+lgkeYqVytrCH0gpNyA292gcmdwQou
paimeRtu1NOPmEqZKHtnmkwtutligVbr28ZqJrHeaJnyeJuWJyU9oQ38xIbaUA77nUsQ5fh20Hz0
B3i6+mYUwGc8uSrLr3MZ1BR0/D6izrQCgKJpeNdKo1N/bByRD1dwCqop6RqbDYvkuYK0mT/RR7Ml
XrjCnyQgmIimHWR98M6Hc7Q5Ssjk8f/Nr2SXgUKpgPyY9zZf+8cZRNW+ZGsvPAxuYzB2/x7QnfQf
Fyv8qS+S4nExM8K7fWxFcEwe3GfmsnYZhFH3A0L7NVHt1iezhJIPFl9a0X1ZW3cWoXjHqJDCA07x
n2wfYuRKeuUQ+pRWYqZCY27gLKHtbsN/B1oxnelOKNCVy0/BOkBkwXNdiUYmSgfYSG43lc8sVL+c
jcnoQUuQC8SOHQ6MCTP+HzjUfgQp1eIjB1fovx6KaNSsiNj6G88b1CW0/lIfYigsM0Af+sWCMpSe
0cL0IFKwXuovQxD7aR46A5WaWWVs0W4vydM2ifJIilNhxXjN4x4KbDQsF+ZukQHeQ+geX1/YIBp3
OYPKSeHHWNcWHDf4FE69rgRDsAEJreXj7dA+Ome/cRUJBX6xEAZdHPhd01yXuM65hFoPvct02H5A
PaKl2Qz/bbWLOhCC/LMe2M7v04Z7bdoY5uEb1ppKjk4khrRW1QR6axCYtnJ0OlG3fhc8YlyOfksz
N/SOugyQvA40ulJ0j8aJ5JLBrpE2m3CN2dCAjpsUrNRedXb9koWhGBBygnqOOPWCQhSzD8rHSLBC
I4BNvSb+jx1UTFxpGUBWIogf9IL8Q8aY+Q3QiHt4FT/51vvZgvtRDt1wy0Qgpjgy9x19DCkKGae1
+GlOZbLQKl+W/BwekTu39n0Sac+FQ+9KVbbtXA7rnrfNBn1PWsdqtO1cTZqeOxlF4kIH1fDUHLUI
c4XUPAPBJhnBrmcfBNMScbPFavQEc3g9b9WY8moSU57JeQKG7tQTodoQX7hm6TtCijoaj5vRwQS3
DjGcw5kaGoSd6G5nc7wQx/bZHPehvHua4iSVWeWCH8PNQaHuV9TmU+V6sU1eiU8vGGN6T65wcnwd
2k766OumECNHY89ePQqE62W1Un3jTUXGfZijAKuBkaTJLsxN+dPb+bvTHrrHMnJIImefz3C18mJ7
mDTb5GB5YUOZVIvj5gtGgF/AC578C6q9FpJV4n8/pZ/7MmlB9HEioqlVJuKXZ3fiJgYwq37OUxRo
1cihtw7yJHjb9CghcMtbH61vjVr7hY4LhVh4vjMpITsszRSc/Ela46d6L8vkBHcwbITfgTx5G9Zc
xkEHz32YUPf89XR50i5UkbdDQqqPVtJib2ksjhVnIKteNHj7c2KotZTm1SuZk1pwG0nFlkczGZnn
b/VwyP/UTYEzNkMNOGvzJM7245KaPKppq7MI8pSKsSSn63CQ1BCZwSKTsBXAFyI5qT6FbY4DP+2h
ZfUXkAypocQ8N+lokI5L8kfTZuCOyUzRWuf7sStcvVDM3lWvo67BYjED3mvktA228NRXi3M4iEQk
m9O1M4avr7kIa5QgU00y2SV4LzlXRcFWUXUgstzlBj9FoUdhkaAjp6s/QTTjIWmBO+seJKyh+DsH
kYcidOR52ZAuhSA7nwKMNss51mWhCsnFk6iyjkWXvLK8eeqRSV0eoVM4DvYTrNZTKguLavryvFzN
E+y9F3Xq9VHbF8k4k8aq1FZxPbymMsFRRXk7EnwsTQw84JCUNVvHGZumzhOv8WRp+nkNgXkkH+Wl
nsuAOgiqOZbGL7TGLYGEUJznzY7p+LtWSjmoHXAmbZRO2jPmF2qcE/7D+1ZrF8Y0MXUVs3+STLH0
aksZmEW4zC1GmfJN7tp37VTKQ+7TUPrqw01Zz0snvY6bNlkE5qKykLzQY29ldjfHhgr0dnTA5+Zy
2vgds5MlUl62RIyQex6P0UgrInNnyydJaSdknn4lpoEQnCRGcdSERHAk6tI1YHxo0MBNddxqtEGY
1i2NyxSA1v5NSq5h2QLJKFjXBdu7guh9yQrZfFTmQl7L8Jc88laf+8M231EUTzRHwSJBwGEXdupE
MfmYSHoNasAU896PUUdBlA/Qu7lbWJB0WJSxoLSC73sSisLsG5AxjD7k4P4PhwdZyR9BWCQM7AP4
9kRjVkNtABdCrRzyd0AQXNucenLBbbvo1l5ztX29zohmKOJ3M28z5yECvYQsBKXsfOQ0DFtb0KHL
MWRQsRF0wwozEdUmOC9kxKdx0qhClMvabD+T5viBvL71NviRdWhyqUo4ugVQDW/YR6PaRHuMT8JY
IRpFnTulmCuIDznIh7PWWn71EEZYS/R06SPVvQKzUhrtRtPbkNWONXyUuVY6Es80Kd7RWP+ubmAb
T5ZzSbZW77l1DXHBWXWqgqlyQdRonffbFfiuFZjWxO7to79Io7c7wL6cbs/Egeuhkag7JAmopH7z
AGtCKaILRVJ4/BKsYBMQ9TqhUNee2S3VAfg2fVeWJaJ3dYfZrJw+W85BaWKfbCjM2EJqVHpJuxLd
D9XjZD1z9I+mwpfIsrg8UXA03c1+SZLioNMWGjBmqTLn/WytVeqL/9nBtm+cw8n8lHWGYeVF4/9k
xN/Fzav/VYKXQzIIyVDGjJBmJuG7M/kwvDji+BYKnJRqc+u4SCxS/fOu9NuvO6HHKvqIdVkiFZbn
oAiKJO2lPO7NUj6QYFQcCh5Y31SorbESycHH1cmqomCTS8teALHP3x8U3wIw7hxbdOfFftS6Swjr
puyJfE07KGRwmWzShBEAccWcQjyqvJzGVdpcJLvPBvOEe2fr56cqdMGvNK1qoIJFs+NHDduv+jGb
fBwV/gHzY7ShTJeCWPAlLH9NfAVOlMvvTUSWkypYDwabDw2DUjyMqUOPVtKBRr3I3omDmIZdUYDz
qMwmqjkNBjjFnTAacmJmYzOUmo8vikpow8LrS37qCP+j3qxQlcznR+a3q4rcznN4M4zVPj5nm9em
7quOVeggCo2uktCPc6tSw2lwpCsGChKmR/Nf6GURmB6LqpzrCGHBGYRzB7QDfhwXODDhg292GMTa
4Lr70YYU2AzXPGkZGD5yNfhrPntHBmZ58uj6gqnTRg0OhDW3JLDVTxB7RaSzjOXY8dcc+qQYCPIe
WNVFOxMkSRJopWbIe6qVwBgZwXFWo9pFCbWeY1r8SvpPU/iHdKUbacFCw9QmFh/EFQg40ACAkfGi
UFQgNKHUjlzh9Mm3qIgoEm4s4MvekWQ0mxAlvCGZBhj80bSbqaCaGuabfJFnHsZlUU7XCSCRTN9D
zJb0KtZvyNN3dLCH7hQXKyO9n8l3xBX4rjcWe6dsnE9ijiuCVhTgIGjH/qNWYuokhS7h6J+9jqh0
X2SyQp8gEpzTqaYI1nGS/o9Kek/oDGb0fIetHqJwr1A1Tjkd1H1oyUVT634BMlHSVL07IgRGYFsV
BtVpeaUqqcAuGu8YKUFbCexq1SgVfGGpRZaDSYu1OZUnUX56MEkT84BVZhJY1qsdWi67Lj/EaPKB
DCPgBzBwbTIWO1jH9N51LTirfW7pquELpaC+NaMj0xc0/fCoGxcB4QvLVGkT++eBPV5QAD3vwcd3
c7QP9uthcErcD2HKubLpbsgFcNT3r3wd7pbyO9v/uTTThVX2d6cB/8vbG5eGkse8qFX0BniZF9/J
TkLm4WoVK55ixxroO7/UBwsaTW0yXab9DuFvM42DX85Rndh87ip1Xa502+9CCAs0umBvGCcNeTV7
2s3mwDyDl2z/M75fZp5dYHHTh5puzjoi+HCXuVmwgfo4wxYL7sW2CRIUAqZtGbrGhuVKljmNK22G
tHovfLkhBaYVpy+hnDwgJ+/R60U/PLBD79+G7qgd6iKK+Jx5sw8PNNz+oSnBQN2QMH67N54Bqrxw
UcQJF7oTMKD+NqHuHEm4zRjgAA1lXxuzIbVkaNdB97M+Vc41htWLKRddaae2H0uwhRWm1Ykg67je
bdWIXDTJfNh5u/ZlmQ+T5GskX4+uLAbyqHHjGLSOPktFIu0zIFvqgZBvMpg043d3lgJfiUH5wD+C
J8SAV0w1oxFwxJhccXIFatzB0uAZSha4qRunkB64PCEu2PZEpCH41IMNrHXQSRP4mR/QC8ugM5im
SFiUzR8xvCR5HLSdUnLv8WxqGXQugSpjrfD+jtbhtcPrBt8//d82UO/LPjRt9+PyP+MZBlSmFq/X
7G13j7q9NmyJo0fcC0kcXAAlwA8ltBxjwadm1zyVq6jxiCyi794FaLsQSeHFcNrZpQ/fx1+7L4mZ
zZIsOkUyTaAOAMkexZJ3g6ODkyDjKSt1TwFO+lGtpoE4XRUXEDXL6mnSmdnNdpMnRIcsa1U6qGf+
xbhbyrMLyO/NjFod51mugPNW8bXLWwyhePL0TEGdFZe6EhNEMBUsDdlSrD4rhdC1dlgQ+eVuPGBs
ApOcS4zcaVHfE5csMjYKrxYFXPKwSUz3H1LLIUwZQWQ9oW0GfskwtwSHXZSQBS+/CfhaL06jQ+aC
tE+mC+iS/Dumn7H3kTZiYGz1SHopVwSBzJXHLH01E46Eci0QwbDRUMaod9XVVriZik4QfjmHzUsd
BPM6Y5JynvzoLIUV11ktcCB+ucm1Hj3DZICi0fNjE/fQNgxOjTvLiuvYiDxtU3vqOU7AAeMWL++X
ywllBHtxxQ4sDtZYfIIRYD1oMmBIJuPCZv29flvwV42XcbcqWepLcHZtoYKgKVmA3hSsF3wjRRKv
FVAkLj5OYHpFpi4zbp7ErR0cRRyqvcxCzUWS+VIzpbXaK8MixkSjElLtafAJEbo0ykk1J/ZXbJvy
tz6Z2rqswHNAKNJiTCZcO/0iJZGeXP47YeClPHFGf5M1QBb2JCt8RVJQ7jIXr0EVgrL4ksn99MgE
EK3KOWaXtesOq6JzcQutSbBGuMAnme3G8y3yXtm0qY1tnVUhqjDx82Xkrwpzk+eEB7qXfuWOEFBl
9QpPzlUsy/RrZxo8xuihQJDxLgVS/aSNrpaCASZOYgkuThelAvMmkSYmrl8W+vkU83tVOtYbtY+T
b1SDZR55eEYK1c0Kwba+ups9kQxCLErCDCbW8qYNCPA+sWP0jSJJlxyKXX5DrhUDQ8jtWjn4f7Rf
Sz0unPyMsI83XWYrP0NhwkiLAMvgn79OrtI5Rz3lq23y+bw0wl3YUO+n0m5yURReeg3F0PbS48/b
AIlAVtUWatW+b6+wqv/VeoFHQgF/RbhmQuAKIjg9dwsE7sTvISD9VTugVID8RFd5GoipQj9r28MQ
IWkKvNTS4gMRFXJ4vlWsSHbzA1meFAElUUnq8oJZuCyMmnxVMIGLvdkDYRiAdy65QKQdNFiaMmyv
CKLe30yORldMRSTbH6uRVf7pI6v5cMDFaSwOo1kWu3Nhx3lEVkW3X7psMPJyoObdD0xqdwZJf2oS
gF8Xl2Gre3yNGv3R95CBjdIu7pFLb1Pm4z57xmcJqfavYHB6ov/TX3rvTaGs5o3jOLPQ7mg1HDV3
iqGpjEgRa7Cl9RSPsfXYcKoL7PIyBEDl8ddHYmFnBeBqeFkyc4TiVnTSxEPuADYdO1wELXCY1+P1
J5RatwlTfWToKSOsp5YGbaV1nIaCBElHwe2Zat/Qb7HcHn7mfpccb7nzBCAEiwoaTNlVhTExVJXT
RHT5Hx/2Gww8jv10fQjl5F5avh2qdrgbh1ry9+ugYJQQUf7cAgPdLJgp23EKMjn7IIizHeUDk2kh
4Ath/PBGKC2yoQonhP7UEDDkSAf5SHpobavxqtKBsLMvQBiqEHNgZF9VWP00ZewGVc1ruxNT6bBD
9vHq1TnBQeUHVMbQkD5Zz4aU/zXemtV4bKkgQXcQZfWtPOUTO2SH3+cbc+ySaqf+5ndSm6asYXKc
XVTrmJpOUjItKHIzrI3/9JsPjSDurK4aaXeXfbS9dhpLi54TAm48n1mVkEUlgHf8zw2Tl0eJy8jq
CEtdVXkk34TVc1Er3lcQjAxe7P/S++5Tb6AV6vMKY5Vw336qzzOHF9heaXuyQbIPzIkumMsJsq/z
cm8DOTRKeL/GtS6THsxLhEBmRVIR10uIUOdcAMwIRSVyh0MV8x98xP1C7IW8KRMA8fin9OWwPaF6
+XBZMDfivZK75UdSEB/qAAAkAMR8bW3TmcZop8us6hgQD2RmcsBXdy47iebfuo6n1DuKIdQcEELT
XRIMrgFTCvuD8gQXD+jQrX12YEnJwpMrtdqC0Rv7Figv2L/f/PTXO48COuTMtpRyahl93LY0R5/A
vaKqwvzpH8nmFRGQvdXZSjcMeyQO6736Xw0TZEdK8MOqF8YZH+wT+FEzL3W8gjPZEjps8YPb7U2Z
SbYJvWYUg5Y5lo+R3xd7gu6Ou0erfskMctYDOIu44HRqyICYeZnWzI/qgXX/r5cUr0yLpAMcSp2A
O4mAurMWIaLOHPQozb055vt2Y7aS5i0G6jOU8xgDpkzUmiMUuXAzTJEfeUoi1gExQ7YIgu9op65v
yv+gtdRERs9HncPMcmCkKP1uUUdgNLqZvLPkF1tODZhCTjHoOn+fHQd4gCL435Ia0cqQoyQkSObU
+u9iY744o1Z1ztgOyHpFFl4wNqjFIr87kt9QCmmKdqx2ubH48g2eNJmBsup9qMvlFMfPiqwQucSC
mQoldIrCo1J5rZRGxiH7sXYlhEb0P+v+1Bw4D12DKjQEwHwq3MZj7Zabuz/fZnK1uMH7PiLag1UY
fhBZteFQb+c/pj5b0d2aQe2Hx49gYn/LvrFdB5iYaFyEa2L2N9nLKyG8PxkwskIoxGvXRaVg8Yi6
hdO5l0Wccg7mjFDU4Qgu1VFGAR9OweadFKSzwUy/Mc8BhSHELC1MxRf5xa5cw2D6jB/EMCMiNHtt
jcPwSUAGVTgRiVO6zn6QkijTm+PJFKCxEPOCFivN2Y9AVFFTiX/0jxSkGOdPl3g0xVLfWd6Xa6o9
o3/iiCWZApaa31AYZXmggIgHzYRYakuxt65ocnwRIaevDIW9W4xVV3MSYYkJ8175pmuA3AdhB1oT
CuCaQWUVvqLbCZDsRuIEdR6Q7U1Gz3XxRdrf4o+GTdetQ+LeZHN/ZcnDFtG25WD9Qk3J3DpcCbRF
RN1M4hVD+fsPA/X62KYcGtAVU5nremXurvH0F2aMxQHPTDlEG2FJJbTcsWdb0dgYEO0X/ATP2fZn
KnV619xyEaxRxdXhvju6qyKFUEQ/xVg7QKe75/DC9DVtmg847npNSCJinS0wr0InQsX1fIqnoMZG
6Np3ox/3PUh3ki53akxc7Y3jZ7ByWqeL/z5XbTykIOrwljj1+++oSTZtwMxnrMRA0mDS85dlQ3J+
W4TEJzjB3ttEJhDXyhkTWdI6zGyLYK5Iv7YmjhAXxEu1nYZimJZyExy95GqB/3iy32RWOhDGYJDp
OCMpfdknrdq7LfFH5pw1qV+0An6E+hsSKHl/UWTZKesYkVNEfrmAUFPDuxzwY8zqh5ogHp4Nrtx2
hmuw1sfICbMjF2wWScUDwU8QOq/y6FOn9C4j5TY0N51gNlxPQ8yqbLr3LOb/WHzyQ1eW7XKQcmeU
0iBwmzte6sFawJ57UZhqFcRtJJGcdj5sOyQrYVSOg2lgyl1QU1hSr/9RSR4cayYxWXyHEJj4zQaM
KPmaxwSR2uEE9LFoeWXl9+lWn9IX9qUBBbtNh7sacp0XOGnEBzG58h50SF9WtqUMBqOxkKU6d4wE
I7cZ8aPdHY/eG+LDzLKsTxG5XM2W9TQw9ctKzgfZN7tJNnI56tVOsQaQnW4iU7VtXojDgBbZe53V
QBhx/RRWdzwjoaClag4EqxnmZuzHfS1oEZD/kNt8hwleeALbiyBVGHpVis2WPbcILBy2B12moGXd
zFJ9HzNGhWEbfbXD2K23pEWxzmWAMx0QBL/Z57cOEqp5yoHw97oDJmXUrOjqFCzHLcA3hpntUHZz
4bha38uahNTre1BvAyQ3+VwDRvlTMiXVYmA6ybEcTFIvkSGyofrjWYEtU1SwcVW5oJ4SjW4PIrPv
6YcvpGK2nrG2KvLJYf701zOtwiytY7I26hAh51dMzBzgFIAPIf0nCBcpulv/NIpP6Lm6I4bRqNV6
fzeBCSuEWmEgwgVmOFXHY+GDCIaDfYL9UBbxinLVv20Zb6W+yHSiwTZ3oze1XlNA141xkJJek95f
IC6hfU7HdaifWkecT31DXhMJFODeK6t7dCyOEQqZ+oJMdIDaQjJDoBbuYG3NGXDuZ85x4RfRTrtY
8zuzxUYG8yVNgMVgotIeOMlYyoDOUpu6405xRrNIkYolesCESG8XvhgD21YjYkRvbeZUL2ZDzwVP
bI3wY38ZOAY2F+J1LhmlkhteptmtsplkQi58nAmwhaF92gr0ZSi2u2FYF2zpKxIZGwMMbnzLqTfz
VBQHBcQPgZO3VZZZkv+HWXhnHZqWbXIcNSsykh0w8U44nMi+r4WZYTwChpVl++x6v+MDoaHSCvpo
nN9BxI758tTFHWDkq3YrWaWewN9k5K2OIvpGL9GD5vN5zjAKoSqIzZzZKOtNPzeoVlqXlU5J8QE7
xhCcV7F15ri8wsrtGCsUCGCiT0etQepOYENzQXmp1kbsnv3tsAsO0KyWW8YypajDRf4s0+aattOh
k2z/xgeG0AfA6n1c3OS4Ju26hyNLP7OzBjJQpJ4TTB5Z8QzHBLo+rL2y4rAOGxFOzCgWu8gSXpNQ
TC4uYT8pTUH/fxSu7DDFuRyHxufNm/ZvSPWfyEi+zoujFjAB5BxshQXXtOV1H4kvC5hnOLVDat6j
/gj/iBhhal5R+dg2oc9+CbxJMIynCAKc6na/vfVjMwiTGgAG0AMM10N2jCnYOa3K0jGugEDzcpdn
7E4tsiTklYzQhy/lfCm+iMaBe6ftnFEtPeCmk0HEo036tY3cu7v+w60hXRe+VITPwkgSuR0XNtMw
PYHQpkK805WZy3ALTWrvtWkvy97JoXLVuQFiWnqjDUXQi5EU37szGPFeXoUlHECl+BYlYvoyMBxP
jCf2xUh//3xj8zVIqsAPi7V0X421AixDL7IYxc3TBnrxDJ/71edhrEP3O621BmoDgX3e+vFQN7kC
LykwLrrpR3JvUeHydHM1Da4qPji3/8IoWj15l5DUd1trCBu9f7B2TNDhFOhi6UoByP4VtmlzWoLR
JjUnm3ZAEnSyMRTMQzx1snTZAXs9LkNeJXiGjXWyQ6008u9tbPMCf5OBQ8lT2eGZTFz090KzgzG6
oP8U9ChDK/3Cd9Jm0ByHpx8TItSGnAjgYrMje/20v3O+AOB9DG/q/joZtN8P7vTcP5iezlGwJUa6
eSn//YV1QkytCrSTfx1eWStJZC5yipTdeR2ubrgaGUTdo4LiI5KpX0IQrzc8ZAHjUOvxYqKAip9A
guXPKDZ1ZUtJsU2QLlKBwDm3yc6SBwQYGUD9Ee6pDH5bPR/U9PObfl4jPm271iApCgfR0Z/0M5Li
E2hBNjUIovveJStSicEcr247LI3doPt4DcjVPI/8h1Bnqke2C7s9JF6BziqtRFVwjLLGh/jhkI5y
lVJQ0uRLjPSpOj0UbRryTOMrG6k076J4FXwHc459Mt+poTAcfjR7Nr2bY0X1oCqUb96cfGTvf5O7
T1H0mjZRqWQulo8Jep6iiTLTA7Vy9AeJ1lnQJdziBlekoP5FXUk3bFGbc6gLxvzm/IXc60OZUx1K
0FtFGrS5/4zQpJBzDNQnASP97RWGRgOo+gcySElFi97yMXJL5ReD0FSsS0lyA9a6t5Vf1hIbB1bI
py2mAvPQPxjprN7cbLyV//2HXKS2pydXceaDfPfAj7I+4lcsoBSWcvTjiaX44DBIfaYkbcJjWzWD
i9oBKeHoA3m5+jIzjZol8Oim3Savo/O2YrWbMY4HW7fNaRq6aoF87PUGSC9HIdkms4P6hoaQ+QrS
4x3TYXMfjVE5OND8QKhsas0WrPID970PabAESv4lJ2ALRDwYHfZ92KLX6MwGm6To+c7GqF1QLbOt
sLG1f1GBzhRcrh+yMmFZGCo0xlRP6eJwTJnu1x+vPCoKxylwaAh9W4scF2IuRomrBDk2Xv3ub8DG
HOgyzCKKM6tGqWyf5R+/IHEzVu8L96LW4PFMEomYANstSd7aGOwJ6e7JCGZQTCJLLcUJZUZP8weE
o17hCSpH+zZrhcighHIb2ZYHo8e8fNPbWWl7xJtoLktCKntyZNSJ68EvrzaUR2T29N6i8DHOvz4f
8U2tTEhdC9sLE86aGLXB9z+D0os/TM4AowIC6h/Fvpo3khTsGQR1Hrn13D6rM4IQTmrXl4SZpZSf
Dt0OpnyHMxOfd15kkC4WQQV8Jawtf+onk3/0Xf6iV5aLsvgTaQMJFNm/G2ZIeuAB9KLCsvkszmcc
WoL/7UDHKTmpHfLroT2mb7MagxBRZDCz9d67g3H8VmV9cCMqc8Lrh0eRQDXQqfECQzEuwryT101d
ZR7jrzNse7ymInkRNylMd4s8GyTPLMmYX9LPOAdLhjnRuyQIMHc9/GzFLNucjh0sGJ5T/hlYtz6S
y62DDBzVGAcIIaDnGBs42rtTDJxh9TsE0ShyIxpqOS6raZuxsaJlDimSvc0Dm6i67/UTNqo2L85S
58Czi70adG3UVqMTGAu/sgaFeeocVYGq1jZmGH8gaoGTN+47gbBnNvn2u/Ec9emuYWmK2pynQhtc
xSttN1ttJoOslxNfRbwAHrKwV5zxgX4CRw1JKRPigcoxreTtv/rVsA8av76Xg9Q2fjQqycludm6v
7kkyLzQOSArdwJ4SwvZ4OF4ucy4eTXQLadpsDjDZNumF4uhu7HsvXMLZDE1D/IKOvyn6DBOvxfm+
25kKu4HfYgzZA+2P1Rd9DcIeq9aNKJFQGwVzCzfpQlKlwUlbyh69ugTZE6n3lUBlamP7lqy30odx
hjmAmRztfaoghDlYmWV/I/gfCsmlgAD1DlWhHwMXchi+uliQVsrreJeLpYqLyATp1BhZas4WUM3H
wOeVGGs8hFtS2Q8lMxwA0Olo55gf3KIclgME5sOFVMUmIDqEy3w6S34KO4iZnbcCRXxZRtyjzTsV
ZEj6NXw5IquO0La417gbvlocN7ur9fRQod2oHU+6oy5YDqr8R/IeTjayAoJisRI+Ox9VbsqnB/1q
nLsH7VztsNs5Hxx1mOnk8foC8/vTA3YOtaEWnDF6FbeZjg+6+18EIFuk4dGrxIK9WztlWYhpDNKR
fVj8VaMUhXDJE/ZMPzETx70khHpRTWdsrxbSwqzPlvfbkbqt02ZC7aRwnTfWiwV0hhZkT8h19WeA
e6dviYxUESTsULOVcIKOIJbinrzT06ZMxzZaa8FDRLdsep1FV0VrE372FiGFX0AjDz7PGL1RWUGq
cm1oLvVNwSxihHToJQTPbWtZ6Qn67ZX4GfxBp4mlTrU23gAvfYwufc4YFKHv8QJSzwjHBLNspHkU
f9LFlEqIKRo6oXB2J05Bw5TDSr2VCnuzDTu7zwSeKdo1EJrnxtrilX2IJtQ7RYqQ/HaoWuUocMJL
HFIISWtzLAldb6c8VxOBJN7pITOuxeLkLX69i823nFVX+87ngMDDyCoYWV1UGic0i7zgnu/cGh3P
2lWowyF4wR/Dt6OXPHHbih7PhUJ/mOqM8+mMwMWWFOfwCiVwhHWu7NLVdkr9jmJXdLS0FQe3s7D6
++WRIPivG3m1hRwMbTig1rQCMXSee/IZ4B881CygGqxUcvJJi5URemscaUffNzpobRMxokb5OZgL
PzC10MLfvAqirumk1NrWRoFu9Y8RBPNaxtCH/eP4w6fXBcxctdncYyUFe+PYEwarUvKQzq8VRyHv
z/FkOHaDmv62vLGnsaDVEqZwrG0ghShq5V2BVC7aDSb85dDDxfw+TdVZEFICR9WQ7QJ47CapmeoF
4iB9MKjrhS5Le51J++8By7NtdWq88GpGOX3aJB5zfZ3vYj14vFK9yAOaKDKH5Jc0o72PM3Op/PTB
EUqCdBM8vD8klFq05Exh3NaGliHXTXnvQBVYyCizkLy7ydUJ2dlQzLLf4upNWtBwaEz5JMMvRuDo
Px5LPNrKXSoGpTYnqXzE9/0UqBUc0tAB+EBxd5rRW2h9J81CILC9cDTilCAYEX65vKtZHJad6iol
AG6gboBQ5X30sq/fOxEv0jZbvpCqHBgcji+95G0xzJrAe2i1U/xak/B75+g9/kWFVeOolPc3ZpEk
nDbIVXWFmLBnHrTfVQj73u8jcjUMyLMtloPe6KYeUd5Uh9RHb+X3NZUwvyJf+aIYLYrMxMDAL5Z6
sdLqNyE4HJqWJsm6qOl1lwfO5RsONXsc/TsEFUrxd951oi1fa88ihqKsCR64prIVra7n+L8T7tOl
1hwTmUVTGncrl9GnwH84pZgKe+blTUXaH/4vnHVJwK+2lEYxC1JLJZELI/TubZT2Fh4Vl9y1iwW9
qAFC0RUrGae0Sb4BdqJyntzCJB0Qb9x5b/lYe7PZeY0NKT68t4T5vPr6fcssH1BoS/oHtbfjQq7l
+i97z1u3MoFXuny9ilfJJGUgeJu+AMs8xhnHb+hyCiS1aTSPp7uSaRUUw3HH/iEPVj43FrkUPZXe
PZDH3Z1wCy6RXUETd49TzfAd1HvgT2m0J6uNwfC6xdkz4xCmLawHj4RDwuqYMTAvZ/rIxjvgrRnQ
UrBq09nD0DcB1A6/DAy3f8H5Pw/BZd4Sxmugj7Ar+LsEC0SnS0wwn+lxv4hWimA3IABdfYv+x2ID
98icTXpRwczmaoZ4Tv4WOTg8Q90CKLUJJey/urYmDQfPNpNGPYcvRtvFKD1g2Qb5mN2Jpt4ZEDo9
jP7KRL77xQzU7UuOtyWWatLW9WW7kYMFmsciTIgfLgPAnLdqRUGycLYAw6I4Cd82wThmqKcsyFGJ
W3unIc48jz1pYcSrnFhpaj7MzEcrY1miWamIyf7jxosJtS79nT7PKTztxCgwA8pkdrKoBCd3bgEi
TYVBZn/zv8FpgtkaKg4uafQ2hOqxvVPg48YGoC2ZgEAsOV8A5JroYY0Sr67owGo8VGMq3mOL2REM
bJJxYq2MAIX+vE9k6Awviuky/DyDi7SHJLXDHGVUmonKV9D0ygBoCTSOwteHhRaXrKwSNTJF9bxD
zTWvuBCSzWP7qojWJzvS3WvNKTxKCnRbLZqeg842nH35aI4BMfs83d1AxFaXajwFlVzb1hFFMaZk
R/iYfFxGhWNMvUTbIZDXsjc0CXftgCcE20M9ynJ2HyTfgwsurCfW+2yXsMfpdSCN46iqp0gb2Glp
py1PItL3cVlazdlNhPWe5TKYZ6U5IxrDvDWdjGi6m89qFLGmo/T5sytNti0GV69zkhQrxQJYdmJK
72XaEH5sv7D8PYIoUkohZf76m7AjsJycLo3fcGpIpYvbwGdzbW00WYfYEIMaY4Av3GH9Kh9dkrd2
fpildrurDDnOHGnVST9pmLme0qO3oDwKYSN65wBQkCTSpssrZIOYXq7uXTrTP6ZWPLYPPWq7Ej9K
zRv6jBKimomXa3q5xtIpMXuA1QXDYOT/UPcx7c1SATu3OCVyecmHs4gB07YAuyQT+GmAlKoueZ7/
4Jmct4OiZ+9PMOAzy/b8NJX+wri2+AB/fzQfk6MyJSUzkAjt8N2Slbr8e8E6ymqJXjihDM1WsCd2
ZQMn3+L6F8jWppdxfdhw490uU48pJ0S4oyTcjGvmJmkiSwlKUYNoB35abo1PkgpJRe9BLEdIQGEr
+TnCgUmrzBKeUwYXPCcLntYLkElG7iYwcnkzbw9PUnTz7UPQPqDdzl6MaG8K1Uu7qZY9adc12SRv
1w5nCZpsEaGpRDvLZSVmGqJRmi+2d67CuFc2b8Zl8sEqv/EjSufYjEuZz9fknpFOW3PdrMGvQC8l
np2L1WJeMHirpuEgQyTVEpLHHm84J1EP2rI+QxFtS5+kR2lxXUsC0Q733IQgSggHV764IGKo5kVD
dhmZNtPJV7IJBmq39WLxvVwREytrYwymvAUaoWJ4O9UVXM06DKxfpUnBSOCtWnq2NPKH4mdd4FZA
3yB99GByrrXCjdejsV4zH7p4AzGuLwtn93ZbJF1D8pRzA1l7bWaURhE+JHU59ht3nBeCezEp4zLy
KHu4SqFDx1rJvdmG2kW9tVkX2awOfgVOMYl9BpRTAKngyR2XCU28yIS1jEuRQrlNLpFfBERFDEHn
OY3pYwnx12AUZC48YdJ2v+xK7QoDKrR8l0SMJS3PUqGrKe64O59SfqUhO7m9H4+G2bDruOZdvZzY
Y4j/kBazRRGoMb3Zl3Nd1XdvkALuQ8imND2hU8+VilyvALviZ6BT7pPiQk+vX8uerwcRXJkjGnyS
MqL2Es+993iY1QLJ46coKOSQBWvo7ppW1nCUnGvWom8AVQnkY4KQx3z54xBSmYIi44v0PN0P9UO6
FCF2OwYepl0COBQZDt6Bku31GqV3gNT33Z9PJehpYDIIsfgHqsZsGYbmd0hu5Nhp4zBveFmNqQmJ
bgLaZCCtMnDW/qV0mAGKzI0xw0H8FNvXD8zPOxvdsoW0mogUvW1OrgPu8lxJ3JYYU4xFvVfxf4nk
ZtYcoW0s3D3B23q1EYhNdkRbuac6zexfA0md5RO4OUed5doP8p3mVS7uPzyAygkonOBDRjpgI/UZ
yfyRKdoqMhIsqj9OEuWZT+1z19K3F0H4nJodwWoQ/mq0wVD5wA1rSqOKhCc61WTaJuQq+pSgF24q
NaJ1tzBS7XoR72qQ5Fh6mDA+Kh4WsaV+eEZt5OrqLh82NZVUQdL/4v1AwYyxMWKgYpT3TQrrsS1j
JErnY7vrstb9X02w43c5OHwOoffuZdRLOfoOvWABYadUB+5eXNUez2gun95w/5rRfU+N6MK1VcSR
l6r5TxmBt+N4OBLBqMlKDHhN/3ZMpM777LdE3dtQEFmuTwohv028sAUbaAap3IFeHvPVTBHqsD+9
yUXjH8UBg4SdNnTO1V9pweqEKLgdRu1qZswDnWmcLUDxcOuO0BMtmuFsWIX08MJREisFZtVWKdT5
bpxJGXfV67fkywfrk2Mz9Kypf9Jb6T+h4uWi01HTaE1K884ZhzoeO+a71sTp0ardFbeHjHMvpS6B
2zng2kjsmfBtpHb8XW2RQ9lUZzGqNqdknU/19c1v5yV1/JUgKjL8oge7Z8vxYI3UkMAhp1KQVf6f
AT8B8SNQcFkwKjTLm5ZN22T2Y4kHFuAAj7A99n9uPLYlkcf8EKkIPAPLWHZD4q9Ex4VgTc4RnQUs
6r9lkfV55plP3CeuBVr6oA/FXgd2zK52425Yz6gU/pfpiukxSCBFNxgh2jGN6kIYPxbcgkNcaBKL
rJI5kYfw2QF3fZXoYShGzuiCOE1s8at13I+LlsJvp5lRjNx3CNNiG5dCnA/mGqxu8hi6eDoEtIl2
/b4KIpOAq87woBXpNyhnLL7Wxsk542q4++Cbo1JA1fwvQnvhgDu8M8UUgVHfeiOzc7TURvYLpj7b
/JShGCp09VJ9nX1QgCudPlG1Y3KD7JTxTrFr1mz/e0IAiIam3dCuYHyY+Ww3MW6G7byKkeWI9dD5
oj3wTSNSjfPITwNK3rUU3fE3HRx00jgFwNZMl0A7qO7ReObV873vxVkdj4u12MCbEVNqSzBx70tv
5Ankl+XIE9UzjcJLs0yn5FXc69GN4wRuJnKJT9h7MUWd/0oidylf9IqLI0Ked3kzYLeQhLL1kQuz
zQEGFFug7jqJdVIt+qtsTWd14QNNyyK0lRE4y2qWJA6bX6hQxjjdwiMgQiWX51cWu6BQQKXvlV2e
d7OElZ4wHqbDuWZm3exCOrJBZN5W2/wufmKyf23d+lM9oXQKAl/06BX+o7zByCrM11eSmlxonLLv
bwnryUcpN8u18Iaw1m/9KSUnn91fYb4Ic+00Uf3chzRchE9XEFg8g2YyXmE4n3PqvdaZ70Bmlx4q
hY45hIZLSNXTLTDnFJlvLzHa8TnMs/tz9dTKeWYsOtQw6LMfCKsFoN3vY2w1V2J7WuxPB7/jrvlp
AAOW/giu/q4O3dHQC2muu3B1os/n/M1TxDy+wdnxyzur2Jkz/XPzh9f4JIVdPxOfTVIV8qzlVNuf
5SaT6pDUZkIfEU2r1dMecHv4gKEXkw7Y7pZNBr5Bs5VPB2jDh7U9o/CKYVM4JHfnzRsxlpXt2Jxk
J1mB91DG7/JuFCFZ0pT3xd20D0tqEcOpRAlAGH3luE6yyqwHHvlzd+toIEpfR1lY4qyvIYtaZyjo
t/je8Fhhhh6eDX7VOl6Azcu9bezVHoeQU9CrJsosbkHtdZdliMgozvMNra1pEqQBXJgX7CultZjl
OiJtvTLu3N7tUDFO4K8+NMVwcPl4JYud2cZaZJOIEWUbE7OnmpwuKZNq2fRUnik82Y1wbBNv9TqL
5S5l0YtMMY1BNwe+h0Y3OAk5Q9Yi1KQbX2wxP7lYjJH2QjHzFwUt3YUEhL+T+zZt/OmAt6KGnyR+
+WwybazjpgZM6lN6bTHsp68V13UtTlgPVGMmettbd88oGsqT5uR8VKxqpRnqXv37yWwUnzzYEKWJ
fC2lK5s78jP8aqNY4dA/UKvEm6F/Tsu//ZKznI2x3W+/RfX/vpu7NbD7YS/dAadilJ4Yi3r2H7EY
UcZht5y0ff3Di59W58d92q+kMrAw+/8b2EjiIbqM4pqWHFc+Hc55gW3xTZg4yzEyHlYxTJ0xNHgK
eFNadKrYZpHFmJytp9+HZ8wAn+uRuG8mM7AblY2XPDz72X9GQi8PY3nMfGZZAKFyESXU9PszRhbs
/AUgq94iJQjopnrIHpf8XI10eYf16dpacAghmt7Wh8yDeg5Ase1A9P+jQCORweUqKY4V41az0fpy
pcbUUO+l6fSNIZsfQomJSKlFNfqUzyw0+EjN6SGVwNSaRHpxqoHES0LxKdWxVa/MqYDG3f6/HwRG
5qPPkZNYMXsIbCdLY27jgb9gz8vf9S1WIv5eaIlAvWh1Orp6IBUGAj05Fka50KC7F0jG1eNoywD4
WjlP8sdSKxks+xWxlLQ2ifXLAsinH+Yw+B8WHUFjOV+CfdAikLkcYQfNBhcfn0nFD81/5CrtIIHi
S/YT7T1v5mtdbqXQisCXw52E5YQzqeVYORWxdFCaSkF0ynwHazQS1m8lL7Pqdq6nPmZjDXInf1zE
MRr9s8Od8diq6IRTbCgEQEMXTV9iR0a0/nSX7mvn02taUXkAoAr9iq308Ivz6fwesv9XBO88QH2+
R+ra/6GW8qm4vICkBJf+cnpw8XzJRMf7w5k1L73gdIbugLwLHtPvAaYgRvXkR16wg1OKKDhzFYr5
6y1D4t1JDsXFEf6DTveK3XN7eweIBcTNo6jHk/U4+7rb/IPX5gOVFM2kchdyezttDM0ORGOyJlAl
B9qumyWQJWHbh8tza28bQAFbR8wl2FhenYni8cAdmaU+l12HSb/aEJzUkIqO166ZcAZHr4Mvjq4s
s5m5od6Wa/U0ZxzH8XFmCWJSLq3IyIJRV70ApkCYrBfh6vpuG1Jp3xeJpq6HrZaaaTOycCRwqoNh
fZcTBqDyImuqEFVaE50M/u4b9DGK7x4nurUhGBc9LMAMYhqUwlx1lr4yoPsIlXpLOdyEyvXGi0Ro
MXQGGwm5zmnHo60s4fQWbC16lVpH/n87Gg+mrMVZ4XnUcZkrEMAG7hvAG+jcY7AfxWmhoM+CfPF6
Tv5Bddaxuri+mRPBjbz1L9Soea0SnSjGUGjmDmNWv0KQyHm3bG/O1VIeuKc5xqO9nX8+P0vQBr4B
V3XI48FQh7HiDGTPm336XWw3fHRMv3UtAVJvGUX4+QaGmJRcUwfZIuiHzKitfEe0pG+8y6nyjoe8
Q1O3+2pGGn3h3xb1LxSxNcECoUD1vcxyy6t4nv3h4aJPva3UWrgpVEnnThIoI9322mVW3DAWQWVc
22gpUq/WHjiu5g+IJMphsKVLDcT4capsKwPZVRgOGMPSqhGEMEVX+KlIDfPLjsmqUTPbbNYz2i+2
7ZDngYIcZw3N/Kx9SCwxO7ggWnsfFliFbrqDxPD1x1Uqc/lGbu6QOGQ5mPTlUaHi4bjXS3HEj871
ZxXIo7qA/f/uT2UuQpcbkGK1FfyLgC16mfQ6vPfJybHl/0yiTv1rEDBaE027uD0NT+uEHIBePQwH
96LTZvQjEg4Uxd/yCj19EJViSZpTAukKS/AofG+VwLz0RWHf9xvzFwYEch2hSCvIa/Agj0oQwwf2
HwJxerQibr+0lffTp62PwuwVLR9Gfe9hkoYo8AHwHscp94eg4nIuF+H5bQqRZZoGgbILI4txSOok
89/zHQBJKCMCJWtx0nzBI5FbIAg4l7l7y8qur3U5YP9oSdMB+rNUM6tFZNhU1sJBtMZKyQNW35tC
ZMRGu0xMwXWjnmYXlSYuCF98U7TgHj2ZWbXYhE/G0p5AQBRAcg9BZ/E76/Ny2hE/6uWKdAeryYK8
jQ19WEs/SgTFLs196RhQBKgI2DGk9vIwQegMI15KOdF7pth2ScFiepbo1+KLoeelIYOOB34fuGxy
7pCjxqJyU/BbWZun4v0aqD6Irgm+WNMbwMuutjK8l+SvooAFBlrJD7o8Ss7BY7ZVK2WB82OMz+/p
55T4MA4w+PPDkZdFLHn8l7FtGPEOxNteY0uIJTTDEClPJQXVXF8PhHwzZY3V+uF1URYg1rG8mTRG
ga/vwpazMLz7E2kc5ulPJjfKYdQTHzadPsgX115EBWMGOKw50MatJZZi8gc18ZFsxSH1FlxumDIm
Uvl7skgHqqz9QpqJjppnKhEB2o5Lwj30OudB4iGOzfx80qVd+idJdEsyamYwYN21t0tIKEV9di5Z
Fqq1xUH5HurAQF1Si4uu6sxh8FTF/UuPYsd0eBty1mRcdLXOtEEQcK25NVqUdBZsMF1fyPhZovUD
zO34V5LLtZg2EGlr+Z+hqyERv//1e5TsPVOClO1nZOoLxcVmuf+hPhtf+02me0zP0qtHLekjgZFZ
00RCoS4ywBQXPR13z3gh/+Ouqbb/2e4k5SPbAahxlDeC8jQO7d3jKubwCAZQr1hDuu7yfiS6E3xU
LBROrMoc5pIguZOq0IS3nedAsILR83gjiVaJ/KvlVWujSOtYSiqhNgIU/ZFlsFvDi1TXScauc3yu
UqWNjhvV0qV4qpdE0JyyfZrj8y2wEe/yZg9Y2aKFwE6O5lWweiXF2ljub/b6k6QjUkmK8tszzXmg
L0oHHszi7Yb0Oynls/gZEC7JJv/c0m1S8XGXLYUoqCUfwgwh9C0PMuWbNVutXqmjuz+pM+t01qI/
FH00VYRlEvH+sRPzr05LNMEp7xz6LpxTWGDqNLIXaH9JavfP5j8zSsrXEd7vez6zeUXUKAXpTFCw
LCdwacE5yqMt7Cz7bhhFEECs+Tt2Krw5qvRmOUmIwKfZa47wGOGVJWx6S7kcIIW1B229ICCtrydH
7MyXn+3KI+HI79Pc994dmaOZCJmTIRFmpylhfSlHWebg/qh4KeEUOcb24qhPEcvUQjpr+ie3IlTZ
SCKku0lzrPHLFEndkRy4XjYvlBFkU1oRTZGgEmrwqea+c+bDW2pebcBTXf2SxScgUBM5PCqoVmNZ
IVWSlYhMe3I+n5Qv6w8cqXfxkwdRbkjMB59ob4iT+x5uOd+S9Z7b01dcesnvrKJbhSLoB9apAP1D
rRz2jGJc2SP9LBd2727b4EXpDulS4KEx1KN7ZopxgZeeSEY+Iskw+faYciwAb5VEIUledyZOJ94b
L/FU9TihcQhylj32wh2mG01lg/ogdT2s4s8unX9jsjUIea55E5eL+wLJqAW4h2vZS3JV7M+R2s3+
DNGkjf0TXli/h2MUOSlHNEDqV9LdZct5ckKzaIlXCr/nJCjm5UDhgcrFRpRB8LdhzfNAh9gyZgi5
YSpyuy5bx7/R5bfoWHbEO4CzKMPuhRjaEHc2EzYvxpkg6O2DlVlcH1tzBYs0DKjFvMNB+6PIerJe
bQyOQdfFnk/bzygQ2LwrUPcHnqk1O8RdVPnz+Kdltu6jJIo3tLBop2mOtIX4YwEUT9lqVnAajNNy
Of23C3M9hZ2xMRJoc/X6AHuN8Ss//X2VZhYLtOAh+y1IlZpvIYm6Xrc0SV4GqGUaufwOPmKN4WWA
3OgVRugHI97il+Fg9ldTF0acM3gaUuoqT3358rb7bCjjNSV7VjvKOiKolnpCyteHDa/LZT9y9yXK
EAzmaSoMRcVOA+f86f3R8ukWr6z5+NCmGDNvxOk6VdA7cGsPy/LFEAuhpb/pe/XzFioOKj5ydrZe
J1dHoK5wfB4vIlW+XNwKy/iiukBnzC4cLXsDbyDWboeZttRCLuL1aBBVyXbLks6YP0INV9KLYA/t
Cw8wlQE2y3y+p9pV/e9Zy9NAnOOGS+vZiCxbwRKwN+hl1h1/34lGG/S0mXAiqcGBvhqWCeEAa4Fm
3vqeCCXMFc2kaiFrxJzszN8w4i0Z9XH55ytOEObLTExn6VFonatOgtTgaHUFb/PwCptt/U2Sfrjb
MzOL7Iz7wBS49I/oIptOFOGyoNJqsdjP8KKhU+mceSONzQEe1x+iIGckmDP6dfGe5kUjxtzOpdyA
UjUCcibHB5CJmRSlTyAuJ4Y7A5TI+iAGvlhFvr3gQAb5lWvO/wfDjevNmy935kdEVeypsUmhLTIz
GhI3FQ3UMoYi8PJTjLn+NWoJFfIkmYYLFnJZeBLIu7dsjxMJA7r3amMvXPtoNfjccVuwaed5254j
W7y0MHoDMQVRLKQl8HOhTt+U+MKP9yk0X9Hz9cpqeI8/Xo0m/4IQHr38XDxah8pyuirXJiDxHjgQ
Hc6thBedB6eKXlCeC7u+mX1NGwsuiWOmCr0R8JPeYRA8rwd0vhS4ZiFIclZMrOdYnyejfzgjME13
8Lf+3TfWpfgxVqAQ7BNeSjD/43qRfOxJvYhLxr/uBbJxJcb0nBIw+jZemGCJLFuP4CXx60Pk+8o/
FCDTqY54WvFcKOa7UbVTKeln/QTe/3eZwAIxC35HqAXRbjkLGZ0IVHDF0Iq8VVYZk73wB10Is6bV
KAZmkzoKMwSMQst5ZjJhKaxOeJgNrU6/RR+q3kocaZlIQH5xNL+vLn5DO6VdVAb6dlh6p5wiOrW5
uEvshoDUkatoa3tAdOuvtl5uugQ+zSlh2/5UB9q9ANEzd1lV34T8vy8oNi5VN8l+uMK49yfjijNR
wKM39Og+pF8q3H8vlozWpLbA3k34S4bJtE/Qy1S14F4u1XqqSsrcX22/8cqf5QUjJwRYJLnXGIW/
3u/Az8y7UmHq7LD9LfgYcxRNQ10IQoAr2nubsbCeyNW9GebwWZnEfSS+ThfjGf92MWR7j3IiBl1H
qm6a6A3CDcj6WmOVBgs8Ma374snV1NNXYQrn3czpDxddkHa4YNFiRcAS7B+NJu0id7+w8IITYXo1
dn6ka2Xn2r1xAggiLiPpMR0ctbgZ63QXRItigUO7CtoPyCIls9+Cy4nd4H54etNBHU5XjHhS/DKs
Qvcd/cAcCAioDmjJHJauNotB3uOeYGJbk9FAat8u0j7H9GEOVS6/50IeSCb21U1DPf/NUd5pd3ZB
/+XPCgKpzneaBgKSQlszIZSTyZ5sn3S7UlcI0X+eKjrhYC/3KD7K3KNag6sAvWrMT2mXbB7//aO1
pxFe85xY1rOypy4qIlNAJfixtFemRPVE5Mf2z3hgrBA983jttjku5D70dRbzFFI4B4CjMcIpPam7
ikQHWxr62Paz0SEjaYOO/yuEGLcm8dRBUbjTbhZXPe9bRQSljmm8FT7JGOQmjJBN0YGpU+9S69Ds
RRXGlI+94/3D7SdnRCRSPuTIjmPKXR+OASldHqsDcRGaBkQLGW8iTSN7r8HH4QzegVFnw4NGKowg
9tG7M25nWda4Jc0Or0zKtPFYMqL63VP+cgatAiDbs4ooJ6tTE988Siuzyq0YbRIW5RUvJ1jXwIJG
0ksjvt48ho56aYy2sMphnnHUvxx9CnZfrq7tTzW7w2zutBajz4GdE2D5KpgC+3usXVt4LWb1ZtGa
xnqIMtJOhOOKoSXibpl0TFpWQ8uPTQNMBlm6xbZQMt0Tdl3+YzNzHRN5P6dufPZjEsOPyYoFg97W
ffpfNKJ2h7Us4Gi539CKg560zPgZzsfnfLrcqYNJ1fm3vJuP5eH0YqLhOfOShCLsPQrBmFHXPHbA
593OVxFvFxxw2ahvvO67xlgeEEdHku3vLjlXxSxcLYsjsWMW8pXjgQjJRnSHTTgL7hdHcNZgCumS
afr5dxhO8/ymsjQEyrKfu6mBTavfixKbnF64diahXEE++WdhTWiJRVxosZRUlQwJoIValloKyXUv
d/sgxU/9GZGHinY43298J1QRDdWQoWPQBJKlVfJIlT2ZfHiIrZ63Ezlnb1kGTLvIqXIRC6JtJMpI
BPuqsizn4U8iDY9bE3v/ab+UWihTgj00wY+c/bWZDNiP8uyOcU9UTE4KbGPAIp9PrkVj5uMw4WFi
0QhnlGcaVS0fIwsU+mRLB1m/+6r2QmSjIg2SCz+P1kjC4HD6QuzHDPswz/3osHqgVTyKwg1tFDFP
n2SC9dM2WbKW8XFxHD8OBf/YeZZRgufffpoo6wyVpLcq3Txljjkz5tbepE2Texn/E/SpR0yLhLAg
xz7IpqGt0l3cSi8Iraj7GpqSURz2NVVr1+DcGfrtKqBaUPv9UQRBZ1f1UtHTo2/yS8DYIFemAhDT
zfnxgvKIaSpzS9meeW7op9ch+wp9rTum2PaM5C5vfNhchQh87pu78LatdYjFFUbnovU/d1Fsh2rX
VbUc6spIe2MkMehLYKqHFitb25ODw2WD8WxYqvtAePNFE8xWQ1q9LloTSSFB9fgpR3GCdnwrw1lS
E+TElp3JQe8tWBbnWgO6gxQeQUZop7OKUl9H6uP0MNsRGTkeAOHpwL207K2GRjouFZVUOBZxpwHi
nm0HOkuhSV7CSf/uOCy5M7q+iXEwQLL/kSopZoV0AzbP1e/RnzYXy5aEXWuZ0p9YrdI1+gw/F16J
m+XxXoCRDDuF1S4qBibqCokUak3flCxr0z+uycUrqzMtkWVfD533LQqH8MxJbMpOllTm03GyB2Jk
nHqGPRb1dsH7qPj7j/BgBL0sF8h1TVScsTiFlFNUwyKb8W14M5iuwVuA4HZWjep+lrxUuuqLBuOp
ZqfZk+JHNCffX9uwmwhDaEpBIc1LjB/Sr8+CkNKGcnA1JgJPw8MEWhMNbzsvjjm1H87/DnpP27y2
46/ryrD7O/+U4Q5wl0J85GG9b80I8tJC3nzXyOvVGU0w/+gnGDOiX851pEzfQJpv5Z+m7EZRAyKp
GPgpKmK2hOGH/ULPztubFaJeOpHC51BI567MIuSP1Tx+FYeSToH65OmFPIep9ANnl2Mx6aEe/SE4
ZDrvMDRRwYT6y0ZsiFPPH/ZDM9V5aLcCWI2LVmZxEUi7dyZUZad11foigUFZeNBowJ4b23B3FCty
RlhYwydtz0wMLO9sXtLhYC0B0vCIcZ6o0gxKdc1qOEfcAgaBFcVGoQj0dH3H1/UsEKuF0OyX8fQV
kxDkYpnJDu8SI6B958+iuhobzdTfGzXedrSF4FioC18NIjtEhql9dEdOlH4L7/ojW2Q1APKF3icm
lD82gmwm+JjU78WIEewqIcY5w0gnjtRD7H2kd7suziF54iWc/K158c6UHwBRLb/IdWucU2DiS7c1
CYqLE048xj3/1s/3qvEUAyfbCwidCGEuMovgUT5f9k41VFwb2Qs/Zb2obJYUrWKEBD0Lqlf2usB2
yS5/9VicnGjJ3kGufOwaereodfF5NHQT3Ff1YqWJgcyPCJFFZxeLLLUO5ek5b7uAUqUvC2dxSnJX
UU6ij3tBvdzZvg54t7XCvZEAljdgvJvkGnKqVYGsFnltFuUGyOKPokMyN8fweczrGs5CCF0Aq72G
LCEHMsMAH9HPkRbza/ul9/HPbkL0x5za0Lx2PoA4uk7mzRM3zhSeJLZfXs9JyVn2LiaxNK10K9X+
DQYuWhXjECb8vz8+7cQ8MawXmf/OI5TnF9LCJMmTVGCYAyj8o7YNXLiEuG5jwLzXPKRQlRSBglc1
l5pr81ZYsyXMBy57NpN0hQG4+spQQUBOu9QPREFfWxMkFJA21zHoz4/udcy8/BGwXS1cMivL0+lS
YFzMxb2f3AaNrqgydPqXsymZMF3PcRe9sZzm7uAWStLRVUu0KWkko3Zp2oat1KhvKBI/HCNCAao3
RmVSnSKr/u1D8TqqikK0LLPWku+phTQNgwsJdHYbtWA05NcnaizhJFBAApnf2CQ0kkj6roq1W6HJ
CQ8rfAu3lHTeAB6nTMJqj9zqBdLwDP+enGFFa6MCA2U8cjRf6LLpMi8ne6C2kbUGa1P8aHrxyijC
zGqqxZFSFEnDtQCYlQ1cLcrjXlFk1vYgFmKG2f6qi9fnEIJv70GiMIzKlCAj0yfeZec6sYQrz0NW
Sw+oDHVW8L71mkBKY5zLQnOnX2swcR9b+YWbqzDO02eDmXEIIlUVeJcgSIPrpDEXFBLA/GiN1F9g
hWaKQWrQliTR6cbrM2L23ZYC/dCW1+tOXW4+fthThhBUqUNhNb6y7nTv2w8Sw7qQyG9KGNasY5jI
27rAYOX4hwh/gH+jDyqae12bMAYmPAmWiBJMTGcL7PM0mCAWYfv0t79kSDQ2d5nksDlyiX2t1Ceg
VjkkRW/AokeTwZiAlQcPGEV0JLAePzf4t1mFe1SCxKd5puLRKgbymqM39CJYVxAFXWWZ1EJgf48x
XnM27blVEkGOZucVIMwL756xlx7p4CIAHplnSe6wrgYClrg19MRsSYjSqFRtK8gpK/lhtEERVmwO
p0KdIO/J82rCW1AcpNxZ3jWbNHv5GTMAfwFhqmb8iXKHmUsR2kzLyqQ1mQ6wPUyJa1XAIcfOM3VA
nK83MM9OBKwFk9INhwO/TFKRICqgNBZbzihk533zvneeBjKNF+zxmUAZy+tTr8xYrYmV6IMrh4jp
JJ99PIi1WTSh9KcSSRKWMRS0/s/b52Qvim7O5hg2QUCJUatWIhyLLyX7HgryRsQ5bTfVQbYAj8Q4
zeUWapV7jHr+SgbDqvWbTXtHCGToy4cD9G+cugyprMkRcjw22DhK1im+k46vPUH3tmyaHXYLFg0I
DVFEU3dGYugWubT7M6CTYNvH4no00/qCw9tCpOvt55TbACkuw2saRVAuNv0uurZfJjCzcuKN+bl2
REsE4bv9yTM5xNDQmhCURrvbJXn7pb7UUbOQgWfqlN70zVOkWZfUlOlYK7WXnKft+bCRK3woozd3
zzDz9FkrbAt38m3wvcaHqtIvo7a8fVLvFttwWwUND0Jk0S+G0O5DNSyFbndNcUe8Wp/6F30MUBRg
BmxJJIGpC7usY3yFqOal115LZg/unsR9tbHJTaPJmVJXp0OxXpfU4/gWWt3o2Qte1VWtjiQZjKuo
xP3kgH4VkNiX3aQGknZd5ovT/x7Owh3PgwlYoJ3ECfGylLU5Dr75oOJAIm7DJEBBDDD/zXpel9ey
Q1U5Sc5754FxjD6hA6vBcNL0T/Xk1c9S8KbeZV16elsXzqL5U1k10StRmkP4IMfD89PtAnQ+lwzu
bpg7+aJiiOCVGtw+rpXosSGHjX7V7ehDlUkszDA//8F4Kb5UbyWBF3L7xVPW8eCgNAWE+IGpEX7j
P97hvZKRHiP9V5O3t2w7w2szL+jzBdJ028s/KF/JyHwwokOhyVriYp2k2Cww6UuXzHyqK68x+ufa
ND+UuAGwMyX4lACAxxNTff1Y0Hn7PjLq905n6sRMR8KUXTOWfjVbbzclWo0qvaLDYQstHbmgxE7D
8zO5T+V+KYExMqUm7DFpw1PR2gd6S6EEvRgNkrutdq6+9WvsiN9e/mepvv1KG9jIPfuuNN0F/YRw
J7mweGhxExZ8tSEhijHYqAC1Ndu0HOYvdgOF02fdQTLSPafLjXeTAJ9d+3cg4NY7Vh97CwERQ+cg
oLxJs9UKOp7zq3Bi15/7mpsTbyOIxdAO/t533c4HwwkhAogFjTrdUjayzhAn0OSL0iZ3SAC2PrWs
W0Xt4RbbBzwQJ4essJfmBuRBVEu478F38XlBAdWvQkK21uqQ4G/Edd8apI9Cp+12M5WjgPx6YX9V
2sWszys3rJOptBspStlEWLeUx+WY57lupEswX0BPnAXSMi3w2uEFVqTj38bWNQ5Fe4Zyw77ERuEO
clmxwGnBB/LzNKR4YB6Znp8IrqOcn5Jqyt4htD4hQvVq4wIXTPrez+s/vhsS/KkJl3xbYQKLttJc
mnlfLQkVw20xQIY6UoM/R46DvY/eDhWRrwWteWlpOUpE6yGr0/p5mzIp1BaiMURiqPd1aKKfq2xx
0pzTZTXRty3ZEHqMONE8kFM/F0ogVKFAnJfrBp6piDrNWBV92MsA3KCmmI1Fy5frID4X2ETv6L7W
5hRyMjNh09tx6FqG2Inophu6UK0ChIdkHYAsLZiSAXR/CgagaDemV/vzqBdjEV7HV0B9c/u0rO3I
0OwwuO0KUuLggcpFbjQ0L2rabLYOhKdHJckPl84ZM+SsICckUsGeSaz/k6IbGsP8EutlOjt+TTQe
CWMT15yHCfbmiTXYoIsU92rixtri7JQUzonHWqzM6cvCddCTzJnuyz7JzJZgxJCX5IxUl3+9+6s2
fPdU9KyGF1y6LXblObxW5ZJOxh6+eSakSQZvTKxSmlyxoeyB2/3mbF1deHeX2nOCJmOyi3/bU2NO
+gFWmJWXArQ2vugCqOY+IUEFCFDWXxn3E1XGZOoE8jvjJLSweKNPm38A7wubyNmOmpf3+7wkECKj
b2TqLrGeIa3ZcFhCfMrHGIYkk+dCCQHVeU7p6YVIgXAFmP8+kXPejA4UYCwsTRerZs/gjjuVSUWx
EbJ+ZyqvpIhThVsTmiSlPU3rsGkNLEk6vfiRhrT90DHY9Qjc1RN1M8nMw5BRfRpvOF8cNh64t77s
32rNei33uV+8UQZdwmLhKHTFkrty3dvmfY967KbaHsLNfFEji5fMPb2zere0cv15lUOt3uTmL91U
5BzVs+Ui1/4gceiCaDgtRGA8JT/OwgE55WedAVS0m70J1FDv1OYy3+dnzSY2k2iP9XSePC1+pfpq
CgKzx98NrBUXVAev9JcsnefHx3g1Fx0juWEdGuM9EdhSdG1vyVbe8uJ/fTmew6+xX6HmX0nD3IA9
kTBPUDPaCLVN0RSiYkHBg/tbXVwtveVaktEPmMMRpPZ5Ejdl6CcVmkSMitz0kjnnaEWZMEcLX+Gv
M/iDxGl4IrmjdnoAt2Fba0g3l6FkbJqGU7KlAqY00PCs9xTnZMOvP54MmKTwP5ZDdmBrO6K3WU4g
ULyQ2aSPLD/WV+Nf7S4Vtf2JuoUkjG3zp3u8enjBN6qJpfxeAzWeHLNv0+3MguSVeAyYzKoDHlP/
//oPKAR/lnJQhJDZCJHnMfNCGTieNH4l99VQ1zbfAYLC9x5gxEtDGOYXpIGyMRLGoUfPa1FuR7nn
/avG4sRaXC++Wv1R7uvk47/+vSlcdO5FErcdHcBoCCJopiK0xZ09/Yy49zpThHbyyytZ+C0qCpiR
0GQ96EMUz+F17gJx+ZfZt1QQxQ6Le0tdlmEtFCynsD2HARl51JAA9Q9asz4HfpQbWqm7mcwgmssi
ZsJ1bVBjrwyRWbVjvlns4stix0eNo6h3pHi2vHMCp5ABiRVK+FpYD8cvA3OpUtbhGpUWWDJHenFo
zoQuDJzf9N3szRVh5mAx2ZyrgFtw6ssK5BhHiufsUE7TmP9gHSV+FIy3Sw549Yrl5xsxJ+j/SOME
Vvbx9wMCJG1mohkeYqWNdkydkp+gIADPDLeXjmdftyD2/t91EjFZog963TO6ryKMbI5hKLSC8Isg
b8KyEdAgTGGrCRDphxyXEbhvBfB4TczQy5FEZSXZU5Kv2P1kZUFReweJLCN59alvI5UFMQ83DXY3
wSt4AWzawjfBSuLqyJ6qng5fIMncvNNJxWqnYvRJdjZQZX3PY7CFvvOXyLzvzUmYSx77E0dCNC/6
KLG1fZ9p8Aj+dxFzas9+vf5FxLuO7lKiKKNHfb1vl+NEgBeUMvwhTrftqhsfcg+Iq6cWuYYxGenq
rxBP7GVwO5wbGmLqkKnVFFLbbnZ4Xw9DVj8duhuqE5A2Bdqpm4vZh1nk+tfQDfYGvxjpgv6HfBJ7
28Gmsj+wfTjGPEJw6Ej54/GT4+34294yOJjhQfGRT+HfqlNTLTzZ2ErGozmVLnOAHwK3aU7InWTB
XGMc7JD0E7Qpq1Dhbt6yh3AL4HmP7JxJkaKdKr7E5lJhOjb0FbQJMJoYDsM4fUhVoz1iQeWHRq29
xk9wO8nLOUf+JKYEN2Iqw7roDn6xeYEa8keIV2KHI1EZEoaPd4boSCb5U6hNMD8aE7ZAkyPkA3e3
gTFSV+NhArJHBmUQdbacEsR59kHqA40eweZdQOB2AHkGJ/P4tKy2iTZhmYQW9RsHowNarhiXMgpu
Jg5kW9aX5UfqDfGfilyLS2tNvUAUR8eF8qoPXMh6YLGSh/zHDTG5uP5jJTb1bjMoV7q6qN24MhGV
nkEKrombu5Q1Q7er92jFxT5AMhUkyYdgajFjuaiQ/NB1QwVMFn/E9LXakESPyXIZMhrdOACJjhJm
XtCx8TLbTKbeuYs31rPZPCtKstihE3thweL0n/1wKvIW5t5pL47MkYXUxzsn1p72x+OABrKx/Fsn
TmmQeLSHRr5kzu0AFiG+hrXoxWH/VYnUHPZysAXor/9hUK3jpZtU0tzS/LXr8B1gH+uTL0vCLwhK
0oyX2Yrq9pH/lpRTcIHvbAaG0jew1MgbGSZfwYzWsRh6cuv8GkWD/GqGCuhp+jFqV5volcdtavmU
2avtjhpm8oSUiXInz4WOP7svQPHwZ7kyNuHq77TZ5zgzaeDYsaUlTVVXlYmwo44cwom3K/Bd/azt
6XU7df7IGD6KcLvyfn4QJgE93Wzoq/aUOLlXZKBhTIGuHVc7WJYBicEVrRKLnXChAs2Ic7FVgQ+4
Hd9RC6+8J4fub8RAfpfUiw0Wmj/e9Z4aCS7ns2Bou8IjHFCkvYlFOUY8ZvwxLXOIjAHYE5PnEeTV
3jLP6Yh39s2HNlwXMPqsZMTwA9o6h0sJQc0Lwt4YAqyTAGsn6TTC9YqNyKnEAIMOyHS6CndtVood
8nHbEI+fRxCyREXinOe5J0fPS8Zw4vRp0JjXCduT17/ZBZVv/Ex+rw0XcaYWZ33zZkXVV8eCcR52
g0shqygO/ghgbusrkgS/03dpGVNAQjrYGsFO1tTCBKzqV+h3J/2OPtsutpKGjqIYZz6lTgq4FJFu
V61o4wjNaLmS24H5uWx24KK9MRy4T8r7dEFeSmCSzeqpRiUEj0nbhZdDl5xFacph0nArWtPt+QhN
fS9+/NMU2b+X99nEbkY3EOS/yaU4q0hXs1PakrVb9oUuQ/NBM545GTMufwgM+F8wHRxCD6i8rHzQ
YFw/212SvIFgkS3StiLNcu9BnOZnzWpZbN5y7oMAjwJzHWL5pxBS0rkrwu6UK+NLtLl40Kn/IxxT
hcDdCgRzoKRWKVzL507ILj1lmCnKPFVd80rPEOzJwXhmz6BKZHoqf3H20ffwK1PKJrjbHt+ZDOBL
r6Hm+0+TiIdNFtwIfbEOPFJH5Ojr3jTKw28FA+EE/YnjShcU1Yj6OqpJYc/sJCAT2awy63laI+Nf
wwaBcyUAkcLacdLmWESacsgnd/nwpFI6LGrBfrf/tzB1lowSVmwmxUsMUcL5H9LiYEPbpQYFXUMC
dEBP+H+5r1xQhLqYdGZ7j8OiFASj9JGdvr3Zwx9Tr5U0c0Sjt2mGABkonH2CJh9se4fBKL64aE3M
kkTATjYc5HM4oJ7IffCyUuAWfqfIdFt/r53k4Yhi33gLgCZ4CyKDSOcoJsOLQbv9XufWQYRXQLDf
N3VFxaG1bAfjTPjnqXCmkmxLKrPdkzPhj/oXWhUzNkbbpuxfISBXoMTJa3234qzoh7uwy1Hfwfr5
sSYJiTPAalg0UzWtz18PClNzcJrWW+O4RCruPyAu0QilBwzDsck/UuE3mCJXaxr0JcMPCTxONGHx
UAxFzpksPx1o3m7TTSWNXEJkT/5//vemkY9904sp5mpUw/BUOlBmQiFKwi5TMkHEPaqVrOfzHNdu
W04V9Buy9Wl5ZkQpv36XlyXIgHj8QRyPI7LcAHjpKEznNtp02MCtCYuGsikMclwrFfHZADP/ar1T
/ySJo2mr/elZG1/+xBrw/Bf4hgtpWqxWqethLnDq4N+gZs2CgMjq6P8b2ynVUvTxvE3iNjULddIg
rQXX5mHEe6MsAXy56O9OXvDDATW7lt2coOgN2QTydYqy7UZ3MUZhZbTsss8xzDOdFaouX6d/rRPu
EIegucD+/5lwL8Y0eG54PQi1GP0m07vkTTx8slLPGJNYR6PNOMO3M5Oqbbli9IBGu9+Yr8KkM4s3
OfJK1xNN7jtF/AuTq07/UMc1Ha3e1/az/IcYpy8coL00Y+5R2n3V3If5XI0IURE1teNDy/anRfZ6
Ram7e7oMcoujaJgbUZiHBqTIL904NXJ0PsU4SDzzQkURd7SLjY53HjXS+PoYqw7T3n2hEmJlzJl5
NCa5ScSsiJvUp/wkt+jczkloo0Si422oTA+EVQvZOdoaY530XUz+FFIBpjDTybf3MHgbotNKHk8W
yvREO7pGKyQ85EIHvM23dilLg6+Nv1XHP6xaAfGgBPEZO5k5xeuMRzE4PkRPKxEeAGEF1wItpwkH
lJmGzcxrta2P9Xaz4fTVYhS+259t2t4DtmuNrXhdj2CRycgMwsxSx92NkecxOWBxPaMbJNcPYXX7
cuckqtSI/9pCkxIiMAUVLO2G8JTUMc8bZm1+LsQNBrMNGMDGmniifwKMH0VY7uI9iZK/9EWInWya
LWaPH/1bZvizJJxdyaxYOAQnjhaIOdlAQENEqk2Nxac8KcdLF0JFvZGF1hplepfSAGuxaKLfy64U
FuQeAZHRioH6wNbm/0BgwfniArn3i4Kp4KscTxd84P7dvRyiAzKleNQKk+0ccsmwiz+uyD6X7rUv
sLMfckVqoVpxyDhW5Sh0tVMHeZ/2xTL+J9qmEzYLaJNu/1u16Juuj8m/0n36KbEsQnISc7u0EVch
Dk9oWdEsYW2ridYLc7Bx3d4CU7heSf14S5GzGhJV+bHVqqW7VqX+3Wyt/jgRapPOTeVVvkfXT+6r
dt9KaGtCJX8KM9qon+vNiuN5Qu2fukqKm9HKPeZQuQpt5oxxpxVXWEv7op8iniPzPH+ev1fFglx0
ETkmppQmH67vwjcchWRNfBdLIxiU5QSzi63pTBjHy3ZGJpRvr+RFFeP71xFJwN/WDxX5mYzW3gBf
j/x1Yi7tYIk3djb1f3YXD+k+4vbFUXlkIu1ZATUMpmpFrpfYYJpFpSZfJAO9lhKisOYn+OkhA8X5
4ZFFL4X99waT/99InnV4ab9aZ3VM42O0ihiJZ3nBhCiXGAwj+2SQCYhKQ1fn7CWi8QwjJFFwVVLG
V8fRPwFqtrPaNgFRUVuztxQlOF8JllDJlldpcR+nP1PVJ3Qe2CDsq/37jN0VFFtumGQOKTP/RrER
VJG5ipSDAK/rPFp7Wx2cwPZT2DsG0aRudJ40M/cYFmaN/VYSxRgtiUpswMCquybtHouRCtsnjCTB
6HszbovMka6UGlCPU3EfK22rQN8bwTfHwDpErn3MOCc9D4WEAJMhkbgmr5h2SKJ6nM5zOOS8+YqZ
u9qCFMcBAmU3mF8TmfAiIACCZKQFMYWMEwnVneKXAcqfd9UaRWpIDGGpVuD9nv7Mq6yo2+n4GzT1
75SO0Xt0Q3rxwmWuRLSkCglNsresXUKEJudI5a2iHZE0NLB1CRwpvm0EHSDGD5GYQrnVl5hnfaUT
CvYhSXu/aNYGH2FMgzD8PbkhgbcxJMTFR2hLr29QEwilXzHyhERO9rGJC2rzsl3xwAH9eGV5LcXK
AJyZCBAoWGwt13nbmukaxe852c93kTtwkunlj4sVN7iPdKDUe3Uxz2JJWlTyS9pk/0TOZ5huxDVM
BfB75EJH4/QjX+Fg7PL3RvVaczvVgpDAtjuTs0/QzG0HJgM+PxkzdvnqnNSQbLSWcxbFtAbs6Km8
FlNF1CgYc11Gne25s/kb1WyA1jwjVv/15kZqPvz6lP6UvBZFpu6guFHH4FHTBPXoaHQhDiIancx5
h4UHEricRg7I5+aTdGTA9FLYGKhMUH6+HKQtINAoeHjXjsLeiP2PAPPR0vEsUxl5ncD+SilMaLgx
RiVYR9dcglelTq81wohTec6q6OKXGF5Ds7eG6LNd5iCJ/5u4Ci2OcZiWhQmzyH5b6aLzBXlSPJoy
40KXDmJJmhwrrrJ3tFj/ufLWG1krzdUbObrDWQ15uhNItgZ886g5NEqn436jaCtkDIsGEaor1Og0
ulX0qxCn/2ZqBX9zuCydJtOYBn5lB6E4uJMpOObHVaXIbCTz5SYrMYJmsCBvm7GX/m1tAnMRQyHJ
uaFEs5sw4mjiPCLwmkdCUtMkw9iWCJima0hPeQCxsNt9/TwJN/K31EdA4/BEmfnFsRn2eP9/QNdB
ziocMkyHRearhHxPxs2umJ1eROYjm9T8WH7COdLkAL9lPI14PR3puRW6O78cPTqc/0gtb3295EB/
ABUIDgvx4y7W19p+kq7Clkx+r/5goGPBDY7F37mbcd+YADUyrPEj42f0hiP3Q3SnROPLMh5t+f47
2avZIfl7WBJTwCy/qpZE0MSG5xZjWRoRC4b2GNxlBUDkzsR6xCwFA81YF7SWuqQDHeSjrpfQqSiS
Ab+5lyXyJJykyM+CLEdqdL6xoacqLUee3YtiV0Lx31OSxUiUGvf4vm8Ft5N/fjWWCm4svXH3zV7d
qqc77Wa6JI/CDqDY1A3oAv/EuVk+w1iqw6vIeQf1JM1wD+sILcR39jZxcCNV5b0XCS3BhlXqszAh
TZfsT+30uzrIoR6MrL+IZ70/v1Kjk/O/i+ul63EbK+JLoRFg9uSGnQA5zz8UMU4cr1amYmsO/a/9
QFyIeM6mRcoLqN6/XqTzjtXIesWsyFLVPmb6t30sAEjChyUpk7nHp3+h+ihgYBNAKZTtKvmG55ev
KsNQ8d1JdbboIOFGZ3JIw8y+aIp4GF9Yx8Vnje5E6RI3ItZSTMEXlQ16LQb8R/rd3sKKF6t1rfN0
HUKTIproAoK5MVJUB0GKlnX8oXtwYRPyPqD7hk+atKglIKWPQXKwgs48bkgc9RxvZwe5rlOfkQWl
WPZFvUMXDnbDFGkiIiIaEHhxsNp5n47eUGB5BkI0NKmLn/KBxdppFyCYod8Nxtf95XxDDGgqsfvW
Pr7YGDpfQkz9YTu4nWXWpmRCADisPmZJoZa4PxSFGptx0btKM4chKy2x2Vm/pvcuUvUOYjEUZlqk
7b0ZaP2tU/E8EPSSWW9J05JSKiTBDyjF3KN/Ds89GeuWgpqWWQKuPVaQNIUb6/Ej2CqwNrQRUykW
d343OhMxYqXNbIpZ0+pD/6rz+LJvB9jrC2h+StX287R1BqtbbKKrOWlJRwgfzX0+5afySyG26hFP
sCuKkEuGWs//amPs6NAJiyRCq/+DUnUBk0G6Q1DG28uuG6xi83RorcLo9FJ31qFSjga5NfqRQ8aG
v5F0tJB6bqrmX3ZcX6hJxIdj9oENlyPR2of4lakSi7SPE4M9+XR8d+gsszUko2f+f8+QpyqaCkhd
B2uMfR+GY8uy8pcric5ditHX34Hrbg/w5KDaiVc6uIcFYWARGqAPCmaVmzBjyIu7o3609hpkDX0d
/WFdCjrmsUv+HyuR/Oz6K2lGxSULMupppEkfsZrqCCREET/Q/yn3tURY/L7mDWphXMHHIbVoetv/
rOv1+euAxs8KAt3wU+Wo1PK3+T7/NtIn6MuWHDaiQsudwqoU7a5vMlCEgXQ1RVoc/sAjpAk4OYTS
d7xwYHa573V2PXd1mUPixDPW4BvPWMdMAFeyuEd8n1zdc+W+/HgX2bkOU86VdUTeU4vS0Jr/tFQs
ZCUIaWvLU2bw/xIzTdarlRpvzNRizp2Mqjr/ekydwNwbhXVRsIC4e7GPSMpyuwQGNZ99x9EFMNmq
Oq8u5bd+Rq6OLyBkEIeeyqvtb1PmFAUvIcKh9PKJrQVmcxMTJ1lyU8S+GvvQZODZqrV0IO9mDr9p
3gtabF79BdFe8E4v86GK+08XVGl4OB6fDgkLBhxr7VwuvOwWG++KEVVTi0vmsPaHj1Iw8bHGfbsR
AvpiprXtyxobVWRrUrw633GsF3nXkibXXxGwJWEev/Q+tMZ9cXTvppE6g2+XSGaAJnGyBXLfaLRD
UEr1mQ7p8TIPjV/tZAi+OKhceVwgM+JUzGyt/AcEwkeiJUYNSJi5WNBDdK+wrpqCuTUiiS0pOi4j
DmEoQkkOd5mxWYOMmEsoig70KCkoVFX9h+BPv51fb1q0ugayj+YuC+3kYvAMlgJANuyg0aw4S92A
6TcKibRjsBBmvc86FIZgLWCvwFs+JAr1pL8O/8ybMQGN7dWyirPsp9SIW+D1PPZkZSoG7C6LE/Z1
wycZAk3AjvLvJFRhfj091kilpbj4aNHmgh7UCS/EyTVRCNgTNKJDZWyga8AxHghJNWjGCbqifOZT
+8EweRuZh/dLCQu/FMr8/FP1GZZzCLCVn8FCS/bw6fHRa6xSz3ZVMX4QW+SYESwro9AQSR3tB2Pz
CklleDfjBol4w+WXYHXi0wkOtjExR270ipsHITzp6qRN8HUEZ+nh8ptgHTQwcB5Ayaqr1vja9M+t
v3VufZaANozPv0R68UwttKrZ68CVTbFPxHNVauiRU40wKBhJkqgknTPYfSzaG5i4oUz5y/JzTz48
cJUXzeiSSN6awwHRhchuNp/6QuWbQ8UmEiEK/znBP2JhcNX6s7KJrM5++NZm9VRuBL4MThGbM7DQ
kMxvGERIicy/VVn8JlGJuTLVhjIQee/sQR/e91J4+9QnSr/PAXcAcqZ3ObVibVijwED3IP+kZOQ4
PZ9h8vTRlEWogkyNUnMj8GtFfbUugfOdqzXw+2YbqA07hMig3fVuCVGFyIg0rmpjSCg8uaAcc1Gi
arNOu+BOzFniII2XGhb08Nn8ys2vPA7vCA7lTPF6CYhl+xr4QEo0GlVBJdySNmMkqxpwbhPTIP9y
3zI0d9Fv0FN81CW9QNTytH5o2++PhAIQoOnvXh9OabauGhspoFrMet/UWh+iWywuWKFqc8WCfnFR
Ch+62FVFkA05h3beiPpFCkTLvl8gWqGAGjBse8wMseDvHNNbsJwR2YomPCilrb6fGCVCJGuQFCzm
+v/SwtgVDL+xWu0OHyNmXXOriozjsZxNORl9IrxWpbbwgqbjO7RA7oom0tr4xm99/kt+Br8iIMDd
z6KQnK5V6Lo238duFsuGJNvWch73sDEDsjV/+uIf/mFNfMFRLD5dYhPoO92wUQt/H2Ynwl6/WvK1
b6XzIVGM1SHJbObnqNPoWB0QeW4w77SKgvcqL9SxtJ5quTD1P6DhmLVMrRuER+7PTuwiRltZ1ggY
V947ilsX1E9/WcdjFoY0/gyyeGRaPVlC1F8WyUYjHkgrfBhSKHjCVjOak/hF2t55SAYkJFUnew/4
ZoDL8cMbFc05/Tb69r/EfoCOmdF611PzQbywpUMnqp1SUcAdvmqI4TKwtmZW4Jkho+oE5aEEKZZs
GhVv9gO5m3xO7OHI+PKsPtlH0nW9XWpLVySbSDZrdIBYKh4gHMv9b3HEJo/+11v48o5LG6NRtVhl
Xj9fVIYUPxxsFxqIfQ3syYM8IdxVqAo+mB78KbkRyaTl3vHMcBO02Fcx1bGqihhQw+dinuUSF2X9
bXOQxM4aFivDAkACkM4/dfRC6DAPyOOlcifc0MgGPh2y0QoTjf/i0C6adY544IKjW1ZIVvFDyyRs
1/CkK+EpNIhGmf9hna9sgK7tpOMhxTF4NLnpeWpVLMqGSMEETxvzrWKhEUzSuTo6zZ4pVeCRK6yq
g3fThGLURhwSvM5tsYPKX+qDnexqQy10vy4f1E5NLNq6b8X5vwV7k9khJK2Umc+iteZItWAJonbV
yE8EiDm/hGF/JXU0X6OyW3R+NB3vQ/7nCRYsi0REWJFpbKdrqzTu5rQ9xxzsik2VUGZjePqKJhRD
6THoO9QCBo+oIAGGOhLB+XgxJO11X+HMr/VlvVYsC7F2Nu3ey0OYrkY7sjuu32rAD7DucxnjH0cI
wf08UUFxwLI9+gEJeTiw72wdeB4WygxZMeGBqHcZ2DONKGazhfGTrgThWJo3QBUEhKPJ2Vj0412n
JxWodB3sXIwaZjma5QqJrXbZKuCJ7HO7FPjBVhQ+/+o0xJPhHE9Q095pmeZ4OtYdJs94lsR6LnMH
q1rFTuNaFSffPkQXrjXdPChYMLPqBXd5TivskStVLsAl3Qm2p4O9KPzMU7A77l1Svmw868Ie6Y78
zYhMZkytRwaBU243G0PG2yrTrqJ7TjnA/RAD5vOdqn/jEkfQlSqpjZIM8U8/7Q2IabCc9PnfY6m5
roWiL9kJcH43M3CHlo2rG5nGuCqA2cLO5K/1og0TLhZfWFvgznTWr4ViZjjnEJDTCnDFSZnVkdfG
Ak2cCrFPpchGnQgKyYYLgXWFUiIPb3GdXfEZkS2UQ8svAhgE2OnHqrTG1k2HGUGgN512DjhDPf1/
RmRxUHYhNpNag2/51TVrNOmF1DX09A3iOHcdwazWUcifUtEBCaDedxc0kb16OxhF648tK2YInB4T
FQ8YBM0LLNV2Z049xH/M4NUZkHZoGh06kMoO9KRBMo1D9hSJuey1lGN6bT60n0V4izUHG/AchIq1
z6j+dP98rLD3ekh5Ejjaf1W0DovcNIrTv5Gp3XQ5rUGIbRvfmKiLKJ217nTlK8MpDdjI5LkWhEfJ
cp3HQT6kqDzZoyRaWkDKvtTvVWGi2dPAvBxCqacnVy6uMaWF55Qagb+zdjkeSWMp/D5GSZvoZnYe
eDPDxkCnXsulpEJD0TJGRKy2Sd5cYrekvo4bQ5znoYKnO+UgU4s7SOGRR5vRGT8Gj5Dly0Uy/XS6
6+otjbgu2jaOD4hGn+af5GLeKdkqLb3LoixHHsimEpnZ9nrIM9ZJm1UrBE8J+ak/1bHhTfxxXiCo
CXqWsw7BE/4GNoN8JCdVqC7soPvSx0Nv62dH/GPMWRetZltif1YXVsngrEwTMjtvDDS6t6Obj3B0
AXnrFvXpNFEKifnzUkXza1dm/T+GEG/IP7egEQC5OypRjfHdiyVluIsOIYNCw5jl7GKrpJZ9Fu7/
+7zMMdjy2GQv1yoFFb+PeRhfZMGSvF+aO+H6hP+Qj6zkk24msRggWdKC0jjbLGIgQrHVf7wkqmQh
CD66vzi/J79kdh2UH4VTTMRgIfAKdfnZTO5LEpHyXCb0oQ0AMYnvZA3GCtPOjbCTPBhKCqBg3pAt
iVWYgpabFYo1XFhR1rOTHBr9vq3b78MJLKWHK3udSVVWg17tZI6h1tcrIwZXifYiaBbxrCMhZbZ7
7mclHRKg+5aDIJAl89HNG5fvEHB+fO+FUXbgbDleMUbbNmqdJjj3GngagIg+EyP4Zj+KnBzZvzHY
4n8Efxw5/yY50pWE+zMYpPmGFyzbQGQvDSVVRcuM4yOGKJ1eHA3yGgjnahKJ4TcBrOAu2tM3oTnN
EXyBxPqmIcfXw7ZJ86hNmRbcgJ401fA4LluMHnCA7K0Meyyt6ER6tDaDxFbuacQA5nb37X2hMQl2
sp2bfW4uYc88bf2tpV9W0RVV/lGXAklU4VZPHB5IQAizwwL5qUItSX5tdhnZnf3gupT3EhDQPiGq
CTy/L/HFcyzVwOdL/2ojjgJ0HanOLB3kROSEWaqkM1n8DYJMj3IAJqVblx16TZVCYDhcJi0N/MOA
qxwFRQNjZ1XTZaGqzDyvpcfMqeANFEmYH2YHLICn+UHFKPtxaR9ESouYHqX4XIPtcdD+afHp+Gdo
vyFmKC4ypK+UB1hVQI3htvkHCyVI8/wsbeFb7NBOcjZRS7oM/vlZ9EbbjBbMBupNpQ3ZSlCgLpst
1F1sOofBL2jeTjPKv8AnTTMFcl0DhacuufiRdclouKv9eDSF0AmQmb0L5ZgBgu8yiOGVQbMxNc1C
EwIYsWbVlPYTInhkSd8dw87GguL/takuC9OrJy24iniMpzBhiGzSfkyGunRCoKK4kBf+E5SrlmvQ
/Hn77nuSkI1G/n3pYO/jCVUsbOcCM74UTqG4TCHS+RaHzxcWrPSemh+aTt9ChnxnlmIzB6mfRh5f
7cC4dTkdcBhNixFwtSC+makmPIy9thR11SN2Kt5uVc1v5uqXCFTE+AFf8xlXoZcx/tFo1ekpkeh3
R+riYXrVy5vzJJxbvPb6r33hNRQxtBiXhi2Xyhng2pfJYFWM7ZQ4VtHB/eZEsJr079evnNUf3MT5
D4lynVVxbX5g6sSZNPZ/nxbGcKM8eQk9eBaVp80VRGWGxI6OXgSV8RaHc/emMqSuylsa65xdbhST
E+N115vAJo6nriRtU2fxCtYqenCe48E07tGx38dc3N0hYanNI1LV5hS50UQyIqmzTHkNxypdaXTE
CoYS7hFKfhSEqKR+hNejHZkFZQ3c1YwrMZ0E5I6jjuu+Coe76SMBtU/j3pi2VGvtE6kjfxjA8r70
ZDxSJdNKZJ5YGyf3VYAT8nP/INmtPuioD6Ez9n8+1zDYKpvrF9oiuSY5pHQHJdp738PDEAuMXtH6
up0xmkbNdjcC8WAVnnCmXbOXHhE4GbQGJSl5QS8wVslCj86gvBIo0duQ8XsbZZnv1A3/l6S50gha
sI+iN0hb29WOlcJDE9knZU7IDek41hlmiFRRo2JAgIz1TOlB5EcJzlmBZelK3Io8vblQK/QRdRlm
Jqb0J9YQxC43gwET1fpKDmkZbc7uTpSavPI2PNgHu8ovAJwc6l6YalzzdvIia6aMKyogw9n2lSmm
6IeeJNnFD54w1E3PB3Gl0yHPBvtanOY9vXlxfxn128JTbW2GMm4V+HX7jibrg4MHTXN/obHN+vvC
z+Zh18Ca77GDIPsoQRsOE3nAabJPnSLgSZFWc9zGyDAyzBKsVY1bJa/1JVsKPJQdobmuaXNoFz/d
j5XD1JVyJI/ysCNHOR/6/mbYO/ExjP/F1CCQSJdc8kH4lSN++9QVzvwHWxMIbOTraQnWHK8VOjhG
Dv/0pRHYhVn9zzo9Io2XB8wNCtRaf8BxxmCEPN8jaq9SUYJ400WBzTiOLWs+iJJQMUj0e3DiP7du
jmaSVxLDJYXeMWqpgPczPBWQOlv0R8ohIrfM/3dvaEUsmF7f/29S3hQI/BKxYlnBx7NBlW/XxdBV
yYegAD6rd9oL1H07tXPid9iAnY7DT016wk/hHR15r6IMNZT193NF5wdHB7ujg56VNVC2WnglPfqj
JSlq7cKQKIclt26EpaaZ/N3QnASJQW92lWcuwIR45ZyvA2GRlk+VZaT0w8XB2MbU7SIekRwiO7xc
TAQWPHhvRytz4RdmMRR87N9EQOzD+P5E4piQFAd8uXTbSmx8GiXml4mtVCdxW7omrZkurMB7VG/D
QLSXYbcXmOt/LgAbhsrHOtSIh2rZu1yK/0IOzAlsMJE9P6NP9iCM7LpfD83bagk2VRGzC/8kOJuT
UDYUB+CCPq/+GRoTmb484Sv2SJn4yibtVP8bVK3TnwgBZ+bgOk2WBFOXHLpKZV36MMFUOEZqfSbB
o4nqE2sY1YcRC5n0iKV+Hg9GIbNDF0Kpxm/97GBbyHHAUcIul+pytfVmYXd9DF1H49UfR2ld5rmA
5Lx5luaQQ41FweK020kJqSEVUQokdfOlHWv+xNdmqzC5RxcD/w6WcvSYuPwBRAIhMT334DRgOGZc
kOJpTuB5sCPn5MKLPZ0y8UI5mPKgPS/DwKoLHXNuROMP/5tr8uQ78UYuoK2YUQ2qtoFlLXwtXl/2
W+j9niv27MBtWQDXU5SkyNxVDOddBtY0GhXEyS+UZty0MBPqTLKKNMD2OrZUYO/dHl26yiuNJLcr
EdLstmdv0nNyiLkR+low1b1DToSr3azrzIlutXbvCd6Kdu4ADEuDgZFXYx7mrSfyc9Rh/16DnYoC
T0HFW9EGJyGqneNtLl2BAhsY0n1qlyaeU4fz9VUUpYYOKSNwba7jWzIr9yrXK04ZFvF4ju4VtyoW
nLUd8sYU+lrnWS0Brdk5F7FWbAdffMO3xpYnm/qAmMuoZfye22QGaqb1IwS+iOBkVzHx8Azsg77g
d8/VOfGl1gTE4sHAJFwnBjsQgb4sGGAJgYL7IiwlqOfkTxbQqTuB90+XD0zCShM2FheqcBLI7vjK
qGkyV+9z0JrLFeu9KzFqE1vZlTiqb3BqCsrDqWHhRF12wS+eGfXfUUTV7XutUXIAKn1ltZzhNE2s
2PdMhQBljb0ikdsz1rg8RTHMgXPncZ6xYKXxAuyCTYzFl/+3T4XUTrbscY2DgkfEQ1bkjEq1/vuR
VcjRNZ5qvPocSNPksTngDvd9s7ehfdHW4xzgRRSJZJv3GVQIBaj1bXjF1cjzzbilYPL8yEOeiZuk
2XCai5690aLH7A6ikZiGm5F9RbrGCfb9plbe5XTYKcGOhyijRW/zaAUIgnRh2wIyk21JCMGqmYN+
0q70v/uk5qp5zK4ue3bUWxF3QFI7t0Vqhl0/16T0BV6VVGUTnRwbwBTvHc1ywyT3INLTkeSg3RKY
gmrXqmAP3jc9itzsJxyFiPt61aund/LQvOGnQ4f2Cu5AnlcMkc7JG+tn562+UbBs0MutNFhjJY4f
AFo5Vl4Q6yLD7sWrXICNqIyiPZ1jwBdO2tL8jFnfdqiug4oDesKApmWwynZGxidlJTpC1TdstSsC
HwM5txVqsKDsNyd2cpgTmYNjGKU1anigmDOgyxlL114lAwo2u/l8jTqKEjwoMdrcKOrh/rQva9Dd
0HoEbBhFfdj9hhBiuykSDE3t6i6ErHBYZmf/fqiDhK3ypnGwkTSJW2fJ2QgOlBh1iMSbRfeSVvSg
usqBz4+hDpCv6ctt7vMq6bYcwEdepnfutPqK4mRYRxFuZU1gXr6h+RHcfhBX1snqhHeRcJ93C6xo
eabGAj+zXJdwsJuvJYZH1hsrtYDrMbSaDlS06PtmVnL/qdPUkflbQ+8aTVkmGmPnRRaiG/ewqVIV
0SoFpjVTIeHtDBTpe2cRUqQ7k/onkCs+b61VYxb5ByQYx532YZAxL3BExA07ciirbDKVHM+hiS/a
YCRpt1V+NagKXqkIh2Aij/tbZPFEWv8cIHq9tvXXjIzmedJuYlSVY0oe/t6IpHtIVWIgTbGXaTm6
yzg7ejOJ8frgl6272sZKSySnNCalyu0/I0iTyAjOqXQE4ihilv2WsjTUpGV9Htf+9dAlG4QDEkW7
K6hIwPEpNvrN562vLnI5U5i/Hwuo4iUi3Ku/8bwsRl10dnYWbxTRgfK0TxqaR4TvEhGcVtOXGBlD
KvX594U9BMsoVsBWusV7V2rmdJRvyrPmd9xCKBSsMTRc5gH3zbzoGEj+nYXQ8HzTF5sWXpF99noJ
Uk+k7AiVpfWWV7QFYozmos6JeGMSwYm1szJckioNNPtUdLEkSNuljXKaK5u6ewqb1G0DkXWzaPXb
PoJyFvn5C019ugbmOxW3a7lEayahnWlHm5Qy23t9FpFt0Xj/LhhFG4Vy8a+4kc/qDS2J9ZGMVggy
xsCg9DVrxVa0SrDa9WuJ7oKrYjuM+k7Q0+d/vYSs7uMkfPRv7zCTkvXrfSsgvhcg0kkHUvFjObOP
EmWquWTIytjbFQ7KdfOOGvlN2GNhipL6vYOQRmQerHa1ncq24u31534ztHrH7zmN3Y3/ad/lphpU
RoydHoe/917KhS31ce4SiGWqhkNGnAV0D42e+lv8FstUmxgUtt3iQzB9Qmi21KZWl4e+36EqVh2J
H/3+EgVZS0UCAvxNcwLVs4tM+Q1LkBNhJ7mAubOBhXfX0G8o+3mKwP2A8pBD783echwzwjz4+wbx
mb/ibQ4gUFsH0uPxLfz1FX9mNJnl8YVrjaOvnsEhewAjs69bzOP+PZlhDVA1AsCrMM7VVHU4nvxI
1C4wmGH0p42Fp5P851QixzmIHbDmAJVbhEitDaNSHnDD4h/1exHiLVB/h4DcQNKENntYkAeLy7cA
SmrS5SWhMn7PMsKVGwmwVyRy7eowFyfNBjCP2K/2pvB9/EvsUMgiypnoHXd3F58cM8EDb230VpBi
kqLCcH3+rJ9mR9/ieMAf9w5uvZbmrR1jy8XK7kujV6YvoSNpnYAGdUsTx+HjkX6dJMeRCFveBJLw
jB/SP0/FfpQhh5AaoCeuBLgOAf2xyWlwIrov11q3YxxM0RvD+RS913HGUtIFIVXGoSzh0D1HqRkt
uFFs7QFhU1EdX4ZWlefeMw8vNx/X0oh6fS+OS6v+fegE5Geil8TghhrwqQIDz/79RdbAiDeibbhX
1zg9c5qYXjlOfIRtj1wv7I+UMF151/Qut0Kez/WeqowPbRBwm2hE1Mk7LdDYcbnpBilUz2GWYCWI
q7otwYTuu9r6RJtFZ0ciSnQQDZZWn/EkORt19fT18MdnWxT1AXXXEeQ04ryDqEsqkF3dMLy9YaLH
SmM3JKiQvSf75gcAO0hwCcL59g3OIbYGKbKuSvE6uoFb67RQXRZSl5R9/78s2T7HOAVI2xDKjgGv
C9PGcws1cpTP9IycXPt5wEnNw2XTPkM1hqx3i8K/nhcGtilEGCysUsg7PsaM5MwkuUOSlLFzMjvF
NcA5N82naIcYn5EMFKfHE5P1QdUIX26yyeMUPC6MSMv/iE/GOW3/2bT22KDO3AxDOmbzuODwrVDO
RGg5ODD0263qUX/BLas84Mo7xw6aPOCBlb1APv8IkpXe/hZtFFuhBuz9CftNjL6O8u/xiYwNREp+
USCwnL7vV0g/u3KTj31BWBHtuHq/Fsm2DIzZjGH1XeZWUD5nONO1zHZQDrBVnHl+xibpg/upHYb8
/csACrluP5qdvYvbXlC6WZ9bRbRmI6BiIYKxs0gfca3x9DcmIchQrC0i/qYh37bW3DDmAKfFd1k4
zXBgPL7BP1BWq80kjFJIdpNiKTZraXi2goSjMXboh36r1Whyz2Mw6X0MdQKtXNL4bi+nioNNZ6C3
CLnxaMpsBKwtdUQ6rTgHaUZwgWcmsAnLyE/QN0S09dUJi17deVO5eY6U72WZlG6A6CH7cw5YNL3I
V3K9dls82KETx9jXl0QrQIH78XqBSMN8lntbYjME+y9ziOXeb7OlxoiDObAhfObrEenG/vt/1G1F
aYsszSeoqga6ehdLQQqqpUk2eKnI1iGU1x94HrlgzbOY5xKYmjvkJkeiaepBiYFflTKvldg1Zud9
TOSeCL8mCZQJlIYFnN5i7o5WHlH3LefbHomJjoYvW131/Lovgxl5wYZfnkBx2BSBEEYLhA63isyj
dxKf4IYnabcOCDPCiQMo50DdMWZg4KSE9kXYqKptxayi+YwQFPvW5Hiez1IOuqX6gobsvVD714KM
/ZFph8Eha6Q8xdPVYPZD1VadaE+E60yG0bYcADkkxgO3GK4J3kbwgDJblWpEe9Ehd8hAn9WBCXJW
T3qi25B9P2EUyOv1jXi6y4mIVomp9u2LB0spZMWjo527/SrEukxal5hdUP3RTzyU0c4Y12vKNkFx
X08sWwSbrhCC+bhpceVMhlPKrmoEce1LCeQ+3yxpFSehD7P4LcMyOo21ohfI25XCWb4xDM8H90Xu
xs7zVae3JvySXAvUxxKOofwCPxbq4IcBZkACpkjQGCI7A01/2arMIzgdIqszLY078MZticcUJX9w
CQbBVK/h3DCTE3v/W6AaeVkJ7GeUIrRxD93Uajlf4rJwd8KxBd66+pqQnVLPbBxaWDRsyYBFlLhX
yN5/iD1GQMrwOs9/aLuLF+KzpJpRmF0sWzzhugocFepC/Yj9plkQEwGZQCi3OS2s2UkEUv5UTN7m
z2ZeuHTjgnljTRZpz1X6nBCmXFp99+WleE9+ozKI1OrPy2nXTR0JehWCqI8TFz2ZesKYmeFgL75o
AC9YA06DgwhnVjt5olFE8gb/kazPiOBohB9PJlAujDdIRpi5gJFSHJDvtyyfcwrptnTmSYa8Mq7m
LBMz7LDTLqPHzKSlftHcbp2QOnyo669XOPbvO8b0ixZWbzsqbrRFjzVyouPXLMg6ZMBj0glE9UtJ
773iuCBri0dS7QRFx9rDaziT5LUUSaf2PGrqNN/cGS9orHg3LxVUBo8W6TnytnhCk5e6Gpveic1Y
iIL1y5VpRKX24ErCX2syi8wvnR2bHbaIAKPnACZkRDvbWJMEmdgX4ufeNfqTUVMwyQ+OiBrwFVRX
Zd9j/ORRVEnn8S1TROkKsRyL/N+It9V68n9LjOtGjr/3376QWLsuhQrXTYiyrFSidN3Tn8v3xWKB
4beN0aHTHdhga8CGmZ6CDU+8IngcNXLAdXlUIRUNl258jR+IXXj6f9MqF4wo2Rg7xkdpCmVDBNYw
UjOXRevEDjAbrmTF5vo+KdlQGCPYUTiATs38maVM5ZN21sDiywTH0WK0CqY2wkzf5SNHWs9RnyNq
UKX/1pomNHCRqyly4WFCnT52uCdhbFTdiHUIq9fDIAUc1ODu7GBqF/nSYdh3ddlodFh3XEaJ3Gnd
2+iZB2e0nqH551chUyXC9as+KElYNwYBkfLITPhK/1aFc4VenagzO3DC7K1rzL9vytTUTHdN59Lo
alj9oULWar7M+PpQwI9c9AOa5U5n+Keotl5D8l0qzdBAWRnFPWnWXotiiBKU+eiM4KeSl0n8KGoT
d9na3o8jZns1+3XsgPwApmp21yhxHquJhzsdEOYfGiyRb4klfeRM6Nee1stOEn8ON6Ty7lElu6J4
q0E66H4QzUfgjVJYa/hG5XxqXqvecHXV65GknaVFrG1iJviyZfS8pKhoVCC/8dRsvJ/2dEafi7pF
fgLTq0E+VJ4oVVABB5p1PfqVB47MWjD5o4wq4cN3fmPnYPWWSZhkM7DpaRvjlNAixu6a/tBTyyTX
kqjnZ/aUsqqruf5r6wcIKYEbgQJLWespXBL3DwQuN5xGOK5m5F3VbLMuREj04R+F8VcWKUaEhJih
RWL06spJQIYDGF3retm9APaeE4Ox1WGpTCI8ccx8wb8P01s85ODIlzqiLyKJFhlwF0d9hBTGumLD
qCHave6OO7HPITSVBt02CPa9xbAeqsCs5X9IO0L78A7/JQCMkaQsLtW7CQKIz4GrktkDhD4DZiDJ
u0batZqBIS2WRVnKq5vyFUAwyVyhJazqWy9fjFEDEPY4RBjbIaM6tok9dQKbybwcD2f2xi0Q03Go
pdYh1DS/tnHDzotM11ifqtSF1HKG/cXxs09edUw6CSoeqpNQtWRBuKyFzvZo6r2gzsV43CYRuvdO
GwbM8XL4QHa1X5Nie+AJCqHZ1Ca6HU/xAM4eUlavy9WDeaBA4UjnLwVlJdFKkNOTbRhUg3fc0WuA
05Zh3+drrNwAZ45acGbTvg/SrOTdGYOPvcVm0A47WGOCIusH27CwrGOYxcocBzu2t7jFGHvqknC+
1vwTFkef0mvHsjORWunyeK/ZmaJh2LvKqXff2wbgtbKgju5uRvzc1rJbF6Rx96LWZl5PPPr3CYxd
HLLXyJ6j7dviglOWdku5OgKnJ486nqa/P4mz5NM+FT3PGodbfbgRsHHUJdYgbLgxE0mwAJ8r+BO+
ErRO16CUYoFElLreygAPvAf41/q3ZvRKWv7GEJsn3/rS04F8wAt+f+udSe9bwgV7DFj/sNuPj36i
fBnWH/LwJRNRHZsuw2xqNxSuY6DByifETDK2X/l/KeDHLTL6pBDcragwOVxPyv6dOi4VO5AiYQnz
G6Aa5uclxnQ55O2VW08oye3ZGmAKWd2G0ZdluE1oOgr9z5MEmtr8vn/JwI9EOLrjEt1FYbqFTuNH
/H8C7e4p2Fo2vxGiELB6+obcojeQPK3PNY6k5N+0XXpCKuk4r5AZmXC9d8HAneL+RaoNrCgYHSNi
G1KbS8c46v6Mrbm3I+OhmgbqijwM7e+OlxFwV3NKrk1s57G+D7lbcCKKY8af0HNygPPuVVn47dYE
CIyhx2/lplFzzIuO9Ka4KUF+FMvAdckpAf7v+H65hXUwJt2fN/jrqvaii9EOBGnQwWsPzThvb2u7
LpZ9/9jUn6A/zoGuFe5nXiDBIYut4Az+0FEyahJ+izFOSJcuXbZY2M/FXFYOEEiQPL+vazPyx0Bj
sa4ErAg9gEymvp1IC2newgTNIMM9ifdWxnSkamfRDvxTWalFJTCD2kfVGPgJRNhIKZD5x1t5dsxO
tDaOtK/sQEcYQis18iFyOy+Ib/bo8YBcwkRzsxsQzAHlUfMnLfE7rA7xNE5SzEWn6yISV5Y1S1fh
qIdCNP118kzWTztzUF9bijNp6+OdVd4473Jl0AY9/NyL7DnbvAWOc9UO9kDrPkrr6sAKUe5kV5pY
s4uSu0yU0MDATIDQ8ccRumXaol9wxMdssmljkJqInJG6CTgerVXEv+Zh4R3QCWO2HgpblOlVTV9V
NkeqY+tFXHEAuuPcUhowHdmjcL2qAMYbnCJ+OleaCLXEqD5anZmBPsgHhMSAFdxA9mmUKL+wZJM/
ml+cWyUdnonbRpizAqF9Cjh9JI2BDnFsKvcnugCzBqir7HyBxLcSlSJJVjc/Jve2MqdLdgYH5uDF
yAG0NM/eB1oNUFSfcMVKOrGBXangEUdITRpOurvpceEiAo7L1ZOpMfuaAjQolu2svxRdq+MlAoZ4
4C6SodrvQe93T2g2s2wNr93kmKT7caPweH3bhRflnjkP0jkv//ykyMt5vZwpgehZSEiKxhTduJHf
6ctstk+Uqun6jUjKnWxAX7Yp6q6Id9ppnnN28rPWerKJaNMOLebS/PbVXi1jn/GA6Wmds9a01ZJG
QfUiIhVqCUreJU60U2GWQTNh8evPp0VqRvqr/jLi4RB07CgJKMRDmdnwjgmuffj1MRJL674SYHh6
eZI6NH0iZrzDD3g5rthsZT5HhRpBL4IPoSUFdpVAvptv961roqfQ66v2dG4G+50Bjuo/JMfP8gIF
WxLvOC4mHHCR6/F6K2noj2cGsk410ov7TpLnULToVRR1h0D66chELVNXn3HQBLu0sFd8KRJxRUgk
Hrn1CaUeEn53O+wxesbY7eHPozQE3ysg1EfSUDHFBsiTeYYrr+ybdqoT8+rkBKqj3oF1UfoGrQau
TzhRyo6cEwWGcIVxzzdbOj596UBZZDaSsJekkaO10qLCKlb9ba1eXJvgeDUWphWpcGESzZRFHu4W
QN2zXdFW1A9ZUe0QrFDi0oC4KcnaYXRbsLz20AWMexhygQ7oW5lYDbNbdu4TwDhv7KLjcdyMSJ2b
9/gyzp+gRjWGS652c08xjEqfMbRBB1NON4NLSC1Ywbnv5NjDIy4QZiQpTCR0dEYyDGK/kTERjcgB
tj70+p60IpGeYD0/vf16YmEEdq9r+8slSm7zFnrOwEfpKzStY4gbnRnkMvZ0I0xANng00sQ1w67l
g+SHqEtwlYxngy1eLP4h7PkDL1l5Y+whp4EnlfwuPgBjSu4jaNgnO08KOjrnlfVmLePQjNzarKER
xvXJLyB1VNgJEIZkcSxS0f9fX/TheoZL6jdMfKPoq0BRmDlEvuoclZl2ozmdW/pKg7lXscoTQ0w/
1ytfka998J8PmXahJetxL6K2QrIVYWZ5gVESU0xVnCBKzJxgXSgGMf9dhwGEny0IdQhLEgCX3uOc
EU66nEDosNYpBy1CTvmCYKfBF6+s7G4DOe45mKf8phr8OqgiNRcsDgAuN8EXjYW5Lmm9gPLnCx8I
Ofq/qy2zDD3loHG+jfqR5LVabo2g7nfKKLIEPNFFX7H+8Vdnan6kctNPg5QjfUTQXNhNbemqqnV6
Rg2gLxiDmb/fgrvZYXc+HrPYtDDbv5Ij6+9SvkmEs5Q2fz+o+XTcvGb2VHKyicv7RmFfNiVOG7kn
Dp/bi2Z8nxkwf4xbgOBogOOTpbvR11x06Ij2xl2EB6gb0/52ONMTrbZYxfhnlaiHjQPtfLR6Lpvi
kc0QZDPNDTEqTbRgNyqes5xIBTnPWk/ZZqvph5aluL9fbhN/HOFIFL018WBNDH69QsBpfH1eiu+V
ylcdW8HVzxHa17Ro5pQFdaAAfZ6jv/b/3wnSu3K719aTzWPXhS9eqeQ5RzV2qEx/KXyQXJSSmL0p
kK/vnIL48amEnQYQiSbLBG/3ecR9qrqNFRgEfLlOvTOj7M5RojDChzkh9u+aKBdbOeEV123VX4af
YpGCWpV5HZzxzExKceyx7rdsnbGAxQmvsg2Q056Mo5VbaH9qEhUlG+4tV4haSIQSvCy6o0w+K+/F
9KrcR0QOIYxiKcELH7nePQtp5Eu6oSZtKBh7fCflGcFmq7bR/q+8zrr3EIv8mvEGg8mdDJEyjTa0
SXffXWNAGnT7wrmHThxssfB8ZxCG8divEz6a6dirjlcaHFeuo4zgUUBWWtKZK242GjnPr2N8CGA8
MOf+Lym3TqfIBgLhAXTMJtTv0LbNqop8eQxWIomkTnTDEFFzunRc45OqGnxEh4K0iLeVz5rr8sdj
SFE95ohqKr0LexfAa3uj+n3podr69HFFo9xLHMWyOX+q/qvmceqbZNhLqvsSDn0phXcizFRv0wFH
9/yMCCRwko26JoeMNJYGtQUZYznhIxvSGELyUFGTL8mX3twAT4DHt2B7LDaleS4kdrAQj3pFUcOY
Nb6fdu3yTKMhwAybPIvMERIcps7Orzx9Rlqrkl62n9v4BtEX75S46Cobwk6a4ULWrMbVi3ZhkM9W
c39KcbZYON+Kee/2tDJ1yAOqnj+/qlzHYMHIehfRzMIAjpznh2zUS7LuMRZiUlNPNC/r7dyb3Gmt
F5d2bSoB8gJWUImmzzfmzFIR3XJIGM69ovLCdfPTtTicDZn/gcV2qnCRuVEQozX1aCsv3LrzUaLd
LEcm6hGt2+0EYI1gWqFij22TscrUixYZD1eftNPBnaES3G4/IaNwAwtw47gkJpQjoaqK8KSZZc98
m/xNbbUDa3kqdmISfBkiUKZKgBn2GYEz7UlM3njiTLiVXcT6NT/hGxNDQROq1nhl/4NOieIBI201
l/e4vX6PxWAsfZC2slm9QZy3wOPctglV0he7DsyP2FG6CMWGg9qGh7zDy+QoHLlXP8wGDq2tRj5a
MvH6AxENE6WR2o15moYD7uUdU9qanmB46FebS9LIhj9nMg50H7fmD6Q0upz3Nw49x4on3wld1BWW
9bbGHgZ8r2Qg8iuquaVuUoELVuTJz1yB6K0DHU+3qaNaF5UI03bjcnC+Db5GGtnfnEq+QoKdgf6+
KuVsG3czaavnHecZdTd6hcLtUqCuQv30jtJEJ/fRSBwL7KQ1jRSI8gGlQOI8QtfomI4YkBdFEYRw
KXNNccGDIRPBQ9L0k89TltQS3GYw8V7YzT+Ed96lQTjb1LhWc9rWqXqEbs/gXZex94xASnTf880f
cT3KWJZZYcN3+uJe0ycOaoD7BoT2om3Z9o59UoPp22FI6w+FJJjv8m1o4B6Kh3CrgtL09GYclAkv
+rRVpeT2OcPjhLpoSMUNul2AXlj9C8wWYBy+bZ9MIYw+7BmFsI/fOTjfHjAGkuOI5zTHkDWlUUOa
swIqOZzr6gF+gK6VuvVrPkG4J8bpdSFXgRzmzGkSuuMooBaOYsRNkh8Fwb9PGG9FsOlgouRBW90w
c3NctkF8Na76eo1e9TuRAWneTWFcfCJxTm4bpK2n1Iofa39GYphtGOIjddrUNCOl0d6TS+eXUByN
GLh6hLfmzObVtLRf8XbrYC7OtmM/XtT9aZcFIzXH/jUjkrLlf4e1LE9El7ARJLi+4mpQUKgJmVx0
mqzK839SiPvH6D50reOkpqlj09/UDnA3FYVo14Bi6qpejZkkj5pbBr/7AnIHtbLO73XF2+lJvYRk
H/bfmJVgYOyAHSXb9cvPhNtON5Jthd1uzm8emad2coQvt50qDsH0CxL67/pIKtWoV+RraaHDx0pl
A60vvxXNkXqwkxma7dC8ybCB0QBlSrG+FdwWXfhIt6tdi8ZRBkDHW7xNDEohdmjs7V0bwvagDP9x
HwFnVKuuiB6MR138gFuI7YiwuEKKwlVw1FV1ZdWjy2aopgsdxfwlMVaSu1Pq/ljn4RGUv4pdEfYZ
g2UoLqpWhyiS1t5CY9BeOKYPMEeRoJJ3LZPJ81hA4CWjZK1uISKGyKh3pzCBuSOw4tu/E6V+NM96
m7QcA06FyJwaqxA6nPHvjOyWmZkbnevDN//Wx/oAzE2zP8U2EsMecyQAaUaYT7lj8TYkSj0Spp8N
B8CL+g5b4ggg6Mj4fF+USpHHLt8+1PV9p4nusrxLkVckLzhcfVLbInt9sTYJghJYXWhyQoKgo3xW
wMha8FOu3H2TDQguHuh38JtiX+ritFbNuzxybIQr8trzOWC6PHk1BJqTWNGeAPW6+dLo/mkSxdaB
tL4uOzGykGaEDFMz5Fh3NWmYkEajCxQWpd1DOQS9IYTq29TlpyPnrD+Klov5wxnhVUihZ3vqVslq
DoWtQnT5DV2pDjka7EkJIDsyY7yKFI6hD8Tf3mNooOE71/mb9PUIHaiyTWolopDTE7ncIowuvG25
y5kYgRNE75CJUJ+7Gm2IyU+USD4b/g3eaXrDZcN+squzEKD3sXWO5E1Uc7v7+CREG5AxKzGdE7uP
wo/WQbqyvxBZmDEOlOG4PouKnysUCF7tz3R9lsY1xno0jaX/9qNd/d04ftiBrWxh8KV7NTUVtR3f
+G0OT62npc6t1jnzpkU3jsj45zT9v9S76cbzyYJTjZ14RRsWDBkT8SzWdoagm/oNiOxygtxRH3Zz
P/dBlfzY7PjrBxHSS/r+Dv60EqRLmkpXebpb7ssgCU+XcPZp/uTW60pVaLdvLKgeQFi6FwXVhrJ5
BGFc/h99gyg36q+oJh0EYCyFN8C4/wnr2DTmWnac5A2qY0k412kYVlGmoVtzn/IAyyoAoM3sokDV
1MYOqjCU/0eIEPolAJZftzVW1lAkjcaOx13ijlQGPPMiN6NT9kNraTjyxXQj3sozN1JWX41GIJ/M
Ii5g0YEgmivgT1UWUewKiYsOjRFZUI8Z2bER38xbSRq9PyMvGXYQWe2QEtETspuGD0qpFGZOMT7d
zNpC5+27oUmJDib+iCS9hBJB0HpX1qg+uyUKc+aE07oQVTg+8AYz7e2eVS/Qctv21ZTfqNtVMIoY
TUMrdBX/xr6Ly2xfA/gmM7u6OGBl2ClqYG2/4oTvdYWZuNt26O2Y5M0/p9zYHIWBBF/y6wIWnj0q
i5ybp7k55llXltoYokH0vGioXBVnF1FVC1UEK5pIecUHNsTV2NsevxnJm3V44rrT0cVxC+WvjxTm
7tc5r98N0DoV5o10esQ9HCTFGhlL6E/HJFM70YlcXEhvH7UQtIwRDWMLgeCRAFek0EWgACIvyZna
aRdhmKAsYXKfTYlAtvEjQrZNRNp7VZMqjxUP3AnuRoqbxw7arg6BatKchnVGBf0/L8CweE3Qmjzk
alvE56y4A4boaZwDOjIMuYx00pXiEfr8KM4hmPDaJU9TG8iTshH/kWB1YS7wsi6hMu5gmVSn6Ml6
yYbqsT3703eZ/Bs8nOc1IjW5hh+PV2vXojSdejqQ1z/OYZQZRpTJxCdWsby8sGJy4sLOJp6er1E8
Q9Pvrnj3gtRpy9oMWQTgu5lGlwIzJKuay6fIrIvhvjMwyw9fo/E8gLSfi6aPtDCXx32Hq4tW55yP
mJCA47ghsuRJ5WmaPo0oRn7uZpzkM+tBabdBhYKMB7/J1YV6sb/iFSOrWUS2AcBtB5Fl6f4/qMOx
bH/PeqI5+AcRKDrQviaBH80bKNfhliMRRaFjDM08spBBthuLB46mRkVRrzfdW1IF/itNKA7DI3HO
RJVtwF2vbkoZEJiPb9Ggi90dbMgkY1JIFqtSB7sGPYurO15fRr5xLu2idz0G2iQsl4McuIPDeEAx
JLh69V8HbPYJFsC/XBhdVB1QsLJ5OY9FQMjRh20Nepi1s3pRa5oN/BblvRw+PC+7i/fnOTQ56xTk
ituP9+sssAumUvITlb1Lix3XYqgfY17tJ+TC56NmNvA1CJiK/mh5t6Gr/ixT9g4zQP1UG+zYoulK
ePVALvx+CU3Q9mywSwhWrpm5BEooDKKH+lMEqVqTM1I1eiAY4NNfeyjQqzu+UZuoHqnsDrH8qOJl
MH1opXbmEqw1czQhRCxezrVtM4FQxJu01POEYqsHU0MRDmu8hKpMTRYXc4HM8O/inoPZR2Vx/WqX
uaoqWS/G4ndt82+Pl6PtEA2wk7NroQkLN42nclCB1J3nLXagurgPhQ3qqeLq5TYVHackg37aQTxh
1VQZqV9ypKeCYpFePaypre1G4Ogxd0vCpllSDP6Nx6zc3sGB8vNZ8QfpuIxay/XsXsklTIqGgAAt
emHZsYsmAYHi0bxEWRvxu8TyiY5spFp6mSqbpPtJ8oKOzo/UCg/fyQ2mPbQWyjgvGcO13a0m5+2O
uFf+D8yTdx2MtDm4HyRrO4QYnW8phjC3VWv6WdUbxc6WsrWN1cAY6pG91QsVVJRDOTVfFcMOws28
g5YbRdUHQx25aqyY156hAjDZ0X31xuq6SyWvUtwsXo8rabamj6kgRGhHpb1rT6hH52qF9V7sF8WA
QwQQgKeWBovdTF4fdUVhaCRaf6udOcYzuer5qjHF6ymZllDnUf1k0FznlKQ/vOu1a7qHC2zE6gCB
mJHFjxWm6jzGRQgwd8f5Qvh3PDn56mAp7+NltEhSMdknBa1po39e44G1LrYSOMPOTJmZzyMovprp
jFAdsqZCj0jzpN3UcTv6DlGKyKREmtPrDiSIpSGfbvx9Fa/G06f+edF8mDye+qt/2NiPq4ctgUsx
TCwWVqRWR1TvGCEHzxyCw8lYCRqrFFxiNZJpIcMfPSqURzrFbuyppzIXwNwwX9wPHEoD850imoRI
5g2RZehyUJ53KeJXHif0APk888UjBJA7adCj7/HELUbHOUB8ONaJSPO7liVhc4E6B57JhDDDNkea
8NtjygALILxA2nxDexjRYpV6V8XTlOdoRthWps3RLnpqxKnLVs13adHkTY25NU07J15PpzFYJzSP
K7KWO84Rles2My+7tysAzrSBf8vwTvE6lZybIjWOLS9BZHpIWoq04xdOiDCDXe3u2m94wd7dNZlM
UmOBOrgh1t2n3QbhTMeMMGv6jPH6oOPGgcHWlej9g5PQRvbk7/ZKt0ilqq+xV1qDgjIOnngJPo9Y
JsvZMMS3ao0KJRJ4W28fYPlxof6NRldVQ8zQvwBtL9+a24pAkQaCZ2xo7cTl0cRM3jgsGpO5mIEl
GibYc0fYyp7KfTatYH9Cvcoy7R6tIDWIt+RdcMbjTYVS3m93pQqgoA+1H2Q3G/+TmFrns7RRQrSP
urbYycRjgOjy100J3KlUDTH82sz3cSgEo3QwFtm6YkpLABgffcX4W70yHQMiHw+PIZsv/77/wH/7
tBFNznyy/uDlAGWNxI+71akzCDR+H/SA/5pHT5JBaSpG0urnOHKhuN9PkPmLyvcq9reSpUfTtRbp
TGrszv61YIeiL3SPRbOV0mjliHzO39voM7qksCZD1QpyzSl09yJFSlbeMPZLXG3FruCM7OvSY0fd
um+63hP30jzp5+JKe0oejQV6d7CQjX2ZMXFmjGJKnmPA/fe5NU5zQwpdiSzuY+jSAVg1cyS0ZP5a
pI7PHBlwbxM5X161nFBDyLVA6YNHVIcx9XL3IEiJvOvMv13qpLsxK8b1sWZReW9MJmUF8QXi+UKv
Q4W1bW247kFhngDbRFa+NRlj5AFBKBsapRYXs0QrjkYVQ80+/wLUSwXP7+lMck7+2iAU2VIrrBZN
yuduE/TXxldiqBAyGF2kr7DFFy5CPv+gpdHyO2s1FqYno1FWL0dLRS2sWl+O52iAGrI+RWfqpEPo
UyA9hsZpjlKczFR8fMbmzgONidyIM2ahsDlm0GoWbn52RjbtJkA4emIpmb1QCcmeXoQ9Ezgb6pAG
AOifoe46NJggz7shqPcEPUHkVgUk5olGmbcCglqk3GAhzfQLf8wmW6dy07I838V0IfBY/4xGq4K7
Xr8aeO5Uu83wBR2ts+RHRzIKcNFjKXWu0yU6xZJsBqNKFEnxQfZzDUmn3C85ve+Y3xZJ7HHwWl8e
TiS2Zl4JOd6D8orVWcYGwjsWUN8ICPzhaXDPUVzsylJh7g4nVuFpdgOcomBu55aR8QildxOZzGWu
pp6Gqsjr2T6QGkZamjJnNX60GjLFBSa8B/bMa4+TahObSH8PH/8QHJmQUNUHe18d26SrPAt///2c
4sEc1Z/YOJ2n8EsqXli/kqJW6UpWQXUlL4BvalIgd8MPbw8C5rgzmzKwJasXOVUhJ2tn2Xb9g8wu
VYa0WDKVMgCY2TRQcagxC9w8C4doOq1QcFhM6/ybCNIhvb4ckWtOjzKqpOQ2mR7ekqlxIojDS1Jl
XTkgRKQvDm8szLzUaYRGWRAugQHNoar8eTEjKIkJV5DH22JsY01JI6YHT1wtpjlbNE83jApwdo2H
bOD1OEXvUbFEqd52hUpSVf8cWEQTdonNo51iNY02ROgrrpahH0LYbMMSHVvUVzy9+exy5ibtpbDk
IS2jSSSDjtbSm4MIuHFlpp28ymMUBTXPdWkzxtEaDOVOcHnGwLbbM47mEMN/oS3flJX3nOhHGNla
IZbdDpZXVJhxEcSfC7vrF5GJGYxSL8jmgoZfBsyO3Fa13+U02xcTAIey+1Z+o0USD6W9ObT5eYIv
bqOJ4079UMScoQjVuKn+Eprbj4LERvkhbk4KIo1YnQVuvF2egsO7aJ9laQ5WNdJ5TGAAKzqXpnXr
Ppc4W9nfXdLVmyOboTrZt9Nfqd0O3igJuXWtG0mitCvi3rNFMaNhDauk4oGmFbRvlFVBmzERf8HD
Dp1cGNhD6hHkc20dxplBlT0zH2gizPIoi/7Qvy4Jgts/+MQBfi0rc9ynQOR1WaFKj+ML0qR2n94k
TInIkI5Hj8bv2vFBYmvNjsQb+cPruQqHG38616a1cECRtK/paG93RxUr6JqnYl4WUCFf4RC6bGrm
3N1pBlYqSXPNXYC49Bwb6wvPWh/RXS0n3FHnBYPq2C3pN1F20I9ud/w3ny0EpxKdUTdidMfmEgNi
fbwD8SmTnREVIchYzeT7/IUvZlh8kTQon5NvY/hFXUGkCy78bWvwaKCaYbzKJXSlq0Z3GfZHkNWl
wTCfmh5MW5BBAn9/oUfs4hc24K0CPJEmDZ7tfcCBTadJleuWv/yZJ51p2tWzp/076U7AJWLdLGR0
++IaH5bELGo23zWaLE8LFPSXj8v5pNQQ64qXnKUkQVIdaQ64TG10aTJsQX+ju8aFnsriQZf25SQO
Zbt8FIhuBPT3+GbwclLehtGDExsT26aM+l//Z0G4n86yNW002IXX79nlltgRD3DfmbcdTvjhPdjp
IEsYthqAUXgz6q4uIerNaZoZ/9VCG7iUTZPT4PGCwC0yM4voTUy08q/2dZYp9wSPKSDh+ihyLTN5
S4dCxh/jGPVau6rPSII9f9UgrddkKYDqB4IfaAlKKra8BI7FYuWQXWcex01sKHSukN0yruqA/DKJ
aA7DlJwGdRDbnEsfRrn1n9C1Yj9S27l9cBfCQtcEos+AfVO3d2IDZbQ05FtpUtL2iNn1h3MJGeQK
+vKf8AiT/MAWJivurIQNsSCr/2OILcIPG/2qHtFIngqj3ObxKQdEj8q9HaawNL40hTx5vz70ifP4
5QY9lBmkYm+StfgyWyTwJKFXIK0YA643/VipEjkjCJRjPhdTETbkgi/AVja4zkIpA6JzG4Y1SI1p
tcBh1YyG4/Qvt2ffbgNTMN18z3gAvY43MMDiduCn4WBBEeXofKkcoluxnWRrYTh2nBOMGdnd15Is
9IEyUf1f2ZxUvIJ7lYhNohRSJeEiT7tnrz8Q7M1xxqzCcuItw/XuB4InGqjDchvNcziCHXOr2Fa+
Shf9WtNQRIKXAYIAZm4MisqUGXPKPXnREglS43F3x4rkUJ08myy1wLjpZX3FqS8b7WJ8oUzldoyC
Tw9lRu5j6G1RZqIUjIQq2j0R2s0WLBKLSEMB028LL0ZQ985I/z/4CtUAZ3SXlOXI4KgzmdTGvZrQ
6HUR725+SNbrhfnI0J/MAtJ2dfCigP6mxMoY93cVB+XHE+8AnIonQWau4PBQ7UzSb15VcO1UdfgE
QSYhcKffrowi5kHqppPQ8FuZrES1GIOnqoJ7mzHmPy4+xkG0PVsfygREzJMDZ5mOWZ7g5+cX16wA
zfAzPZe8gRcDNMMJGxNqV9696xHmfJo0Xik9oeqEvLJRaXvcjjCNAClcKZXC992X+2wHVspCnKDb
bYBO56bat+ndGma/uoyZwzt8vfRzphCe+Ty0WRnVEwOmPmBTBYe2PpyQaTPcJ7zU3EkxMsgM0FE5
e22t/VDC9oqsRMGcJy7/fOGwn0Zqfm5HxcWhFZsxrdBxoyAMEmYrpN2OQHq4EkuOSbaZe96n9mN0
Cw3k+MB1h+1Uoo1R1rpOWTA8sg0WlZAZaYb6EYgiGR3CuQfzlh/+45T5U3XR1h+62Oq5rSHKZjI+
ZheNiaeXiEhAc9TRDw5zmbKvkd1rJuyFUO5gSoiiuDzMmIAYCaS2Eg5jfKHwNcE2jhYgkKbpL5QA
M4j0DNhtrD2sRCU16in3y4xOJg0kndvk1BCU5fOmjnUdDlee1xGSFeR7qORvw2GqOwgVuMSMaZq8
yBIngD1wDsnrWtTjAKkKGm3mJGWklqFtMRlxGo8rewRPImy2Lj8Isf3KFhQs0qOVgd/+6Dnz9b27
IU4DgZwwSuFP6J4SbFCi2rCc/x9rs0BWwWkwisl4OJIIO9MYfLEHfybJouSMzW3LN1j3/TJDEgM+
Yt+oPOuY7KpFT30Zqh3E6i6w2Fs2SDmzvgqGSaNq9DAgIP3vMVNRD3+Z88/K81kKHM1E+ls0Nrbm
KzrZsSWw1E5sfogXxsXmIPPAeVOYcGw57PANImsVlDVBGQbeITPgHnTaS7FV0PIF3Ml3b/aS6LI1
hggLh11qQilI9PdgUPfvFBqd2f1WaIefnEIeKcZ0+1GuBv0HBSR4iFpFtBOISQqglet5kDWMD4Ny
N6Ioht2kD+gBITqJtToneACaM+WOSZxriZ1C9Q8dt+ZQb0eL6hpbRexPZ4wqdP+Wy0pvb5KTS4GH
V6mFviRmEtsWw4eCVml3E3SyTImNy61WU26FXC83Q/uTe5Msn1Q3ekF1q7/s9F8xX1Nb/roszs00
hynEi/abD0NA2f8x6ij/53Y2F8Ekszr9DVTbAkziY5LTF5w4zXxwgbKtvf+/e6qN0CiTsVZ9RWSR
NLjDD+Eb+R8ks4gq0cwMajhU9GUqQ/PRA1/xa4kHHPMgLkIRWw0w+0ExWik0mgCyHj+Y4d812ZAz
UIAaPHF2/x2A5YU4NBQUPKbxt3spmZn19+naK/GuWw2tR5zM438ON5h0RxBZ4gbCisCHq6CBhcO0
PXeog0n15p6FYIQeC8Ayss0umx95hHzoLsGCmZYnb7S+AqXspWZKYJB5mEoURgkcacRR820haiw2
zwVQUx2B0k5BVBpaB04v/PTCAdhD113AuUD/wCFxyEKblCzfFEbCFK2Y+Ya7l5adCfcjz0+R6KyI
LoqUdL2WwpJZjl+6/eEDz6bEIaDyGdi/w3yKytC456uy/TlkMRzWSy4++lGweRwAXE82Wq15aLOB
ORc5eh51LvpI1ze1MVMRcO4N5RBv6oNRwyQPO+HgPTARIlCd4xdB1GGmyxM92em+GEg6huBeIcgE
b20z11LBsCE142rKdyI+i3Kax1uHJdnPqzBC4zYyMv+j8EhktaWNhoXlCNGA9KUBrsoVqJwlZsSQ
FO+PfZMBpAV8lmdmYwZbaRYn1OUqrryCNi5ptCtPiicV+BSeAzTHkW7Mq7WpPwFUvfiR3tZZySUA
iozWur7d+GQyMcLhMv/dMV862OuSYXn2V/dd9feg5CQzhOkhF7pwah64mktvxxeU661UEjjITpxm
GonhDXUzmi6aYsUa7A8fW+DEW8VMVwliT8ZJhCXnS/pNQOy+LDFtyqPhEP9GC3RDt3+Pry9aozE8
H0t6tTpaGGXgZMhoavwvtH8EFfI2K6kA9u8oif44vyBxQLsm/r4QTGmk2MrBaNSCNw8AoHNdGCmw
pkFhHxugoK52qlrTwnqHJNw4CpuqfztFPHNfZyvj5osRcbRrdTYBC9hzf2+hvIdfChjBE9ImZTXi
gdowMluRnwdqPFp8QC2GudmqUXumMjC/faORmZoeEt/M89D/bsdl75y4nqN/2AkcsMFY3gjHoaBX
xVrRYzWLsMYFcw8VFlgH9qOcYWQcsDieDGGwlmk+iu4YHz3hskQg6Y1NU2yW+61tykalEyKYidYX
JRdC93vUmj2+6ThczfLoCaVqYzct161a4ZHUrtVDuboU+9l9XbmrjeC8Ac4IT4Dp1iFiMUeNMO9G
QV8GavQ9Nv0fc4ucyVV+oTbUeKQ2ZA+MpwUGY6Uaz+vTVY57dTTJT5ovInaI7G7iCa++YCoZkNvV
uZxd5O2jQr0l1W5Wyw9kGHBdMi2qa1S3y11S3YvOCCzUjfG+oiQ6DQZ3BnC3sULDNNsU69Zea+vI
JSx0ttSE7xKXCEq8I6WD6sGO+ElRfBeohBNnWvegvZQVQ3yE2NTiMId0RJSQ5wSzSdWZ147jsHTR
AnC1zHuMaoPXYc9h8BTEYj+XRqisT71CSFVUznOOOFQwgXyWEWZC7ZWk2IJeg3pJ1vnUULOlfMj/
/l9CGjDkJ+fDovHjz30f8rKnGFmz+j1Yy+wUN9UXkdkJ/XTU+G4ZscPsXpPV47+dPmBgeOJefiI7
0MgBEqHX5z9eieagjyMkWZdOawgtSlAltSqdu60SI/Qbkfrq2RBRRuyWKpNwqvzzBHsDnKaa2z4J
MIH0TNZvJuKjOxcLxc/0zzdcal/NRLJpv/jbJRjhlK06tHROCoex/5DrngSMA/VVG7hZ8VGcjv2C
LTtB5a/PcOKVkmPT6iMhRgOamsW9xIutwhlZRhDpRfYrAJw9AJ7nT3he0rHFnlY4NBQWYXVh2Sk6
cvyGNSeIoW92+Xc51rGBzKLXGVr6O66B+kxyGtdXRnsztuIx/ktAjjxv32l6nTZHt03aUYAzvodi
hdbykHPkbj1YqL9tH5JluBnbBOH1pqJLqsSt4RiPIr9eNZ0HaMHWxzKOzzq8WdoAFkr2f687W5DR
5FhY5TesjAZTlhBZ7t24tLmYOf4gKw6gki0auhGc27XjhX8w/nFJMkPOEoi+r3SdbnC0yQOxjJ+g
tQu7W5l7kB9Cmzjb6fNl11lFYMVQZoObqT5gz9fY1mMXjMc4wBSPiVpxNTmrM6xOvqC+SXdDVWwg
7wcwDwg5xfw0wsJpd5LYoPUyMqe82o1nTDiByWBdPp7K2tlJGFEGdFcVctpINNPZKm/nGOABMDiI
KpLJQpo71+wrQrsRM1jZv4SncShLdIn7JptFtjX/xmFbt07+9auejbzsJhEsLFkPFSclCSMRU+uD
OR3yLc1qFMS+hBEJ+rJFqPm249CSdvBxyteA24QbzHNK3yCCcQfeiuoMK2F5/AakRxe1rKWWyN8r
n7OVMpZYO8INm4L0Jp0zPrkOUrglw+Os5XV9b3wVeRlSTWgTJSaIlgKKpcKSQ4PqxJN4/n1ZwhG+
Lv9C3q2BABP8VKWM8rrRtG2WwP8ALPNJTPyB18qogq25qxqauQ5GRaj/D9JPMcjfHqIsz56kbbrd
vYNMWx1haftoEYxnijEGdOh6YSRIGkCPZw3QOEw/0S3vTLCy+MmYegcNyhyF+jPvUdswMNavbZn8
3KFBwmL3Ga6glp4OXoXURCO5H0lEa2IkPMY4ZTzYoX0aexAADHKCXCdAZ/nVJyb58Q1NMdOSX5a8
Yq9Cin/uXYI3OOQIEx/UGANtW8BKyKaE7XUons9mmtMZ3jzW8fjmwXV2j3f4yKCLHYzHKRgLOAdZ
QpASpkxn/ClRWPIz8xbpzdzLA00iDpRgbvce+PDYCUQALnbJUjSErk2vbABhOBKaYtDy/X+kHueI
9Ldw2BKFrS0c/n/VDj0y2+pIFJckEhwwtbUbB3uVjUCkPL2uMMcNhtbEfxyqp9dbh8dcJlihi4Ww
NWtj37GRz19RPgA9onIgpPZCXfPCYXOAtkDTlKyWb6xRn2so8l3mky/CDFlUogT7/2UALVFegRFz
UUrkKO0od+UvfJDNGZ9+4dQccwMQ9aA6l74LIkQ+38FbnwYuq2VGqC4HFUrpmuO8E0rZhsrNK9EV
6PJzf6PoOnXkRmqKSrYetkyRFHW7refFoRuSKv5nH1c+7dTJuATUmk9VSab2CKVMfw720YJcs8wt
epSKACaFC5UR3ONTMfFWVYNGUzXROVcBRY35PVo/yC96ir6SCP/oX3aAV3FTFDFkoKaP6Ha1fg9F
eO/orA14HDkpOakAXyfW2lz7xCG152AkaPK5zUkQ3biRcNCdAbW8Mwso2Sdgbe8hRjxKX9fdi6hu
q1uOE1s49Beuw15gMDnUF02M1HQ8W+q8oTySkx+0r1A9vzW/wW3atdOszwxNxL3ZPnSaASxUyvhA
xmmE7tkh0yNPb4AUaBuSy1/sfjmiVk5wXawCSNImfH+DJux3tQm4D5+4x9v1phmiuNmUhDjHOtZv
wD34DrJSuT6yAGifmnHMkqSvK7cTSUv+R9Ly47qD7ck0GghQRI8ANqob3+upl1K0V1TdlsECbpzZ
PgIc4mJqaSoT+cfBH66XjTMl+UHArp+2xYcFsjdSaZiyU57EDca4fI93pKfcgKM9T4uQx6XcSAe6
6EwyKMgrtYatVRyuL6qfdYUzOdhFHwqZfBT/KxBQ5sBacdKH13r2kNGPh4cKdVWiRiajFzaDoLEH
aFKq6j8H1Tr3+WkYG7WJAI68os2G3A5QICORc1gQhldpJQcV85aG+9C6hmwyRs2+gNdWYoVqn7Y7
H/91NEJRalXcF1M0kMUdzbtagwiw37tV+ZKrIozVo8G5vFdAVojKcWZtyvYPg5JU3v5hOvtG072x
xpmGfkSlvhJxQWBX4d+cxvab8EC7N005BDw2MzAyoDEVjb9DXaO4bCsLjQjie/adSHi7hH7pa0ah
IiporJFweID7kP7k+ZJNCUFcroCxGCoAnR0ThiryMUrSm8gpkjyEfyFh8lPhluTM6bhuaXCUqiLD
/cxMI2oaumDWuvstShfoDutwkMCfvGdeGqXLXfNOzgR3Z2UEv02RLA6dBq7X2UI4HIr0DUtZ6fqe
Pu9LJqbagANwcf/vJUHPrtv9xW5sIoIkEzouUzQHR+zcTz0VhF9iVQLjCnQIJoRmT1zmdN6MbGeS
jGzczDhbK1lMN9gHiyAIGBh0MZPvEoSONOan0YCzkP9fSmX8y0i3seg/MPCGPWVBz6YM/2uJisfd
Kur3iUSfOEt8tJLTOT4euNtXBm5UowS1ECB11h9hM4DfoKfai+kDN9wgWlaMYxj5erqB8sNzqkBq
DK72WVG3pe+sw6m7pTPls3BaFWB6+Ghryjlu1c1EUWpTmrjwSIw7vQBFb7KsABJVyd/URLOziwZg
xVhMHuN+IE0jqCytHMIRijyL3C/qWHXrbMzHSIBpRyiVY2Ao5SlPhpeb+tXkwQqvhbtPN2PvZmvE
2DBNp6LhUK3A4BS7J/JGDoqr+zMcS2ZMFBNd4n3H9MWDb2gGaGosF2LnwThLhy/K74BEFk1UpgVC
R4ZBhx2jIKhQxWHmZ7PcQ3LbKoz+SyhTpr8JU3CvwJcJbnm8afhSS8Jgil83QNS8OtfbRDc4J7Ri
4vFvlnIjVUDPnfhUS6LOyWslIamXvTsGPDT32dy0YR4xsM+XrfrBFd6ClrVoBkJYMKAl8hR8GbSk
D7onpuZp2azghn0LtMUL2vHmxykI8CPddSKmjOs4/VyoGjsrBXB+igol1Rc9Yg7S6tAWKpQFthLh
iPxJruvfUTvZQ/n4jsPMSCh/QxB+t1EfNmUVNAPXT9IJXHswcumaDGhNV6hN6pSTcg53VFZQfEV/
DsN/w19jZr+JgO8uOq7OpwLxXbpRUsoDnMxI5U/XY6l9I/3hdtD5HkUgmWRx6xi+7ZO3HYM4TOfM
wjL0rg73nuiLagd0fSjN5wLzzLI615OZPIiSVqgEbpHZpuabuOla26Lf1+rtVL/FkhcQt7EAkCUX
18wafO4C8l+iKSsfD3tDA095gtpc0Qi0kRTg2rNz3tEYPmmwWFHAxwunjCU/WFYRFDyy1uvpP2tE
oQlSA+dEYPJZiy/cBXogr+Mjv05Tz4rojjEJ0jVyHtq2qqBcsWh5dT8CuZoXTfub1gsZDfcMYD87
74dozFPVM4ZF3wM9WyKZa8PT37urOdWZkpjC7CPvZ6WmKH49XnXf3azKcjRYaheKJu5ijts9d/H3
5U4eB8ABfYr8QqlR10GyFAKsbNVDBCzePlcajjnSmuIqwHBnnfMTlmOCjrTNkUBvtMEbE9Ud9FLE
K/ogqThjSCkjfw5vqKIHo3bGaEVVgTdQ0uBRXeiF/ZIlWyLeidMIFZWRK9U8zpzOgU72h34VI1tH
3STVSE1XLpUdynWx1s7ZjtYKm6N8rPHjrMAMpXETLLFjQBuyhC9YS4Sv38hhwPtwvCrAokZRQBy2
UQv+sTffGXfFxe8QAdeo1lt8rAqI9fKGcjwdp5WwWf6kfmO6qP27KyJsPTrqd5mjuR/P+Kua+8z/
QWjw74dTuNj9RayQ5ZPhd0skaSArZTN7iOFPkUgNLKAz7NeC1My2zlxgvd/PofILBfpZFhoPP/kP
9y1AQUTCAVNl+d4rN9bEtPvoPkdpg/FTu+gw4PvQpkMMt+bSqfN9GEWHghJabNGfi6vMoxaAXnGE
oIOaXMHSJhJgPNOPcZ6nXs4tX2tDqn0zr9YrkrPf4MmyoTm3ulpihNpl9sbI6JVQfvDfHydbtJ3H
EKWd7Srh6yXuT7NX2ebk8/9c6z2Y4A62sQNhfxbWyp/NH70/lTSCW7bGn/xasZh8V3MwF8Psovem
LNGR0xVhpknAPVcHb2XgEmlw49VqucXHPKGZMr3/0JGGuDoh4gDwi2R7vQYTUWSEiNOI5lDpGLxq
1AOJatsaEqRPYz0CYnnKKYVAAZMEzGuDBJz7p1nW9Xh+CV9WhFyP9CJTFwJutwETL0sAgXaMRVYR
8sK4txXDCtNWD6/E9RX/Z8K0n028CzTWHagI1Fyv9oOS3kZW3x74KF0iK2TR1irp9wBJalGwa3n+
gySeoHmDHH99MCrEMbE1mFtX77F1GIWOAhYMzt4cAt7dl9WA+dC67cJDMooM5gDNK48HNCTYbz1a
7+BT805RN2eiuUoQxAAxu+PTFuseQTvPBAkkii6QZf955L7VQFHiq7CdAFfWuAnhIRt6RJDBWKzb
e2qPWrEz0ZbpZFxz469v+IqkpgybmZnQEIX3/UZiGrZu/TayOBaLxFTJS2+DrWUl4xIrKet7l3yF
mYOey0YhMpMyzwZgoRK1uFZi3aLwn9b1+zMW7D8GcepJ+RIphmIwdMLYnkOihlrjCitYDwA+Rrj+
D20hniib0vjbXMrXN7HpCYbcWG+xNLbqyXr61njaxyClPX9OZntnfkML+Cv3SbxxOHu6GhJWOS9r
Y1hg/amSUG1h3p4nvw/WnbjSbLOxZ+ej8Qqyu8+NLpP3cl4x7QOqk6OPGKetsIgNelGHZSzMC76o
ICQtM978JEE4V/I92o2NB5d1zromVgDkUADGrasscyZWCtBTSegJhqYj/2QmPHbwOyKNLZWe3jrK
zKEw4wjhD2du+PSF+ib/+uKuElPVdqlsNjT2uamv2czRK821g+lrzYtB2pBEc+/Hg6csAMumSF6X
cU1zCUPGeUIVFEoH/gg7rkzbmqJX43t+hnq9rD5dpifnbweC0lV6IzLUOS0/15yxAn5fideLQ6MM
jUEIC2sj0Q5o/aHV5xbcecFsiQaAZUP4+3m6s8xS4vMqnPBiiBSR6yDV7BQ/QwPIBdU9tKFwuGnI
zeNv/ug4apV+GCeKjA3MVJKgzt7xSyB4IGeduYGPCU+ADj/mT2XUhWPGR7YqI8W93b/4u7Z69Zz7
bqUx6BiUt02waSW+yrI1B+SL3FHCe8D4Wg3BISpkf316szxGtyuqYjAGdoH0ZYjqfqek5am+t3Om
1jW9oWpuQSqK7VZrGA+n6CuVaTC9IBuYL66OkkcmuKJKqtzpPc8ZeBJ1LWN4KbEYh/6CA186i6zR
07K+CUHuzlnciwC7OQG4ZOtnOKNS0Vj795Od9T8EPQCsh5nmk8WDG2mdfl7pkeQcRBhn9frpNxSL
aw8M1WyoXnUBxcmKT7FVQZNqAsei7Pi/MJvXZV7gdmw7wfdZh6BNwPD2XaBNEPcCemR+oIhoFxDJ
QnJfeCCPvckFcCa4nxvL7F+MnsvJS9npW6COq6T6aoDrYm07WehvdTBvQh9aaPHfC3Bsyu/B7iVI
Cv2Wy/USH4m+FzV2Lkc+sZUDTACXV5NCVJwzVOXzydhab3tvY+3oBgGyl0U6fHo1IZGZ3Y9LjqCw
r1lJzW3wa0E30rtm9j3Vo503dAxEp3CEP24GQRYTo9MJ3fIVKVgRoGiw8rmBpJZO5UsXZVTmAdGd
XunELVu8UdqkhPaXDSkYqHva1uQXTpN+mAJDSKadRpAuXtcFidJxOJET9vwaB9RwaCOOaY9+bGbk
IZOLRqsVsO8WI634q+MRyAO/fpIV4izbQT/iGAhGHw9HMxD2X1xEnwCQCmyC/9xE/c5TOPkUZWuJ
8xiCQqGn2fVQgYWVVrTK/BmgTJpkPv+7gcAyKZf1P0nLfDXwZ6X2wjHMl+5N+F9O9f4m6c0jhP1Y
6MY19yfnKT2xwsGd6zM1o/FM3qKfeIt5YhF0kx9yGDhpgZSzUqHJx+klW0aHvQYuIBT2xlEoyWJL
mr98LjVHalCZa2aG+DmJtLIz9BBNEdwr+ZH5sOZSi74GDvf298DHNYyZMhGShvdUc/QEfGpgBzC5
gFZZrrtOL7GH23Dvp5sJVuLAB6Dc5Uq/o/dc1Gqu8N7wR8/JxP+H0u61I9eahIwzas3B4D6h98ev
0bh/vxln2cku5fsZbVc0aLHnjjBh+JODSsPs0rSs+ydYuErwWKP85OyhLEk462PDCqoUQM4uANrK
wmIKrkh1i0hcYpFJ6qAA3UuQdqrr6AEMbIquwd7ayHlPVtKVNdS42JRmJseadcwoN8AHIzHjTIYn
sdhJ3ams2wOZxwFkxVLJcMy5zqe7Z5Jpky2TEpIA3Zp2Pe7QrDNKYabdhyg9Jf9iJtBmleSQm2iN
5CMkeRwTB8wzp1rEwxofkpKmffUvUt5ZnHLxbhv7UC/fUOTX7RchR1BQF6PE8Mk3fUbkn3VzZ7Ma
Tir1lCgg8EOt0knoj0MHMp/0IwOjGO0bpnHaOOLYk8ED5PRN8UtdZr7LyxMYO0w3RmQ0GnxXitsk
t0uJoHRsveLX+y+wakqgDC+fC8rI6FKeCzl2vuI0lX+CM6EZGbYYbyOrRU670psphyyIiFII4dYc
jQcDTNSDSuJmQ28x2UqKeYYMQs1abEPPUV8NOZPjovZyC9CpNFpb6LbEDn8oKIe9gZUJAtYq8BRj
OxZHS1EpC3qj9p1aMB50PY9bCC850+eV633+tygli0t5noDSETK+fRCSDTU/lVAk6vLjWM/a0lnr
L4S/CTT7hMJq/PLnuCIUQi/ScisgCyMd8Zgdbkbc7VPQ02zmxoV5DhoPK9/Ohxxc39c1ecTaECYl
SD8QHtHcFQ8BI1lvmk41RWY+XxmjohxW7V7RxaXDRWkFEt5ThlJb6ti7ffbQWRsY37XhEV6WBni8
jWmoZIpoQZN78Z6wB0UtawOV4uvSvxWMkBTi9zxStgEX2bU4ACT1wlxclCXEXcnf/ztiMifr9QFC
hDfZXmtjzw2pwyOJMagj2OAGPWaEha7lni3CR9eA6QCW96rnQ8BgcYLtuLJQjiB/2KczCC1lzQSM
w7Glh8XKMMESHYKHLHNaUX66h7L7BZflZjAHgcrLN/3KuO/kIngxqGGjWKf/ThmvJazEdIVIHNIP
qYi1iLYJjAVyQ5x+oLdj7+Eb/G6UvyU8ZSsQG7NvZZgD6eEvbgBYOH71/QM4UAA6JEx0HRkFALnt
3eKcbH9nG8ic2ruq3ZqWDEpuFas9fQl6mHkETEg1LWcXy1kV8wU6+QXALYLYJuigPxVecddFFXzp
wVtIusosZDrD7QWXn1pTlkizQCIxdb3Z4kNKXAyqN2MEuEsgsQxAbJ19WCC+M2WCjNCKd2/ZuUCL
9fa7fmvhL0MNKz5nYfeShJWO77KpiOmur2N2vHOyBUn82nD1ot/RMhHiPEStjH6+oQ9kurTPB+OU
S3OMT5Rx1Y+ehS6liVN656qv4SAq5MEjEYCbm+JaDvbRDFWMsEq+nVex+r8QOwjOfCliwunN+WZb
oshmvH49j7KyLvw86CY/+FnUbe8ZXQ7fvS2P6geoe45eRLI1vLSkJM4jxqCCRL1DGd+wjZG62csq
sIM2CWFh+n4/fyaWx67aOsPlIKYv6BlPsTa7M1phCl1RlkHwq+PX95JlJqZgnEmE7QzPAs0lGSxb
1kQP3i0XdIVtNz9TdzQHzOsWWtc9rKM8pVMjwRZi1JoZXyvxBWxbkarc/6vi3BQ+aMFRHZoiB5yc
3+DKA85pouwwNFxDHRwJhhvqwVLoUUwLwx1vfXlqHWPzW67aMKKw9S6bxx4vMPBruETIqjg0OGUb
15fcPcKtMArhUVe48NYG9BCf/y0NjCaX5rMgjtsaiEZ+oSJQmlBmL0Sz4MXZmSJVO2IAmyatPFLw
u2iLD8BabsOkgHobKEQ+PHREJQWaVmomLMYsSWibvdKRvODkaFWl2oEnuyM3BE/FCxZ+4EOe90mA
Dtj2wiHcxAu4OqtCtUSR5WW9pq06xwGQKuv0OReB7AGHS1+cs3bX5Rm5PL+iQsWs3EkLOhMJOkLr
I0rr3CTHs4sYkxOCqEJTclHqcZeCz1C390op1+FZrMeR3KguwpacPOAWywvjnJpIJ68yESu/t6R6
uh7fWRWylLfwY4p0DeHbUa0RlvpTLzepx+54qRgvYe7K+PLpKl1xt/pjyxDnEPhlRdBddFyoNnH6
t/0u3vWJkY+Bn7xCpcrPFqCwrOVfHTPTuspfGllFFuEC7r+GwTDdgNPTBWY92AggRfWef1+JACRJ
S0znoJRh0MqkwFqjyenT9FhT3qQeY32TCC9+RqBJYBqOdfbtDo02VlfauQEh97YzqkLCdo2DEUs2
OKumwWvTvPatxbJvV3PDmNNgospPeAKckHK/4Z88mnT/HyJthvrJZ03MIF/m8tJgGyEDYALVEdyv
n4fWZiXyuBqiYbjdrgF51hM4beWAqoa1dIxWa83OUqdqsUPpAFDoMLr87d0Gk/mOEni43A5qGKeJ
7ykglsWAr9KQNXkKNZptmFoB0qdWYnWk2aFUQSGrTI+OtcwBpM/JfMK3FtsTMEWem9SAK5aqk5pU
OjJlM+DW7w6WmZalslZh6JgfmytkcbAE929MJfWk46W+0JUFBUH/vL8GfkHindo1QEEYdTmspICb
q10+jBvyH1YaFBxO4BDKhTccexHUqJ8mzPAmp9vW4uampSmjOz6m66Jxb7JMJKVPuou2XnNvsuMS
dYayGoUr7Xs7YlF53Yfi5IEL/VSzqikvw/eZX4VMgtBTze4D2GvimetoOGdumx0buP03y9QDroqF
40Tdotnh71aqQL2ZfX8qFWMrNtG2fUm1gh3oK618zEzhq3IapoQ1jKlzrWOamjYw1L/MUYzZEAPX
OXxSCHT38tBMCFv0kKG6nbDZPSb3VGJgMadeIav33wALO0Kk+TuBCM1b6kCWyzHSlIDGxoBKFfxq
i0GROqUShJVqboWg4K2iHBygU3f9RYuwZ5dvOAHF3c66uaIREMOiHMlxA4pEn4RoSVJI4pRQJtLU
J7pPJXhiBHCXwRC2+YYjFxtCrQi+i04XY2Iwq6O+ghKbZFRKpeB8UsYGlG93Bgtreq4wfbjuYuFA
yVJ60Q3BTaqzuH8zEG4JxL2zXeO5RWHJ/OLkG9KDao/pD2KfNJ9M04vCSBGLWQG/k6SlcPI5WlM1
p9xmQX3/ezMy9dibh5Z7b3T8hVRmvHWVB4APe+pn82u0+/xGZ5GGyJWi/NzuiFivh0QcywzG/cfh
ux6hLCjQLrxoifW9b2X37GHl+aC1P59S0cwIIqqlumGZrcmOBhxZXCysRdVUHtZffsiFwC05Yacd
ooc9TM3CSfb5bPSrSoWsWnBYoWz6cYH99pqPxf22pdv5fpA5+snVz1J/r562C+j0iTJg6mHIS1oq
7um/1Aqm82nMHTLyjXaRA2t3kphL44fhPBd0VcO685T3dNexkB2190Z7SYKEENbanJv5qMMpSSTf
XhtlxB4gkWot3+t69TPIjpH393Tgywg7nSAU0LwtBLvqsnGKvxZ7pB3jbjwhsf/CrYxx/x35kP/W
uy8e1IA6fB/Mvv7TRUo1iXjPng9/zu+kdgbNTw9YwFcFqTtYWlQechmj5j2MzdZCbKvWen8aK1tN
y2sGIKq7xof9OOBCxlKWWvZeuPfYpDJLaqMm9GBWGXTMuSOcO2IGjOXd6n1PmsPSlmYSW5bL0iDg
WGtWc1oaaUsKMk7ADD/UftITmWz8zaLmNlPxuuNR4SqMZTJFQcDf2Zqh360nDyvrt1uFk4gWjSJY
N+y/dMdrhzcdRAHXaHohwZAVHbKGY1oC0OvCi4H0I+Mr0czIBy+qgGWmfvx6u8NpLEZhrpwLc9wI
8bDMk1HQYSpScNFD2gurip8M1tgdcvausN5yioIup5f0J53kCk/GX8e0PUvPi9bkSQojzWs/X8yt
eVsTniSRZ8c/Ie9c+qqt7Eme8CIlbulRsimp/tos6FZMip9D/m8Lt917Vi6EZMsDuXnOAOp+wca8
KZ9Vi4J5AMOtvvOOiNV6/kFR6DLBURn0Hq2pWILS+LqJ87OCWpScEfximasVpP7lGq4CrmZZNwU1
+BmhVFE50js77BA4GPiGxbhMb+aG8+EJtUF5A3LkWy0S+6YG8HpoHgFvbMo18uo2WyFsYAVx9JOT
j8BSoPjfL6FyRiMAum0yhi2SNM3bXV4OW27Oiw4zWZ0qVE3bVVahmNEyT4ZWMGdiNWAifuY+PA5r
HEY3ySPGIFn75tQVcQPO1paggaLgWbhDYOCZ+OoklWWKAybqNs0d6oNgHy5HoXbZeGRr8DwOOndx
rkhpaNhyGIGztPH4XCEtnz5ITO9EStzy2VQs+yji5kbc6l5ApSS5WCCr5Yw8MdTrNpKf4Xb//5fx
Wv8dlt5oZRuDLhSGs7MEQJY8/JOTpoSzDWqI6Z7krwuW8tWZX9J6qw24vPkMPAWgG2WVyo/qr5Kx
5eDPO+PYSgxJfzChIX+0DT7kVcPu0rYW309h5ls02OU+JqM66eC4LM05fE2b4JE5so3Kr+5tDs95
aH7OqTgt29Z6aGcHJcurpcf2jDXwmlNCP6kH880XDjp+4NU9SxPbJ2EmkOhkhgVYiCXGPfU8Mr6M
of+3kPHZc7/9j1TxwolzJL8aigBcuWCt4ItVQIDO8x1YJtmYJ6CWNS5+FiZI5eR0XwqAL2nuUl91
80VYdAvP8f5fbeuX/VwlpiEecMk08wN8bw4uR3TYoPoWb7uf/eQy4GQPOPJEy4L9jUv8PyWw+EX2
maPPDzrPhrmElpJepBlhtD3nIDAt2bOyXbd7UW3auy114htTHh8sRT266VaD2IMjwv0Nb5xxVvLi
Iz9bfYn89Cw9S+67H4QW6uV7aegz3wXqLuq8bXysRqTKBYYM96YCnDNqVTMD0vhNbyc4C6kxVVwE
uIlt3vz7K+Fc5hgrlsQT/BbtwoBZN00zvlPq5TQDWyvYZ7phgnULgCp/hJb8H93fTu4ea4wvWyef
Vom0S/1QYS2P5w7qvQZWnXG7t0fQAjHn8H/+e7cwVsbSAuCxN38BhSOFUWy7TITPus/+nkwG+M2p
2EPYEEqw0/mreEmrIGziZ2TRyb4JavWR7emBs5RTE7eUPkSJ0qCmTy5yaDaZvi5VmqsAtJ5SzpzQ
QgQvwK14t99R/uJykV4CmLpKwohFx6ejHNhDFcdk6goTJs98680ulhOLjGMTR0+rpmun2tMUPvYq
BTySF915iDjwwli3m4+pOSg4Sh5+ahkXGXhX6c0d2RKIdM/BzY1aIzpx2e1BR+iqLlnqGFagKgmW
XZFxY/O/9iiYgl9VekDG4pKAXt/TWfWyPjAzLgCv18CQQX6lVvvT2HD83IWqb+Kszr3rzuJcDRuz
bF7PqP29+jJjL+8DofaP3b6u+x82DU6Om9pU0aIqvD0hKEBueGLziVvcrLEBcwajCiLdz74fX5aW
fd6C5YrfoP9MH7uXp0Ey56QH+yym7J61m2pB5LsONHIZFQLTsKMLbFHcVnK9r/9bIE65H11u2VT1
64vJo4jwYJJCXxY4cAFsf7DZ67gkaEfP6X2uPrHWsO/SwIFp8XWjnHcYpjrqF1w06KfJCnnPVZDy
0qKNiq2Mkcnk93urWfzjxx27sLjmvw8sjPcTxj8LhqGJNcC3VoH/kpTY/mhbXjMka6LnZSEhRhkw
8ypN74RccrFGFCH/gJfBVVbiUS9GmJKK5XVnNC6WShz/zBw9rKd7GzTQN7OvVhP+RlGTUnOMsUhA
8EKV5mj0u4ky0ds+xS5W+hrpM9L6tWZuZ1ICwe0lAHdB9Ry5ZTe83+iud2qPIwCjJqpPiCPHDToZ
5w8X3rz7G6Z11PY5fsDJJFyxRS5/XM0ZERnVKj+miBM595ImBHzyC3fO6Sy54BT1di+3QojuSRUQ
mPD2XzHmUJucZHl+wgoACVsV1V5OLAWwvv1E7qzwhjSb9lbhLMQRcvX6HVYX2JuHyyMxFRkdLO+N
cJWc9Rfe/f0IpVy9IYLMA9r9crHzK02XcEdT1bNWbH5ks3/cjHpcNzJvUttckkJVtHft9UndSEY7
LzY0SaYDtGWYnvZRbijfuk9eo3ZZ7cWuMpHYgE3nFKwaERZHMs5Jl74CoG23NY6GGGvDhsiK784T
aXjT/Hy5GhiSOaSuWWNa2gEcBQ96jGV+bLyKVCqU3H5ZyeRzaygA/kvYsW/vFASLJGYbL0HW1oxb
ksJUGt+0iINiajemQ/+cBRSYN965GZFgsZq5SmZYoD1UUP30RsXSCMmKDcbp8w42DOI/jaHsIz83
ZU64mdCOmPJSttni/dYcNQg8/w39HLXa5Bt41WMN8lSjTxinyV/EdISzxWXKxtYSzlwcSTXP6Tll
2Xy0VCBv+bLqSi+S7ucsvUCgXugB2l0IY3XP3G3x4hmmMAeLdberfJieXxuczThcxBlBqa4atfBC
0wKVOuTSbF1+P2sSSsTTdjXScfl/ZW9I0/k0/HgFZG47pkicUX9L04XTG+vwC+D3IGGLmlcR+HD3
Y4Guy3HxOmMAPppnOowZ6ny8Zxw82pbrVdYti8I556E+mZTckoXwTM2TYeGeHU8td7gvafQ3WlTN
8mVw2P8bKDVpkm8uBWeTQgB7D411bCep/UweA2PjWtVHKTl29YwhxpgsdlojMRpVKPva5nqUJ7ee
WW7TuRhs1PlYNcQb/EM4HzuHdN/oufZ350E477T1YuF/MrcLVPx//kXvO/ENTtPafNH+DGe0oZ2y
G3oiWzWYfkM/k1I47AWuCjbacMFGKjkiKkiIw67IRM+YLDHxBuP5BQ7pVT0EKz7l4o7LEwQaKIK0
7iJWe5r6iTnU36TWkp1p0jpMA0Ved92ctz6dTqOEuAYEoTbQGWMMX8rukS2qHJiGXjrgSb+RTBgF
m4AokAnt8avWMQpywiQtuuBgDA5wg+UCpB4IfPklZWbOStGRMB5nqmy1XNmu3FxbOHQUvDog4ABW
V7Ms4GJ5RFu/4Di/4bJ1fp0pdRmYrjbaVcdiZXWkFkRwHBLCRFaAiW1daXNQqw1VNMxB1AKrMFk1
10M8+IZxw3DllFsSTtup7vzttHUZpAJ0ldzmlgckWhKBuo+WYg10/qvvkb9mnwTsD3/3WytYmQWI
9RaHAEnHP3mK007d+6/2hNglh53fw6fLyXQL/awT+2oiOiCerYl8pcs5r5dtUjEi7CkxXVfhN9xJ
nmyI9d2nTdLMcu/F0pHCfY/xkuY292A0ODc9U5HqewLTmQCqxziYKK0GR/DuJawpPH6qMKFlTtrf
xQw3XcxAHv9riQXLjgSBmju3e7GPhbF+BRW/hctpdDyOPsBh0Tr+47lkxnqoZZ2ntodIUTuwnWVi
RzyprMI9PpWHc1JMrVNt4PJSYmMpSNwrL4yOyT3s2fH2izdJxeomgUCgWTqoEAnzTZQazphK6Cp/
UG9bz1whfPmgUzHpCnDKjifB4FSAPSeQMJYWMkXmt60qXdU+QXMQ5OMyYIu1AhdIYRuTPmibMH9C
HXg/aSHbJCut0GVW/1aKSR3tK59SwDrxePw2oH5Q40lPHkxMJtFiIZAhINktoONVO4+7+e8Svorr
hrmaIkRfwB92JAXWYwRf5qUWpg0GJv0EalUPlAIamxhHgjl5zRvIoePlH1pTVA+Ko0mTWZ1SKPRm
PZW78bYPT9EHjwuVF+cJD+DiEk+klMDgtLXxo5DP1cYGoGR7AQVbl74nuPYJ/X3aA8jR4Ma1XN36
NKHhhpxm+LX1p1YXKNVK2gdhfeYBonbrmu8XWWHUuwNYex0piqmljRZbl9PjpXiet3R6QRBW/qnu
mJy4jS8QAnqy8y8/GYO3KSjwqCA/dU2ZjPUzziZ09WVX7yVJ2YvTi8EgE0frVJikhiWIbcM8y0UT
GKMrDVoVZu0mZvNoP4fOTS/dh3NFHoeJeWf4kLXzdMFUlVTXyS2Uv9cR1MurkJCk1PQjwJvxFZ3i
RWPY5LyPBQW7hXD/ZSmguO4f2Mdxt7JQGe3Uh3jekE9cBv+mBI28hZ39i1Nhw66kkPJrYg1oHb6j
VnowTcVnBWHqmrlB53CREHYPgUdyKpEBhjV3bg70hfkpbsEpFmqf9RO2+Zl110TDbqDamwzDUQNA
Rh47k+vFsuqc0h1JCo6okAHZfwLA1ecPdUsYZmff1WJasbdwEgpkvuJquaiZ+9LhJiGR/TSJfNrV
9b7XMwXCwQnAaiisRU4e7/57zvLl3AvIYqEO7Agp64oS/HUkJNoaxledmGHc/JGtTrEujB+FVBqj
kf97J1sEzFi6CyOABlUyBGvm43o2rvavkNTsnD8CmgCIPICJ+/PKC/pB0mRS2DsN9/s2eNXbrqd2
O8uq8WvxmJmpc2KZuhKyUIlOeVSTSm+5leeoD5KnNDHBRmSYQAqQZdzZGkXWm5HuVB2vneTsr6cj
lUhfwv4SzNY3EJpnRy+bW6M+CcQq+UlYdQ1N1aXYaEolO3366yJMnLK+QN9otHNCGljAMCW3AQU4
NHvQUQHC8r6RGZJFW8UPZ2TvYs3tidTDR+XVpGKS2S0AhoNrCfRmxmvO1/XSKjcrSqtqVIPfH3sS
J4POvCoDso3WfNzRUP2Ww7s21gu8FvDhB1YInXfNSPYT5xgjwtR7Dllva/E6NV3Keo4vlhOxRnke
/UEdrsE7cn2Jx2LUfIn7zP0ghSDx6efYW0bHS8+IqK74UkTKpl724xqV/gixVMEUOjRFxiAYYXF/
GdackWuEBOnJ2phXYWbnoww8M6arVDwegFFoukCg3zbVfRJLw9ieLGIjCpMGQcbp5P7TVcsqwPsF
5/ms4q9qs7tb3nO0eonjXVgSzKumYBO9Kbkm71rb63JFrQ4EaRdjPcQP05PJy0sHr9LziorKg8GF
eSB+wkO4MjqwUUpmwcOmW4TZo4DDYQpjTJrT0WW3zmAdWlgQscwrFoVKzhQ9EUBvbAosLi1S4Vy3
1WDxZC608JLwh/FB3nHlX8rRvbiev9ysLjNXGR5dr89EWakxAN+MnOFsBgVVcWmLyqrjBpK6vl1M
el9jniaqyhFYPvIvoqq6c28TvujR42MdkY21AWML8c088vYkRg9ZIeaSwyZ8hh9dHOrbdipE/Zgv
3KQqOQy+oqKV61QEZgmqGGfZsB07krWD2LcsZkRtyS4Na0j0Sn/w0k38lpFJ8TJ0txtbysMr53TW
PD8iPAA/XK2vd+h8zMLODZny4R5gdvJKxLjFTUmw6ZQETIsYJjI+ykoEAGfMMJ6c2b+T04FOzpbm
Y8S/zQQzwbJPFssDULe6F7LA1z9CQWjF9cNZu6Qzt7RuM4gPApRTfoHXIGOf2ZzFhZBcGgb9KtBL
Jjw9GaBGEWvvIvr2Nu0dq8zQDN1N/9jcBPlJh1I3mcC+tfrw2pkHENPF1KPfaLmC9+SY8FB3z/H0
sALSepVsOtGsKgr4/k9S96fncHYOctCAFADR2uNBlGm+jxOvpODfhPjsff1Y/1FBMujwfifwd2FJ
KFrEd4mFFJyHQSY95vf21SyfNkzz6BUOCZ9pXX7R69S/XIpNCaH4OWg/wvq9ECfRbv2UK8Uwd3Zz
cAE27Dvv/EY6V6+tSiA2yygJM2GIjih/PsRKUB4vUNQJ3yjcbVpztt+HszhmabXhJpqLY96LJYuA
cpMKmJbJ9FK9Vnnj7bNVMHVgkZJ31sox70oPPslSTXOkzlFQ9pvUqtCtSvDLexgT+CMXsJuIZSLf
yBL0x/c8j6KILTM8ppkwgBljUffzucy39jrxxQGz6ibsV+AJ341DEKGCP4Ud9aSHissz47XDbVSE
zFZT1kM4jR5tIIznEz8Ly8NkYNtf4MVswnD633I52hLhnwZkOH2B7Iu5py+V7Du71fGplboYrQX8
heSo2ICUG7Hgm3lkbk52qhx5LNZueJUXMlk4OUKG/5bdPJjukFKm7esMmsWsQelJWir7jwar/3Qr
RPq5MHpntYaBJFtkM/S5MkuyHZhxFpK41rPRM+Oh9Sg2c9UQ/dJ5RHc9AQE7TASmcUVfZLkdmxgx
uKgKI9Cz6xp+zaXEXwe0/GTDhwH6qJcpY2qrI09uuImsVuJXpPsu4gzbR1lFUJ6uc/uRH+pafa8/
Ec0YUKBchwpSv5u/Gz4I/SnjEdWfO8tHmNabkAQggx/XR1zLMG6X9VN2ERcKaqHbVrvpkLrA4CnA
mKsZ4T4HBu97srhL58cGlrAazN3nQAujalPuH3Qu9JU6LbdJWu3j+ehUe20FEAFEa6qITFf22sP9
28ml0tmnvDw04tf/daD+W60jr2hj+r5i5tRvTX5aeMk/AuuPJkvCKVsVuUO1BvkESDR9srZoMawf
pp67QUGQ5GZBxCP4+hAsAllmXB5ulvwZ6J+mgNPPXfbdly9iEE2sonEXMxkFTYaEzNAKk1v33jZD
oOM179XibreW5CAjDo6cdvveYAucUJ13ktBRggw3e+MTlCdpX6QkR4FaNlBqirY9mv6iXEdZ7wWI
XN/EroelK16xW3nygpXsB9P8AMGP3j2uxVq+nS3KsuNV6lhtLsfsfHJfqlZDoh2i3S4IlQujfaGI
QqgnTPSRC77mkCkrIXlxBEErQ34tsConW/yMCb5p4pO6PzuDqA/WHUSeQ2HS8VMrfjcEiOYuF36T
Jd/lm80vvaGPSjRqkUO4QaCLz6Gulv+SvNYtWcxp7nPBYOIgGUNA8AIqDDNDwvDyFt/DTEdP0nAU
4X9pnj3+GxFf0Wax31dMW/SEdOYGM5T0apAJtl3v8nXHf22vZPjWA+FgGUN519cQovUG+Hu75yJH
MZic8JkM806OtKDAJSMsX0TLOXG+WlxDSoyW1l5FnBHHSGMGSgPvybuFnwOwxd1hVXBjV+EiDwKG
xd/82IryAfIu5unLlY+StY14LXWKcOpg96w3EWXQsSSYSSdnPts82Pc/3cCqCJ6TnBo9TjQbVjjo
paF2xOIO/ggBL/KNC4QW1C/QFkHzTkx4vm0sjwKvPrf8lb4H+mBE2TIjYN+MSa7MQgLV2iehYvRm
q133kfvl+671BaqiRbhpCkxzxdkjMfP8bX0F36wwtcV/JEZSEZhqV7sbP02TTVW8Fara7YJi/nCZ
Ydhe1PfXMUH67UVVYqwif3jzBMh3lp26pMiyhCL5BSL5C9+NMEU2TMaM8QyP9MnXtxnYGP6usCGO
/+nRK7568/nUyBvhCdRRqu00MwMy/somo0++sfGkQHWmi1r12p+YNQ8if5pyq2VuegMFafQON0KG
GS20Qi8FLpP/5nKvGtc3iakMVbL2GV7KjjpDbwj3cIKcUJuJkV04p7s11DH8ZVn2y8SWHkY0XHe8
XIeu0+xfFRKo6mWj12VUS3OR6EcsoAq2wb0SFeHGD1CSVyMs8vxUaI3cCo+wUEci1tcciUc0llLK
GCyl+pLAg5AzA4u6Y37ct9xTdkz2iqcVb8PO9FB5DwIsoLh5FzIXduz2ByaY4tgq0zSo6faXk2sX
E4uK9mArK6C4GjgW2UudeAi6/RY9DFKogjmDCiv+EEMSud0nGhtrbLkBP6du3Qi4oFGh8pkn1OYJ
Kar2Wme3KZvqVbVdEGUiTeEKRylbNBMVM3+dgM16/qSu1GSy5BH+n/MB9aNeAtOz5YF1ucmKQ8Ha
uuFa/AsaVwnetnc8hxLYeWp0gNRx1Hm61X4JAkisPZxQLKO7c072YpbzN3TBWQYGhN+GTteDa4vO
G+LvhuUI/HLfhOyLyqw0UAStsfNQBznsO/5Z0QwyNiBlZu31wj7ga8auvIFn6afeFqAPtO6rSqOB
i5zx2ad6QS0WIXJCyArnMa3PzuKfguPFeJZ6mfXw3IMelgL1d09VNG4mKENsTWsuKPhwhVeN0zM8
NHqro4vJQMcoG3bySWFjrbRw6F9hUVtSxMhYaRhhIVlx46D1Nrav+GUXYYFRlh9946JbaMnXiid7
My572WwxElJ+vFAito3l3g8yeXZWLNYiqGXntLTI3pBFtzYkmRNzS7uuoNid77zmsD6Po7gsxv7r
kSjBzMydC386cDryg3SzUH5GlSYgXVoGGlni1jCInObqB2pQ+IMC/0PoBi4VOhmaqSoZAh4jcVOP
xsV/MbEDe9AwwthMyOsaxgJTxB3EXa5sPhTrogrZaADC3cSqEoxiHJt/KYn0KfBuPAeyVagDK2IM
yWcaSeYlZ1RGVG8/HGdXsN1teKBCkA41I3obxcA/qwmA/xiarUMPd4MgqgZ/AhaaEh4IxEVS9e9+
Ee/bOIKYiHnLQUiWBs9UKs6dd0Ofj4nDrf+h5UEFYawKFjxC67znUXsU8C22XKk6hGRfK95W++Oi
YhXADeQrKQc60tF7JpQMKhKOK2u/l6XZYdoxSBFivYA1QheqFV31eXlqxq88N2ytiuWk3dbNlahW
1Th2SbkKiu79TfP5BA+nvRMAqRNFvV/Tf6Hsp2n6nzwSFj36bR7CVb6IlFi2WeAsx+auKT9mHvTx
hSwwllFBk5PtQdnKPZy/4/MVzt9Ka1ZIj1dDOfcVioEIRbYheqR1+dYghdD+ErgRqnCJsdshdHSL
Fs5vEsCvj0nhXjS2gFnqN2OQFsz32tNIdHRbi1H8CQB2c0lzgYUzAElh8rxtUs6Tipwq8isjuecy
bFuCCOqS8M42rq6p8TIKEEB6sW1dZkN0wKAxmE8JKNNNyzO+lpR8UtiHinbS33IzCauqZkJuc35m
t714utO/N8aGj99dqyCoOLnk9jF5DOfgSHIj69aeOh1VQ8++804YXJj6QOrzpcSyORauNXbs/FLT
gUSYtTaR269GwjV//ZUM6kIA4ZKl9jD2W79RRAFP8sLm18IL2/mLw8jDYDoMWxvq6md5OWBXVb4o
RWSgPtWrqDndHhFXRcjoasELZw1LhKhM/LXaVMYkiTeZdgtX6wzAS/OpFmrlcKe1y4c0rm4Hl4UP
nJZDQJzHjMSNAV7k4ud1qC4g5I2vXevsdo7l5aZoWQsYmwFiRiQ+5nKCVkndRgQTlQfBQ9y1DEzx
UzBRCMBdBVBJqiTx8M/mumidAwB0D3QsxHfw1Q+/2eA1Oh4yFNEymNFb95066AKySZW07mZvztXu
dqY7omM78k1nZONTJEmeIUFow/cRw1MrSrFG2fm1Bw1USaub4xosnATkhzMsXGVwmbgK+SIOnYca
2EpPaRjRZBEyPTc0tp3UPwgmS0w+PNPcfevfXMbT/SIxhwM8JHSAkxHupawNKYdSJDlP0rPGc0aj
b2EZI6IJGOMr7KTdaurI+ISGbPFGYfh8Roe/fjqgppmyATLKbXmAbi4h1p76obpYcmyy2xIiLms+
9B69cJPG79hUwH4TUJVNrDho2Q49PvSU2qQTrfPegTUa2uUZgLGkYm/Ax5ZCCQqOiJrJx0jP6bIV
oqVyz18NvTwOSI7Dl2KVkQyAxuI2L+pl21mmydU0GDZ5p03uUUzpB+h3DLkhiMqHD3Vq0CVcRcRQ
CiJHlpaEGFVqQl2giEaGzDkStXYcvdwCTcaGG/BdrnGWwsn2satRzxA6FXLqEBjyBZv7fc6mAkJO
h3MNYBfxgUZah/+u2fc6iXtcCpI3lCdp9SqpwFawhzMzYi0D4/q0byIp1thUbkwVoYC8dPO9yMBH
FjWb8NUnUBDsgUDn6HPkEAEyT4wOTnjz1VHSOs8MCKgBnqS+nLMtbdLmoHYKtv0RyVCg1vVuSe3R
cruE6vbBC20wDBtGBkgqr3/pUbnMPyJHzhdev4tNVvjpS2oC7tN+OoTflJXreP+FJWHpxBYd0WsD
uh+0FDQJJWoVGmKVkyHpMUn/IwifPGmANExtCENBBFY9vvvPuA+Lcmkg01Mtb1QGMLHsSoY98ByO
GdAzabwERAW9xB6bbLLiN+zj4Q0ax5+DMyGZvaGV97dkXxENUic/3cMgIkVLlgMk/AeG/7HMsBhl
+ocRFCH5bV7ZCXITHwf7SecsW7vDnmKOI7iODUexErQWhXTSPHcpuB7tG8XxwSDmFN6WNhbpyWaz
w8e1wbr37p+Gycksp2BlR5ujdM2IEdz6PrL+3KS+pgKp86lz9WgxDldO0VpVJPt7sI7/fgYEv6sB
BMXdrDBOBI3SMUxzRMc1xygp251BeYB/PQZh9VOs8T/ka3E5g+uipShF6Y7WWdY6R8L0dwSHC1BR
CD0E+NGfvzthZYolA6k26p8srEDPdHCGf1SwkWEm6P2tgkKQqcB4OYdlUf5djZ8gki1SWmtOgXL1
DEFAmCWOKEXqsqVsuLuyB0I7bzDMhxDQJL9mAP8X2XQe9h/Y9xTIf9mvi7lGwr72tcnwJFhFBRwk
ApYWYubMCnnwYZvGaS1zT2+4d3ulVfFTnq74A2/e2ReIlFmof2u5XLcwCCh+vyyyG773pXO+QEmv
eLz8sqT7WdW5CYX7Mk0XtegHtmY5v3QHIQQ+LlUkW1pi48WlEhnzkqRNaO/0+tZvmyij+UDpiAZ7
gAd5Fk9TnihC2qpnID9bpDt92Nn0qjPjcXoJDWt2mxgMacc1EZWhjNlWBY2vgkqdhjbj3SBmPKcx
rdJhe/ZuieCeOxOpf0ZQVdWGFTxZW+SYgeiPXF0jaam5Y8g0cNcgph9qOHdUfs9NBYXYvAYpzf9E
Nwi3FuZnNd2eN+OiUs504iO246lCmnJP8Y1rpdpFK0UD3iudIg08a1X1OttiM3d683Lt8SpNJetv
Afd20bO/F9uUfiye/sKDHJVOGeuSqwh3CNZtBiSXyhuolRKf0ykqvEJ/MxnmhOW+WJUwNzuoxT+m
lKlU75m/crPo5y7NI1MjtsTmwTqGb4qlpp3TQ/1vwhfxoZKpu1wSaQxzVqGncSnerzEQT4/5G8DC
4NKcQqF2oxUbGasE7NdFxhaNnYEzP/2Q2Oaoq95/Dquj6GRuMe8YGcqnbxb/rjOLITxQ0kntMqH3
x+17x+jF0Vr3hHtyjPO1VR3WKj37BszUGsHaWidETk1ylqc9CBSIzSHTrgrC5Q8beoqDdDk4P5YC
wWAsAEh3UAL/UKsvC4OqKHBn1bCjtUnFznD0hRGRU+7+ROTkM84MjDRNhIpCvW3jgE72pLsHzf2a
rmMxub3DdvNKPH9P6ksi+7eVE9LRShQnXpGiKrYLhEJLl1LIeAngk9UpvvMCUxhSUaXNMk/O0Vdx
36eAQmDUIjKbLUwy3aB4ctcRF4Nh11OceRf3Z6NTEIqdfU0ASmkJ2ZCohh7FWb+ekvCHUr7F0aZ5
56KQtRyiEBAywuBPVsFm6oFb2qpxw1DPhQ/XnrHHdVju2fo2S5ZuhLO78d5X++N1T4lU80cxmWPb
w8q8AW248NWYPBo5kS/8JWdUgNQsbAr03isBwMAzL5u0a5EXa+8QWRpRPYIdk5KHvLkbfCBZiWZk
rv3TVpVcbMP6oVF/eWI4fHhkk43JiiACMl5ImktTMwcUhrU8uzDLt7g6koz9JNGYA5chx2+eKr19
tiQjQ/yxQAsOYQFW9mtjTyW7PaQ2mM2ve7sfqLFlPziR48KoAtYObgOTErMMNowbwHnSw5qTSn4h
lMJtbR656AJahEZ6Smmzx3oBp5Zc8QtFvPgorAEsFm7BNF1r/XRg9LFXjiI14qPJisORifsFzwhS
PgoAEzlSHmXy4eDa0wREJIKNJMotm+oAo7mZI91qVkAOc7Y9XK/09EtYT06DBKT307O11gMoHP61
aKEM3sSiSb27iJwxEfeMrAL73ZQFvyqi47XOX2DLuVeHOwAsK2peE394he46fYq66tjZOHP9YcmU
/VtQB/mwu7mNN+AjiERDlYgO88/NwXDAkQ27YD0OL6nbfpavmGugByuM5U9BPCrdsJLkj8mWXNn/
KYRdj7W1Qh+hXHn4Iq8PH7a5BH42NRNUk8muaEp6u9fXHGrW0mleDfswlgZGNy/NbuXe9O59uBrW
fjXxkWt75W5/r2buXKTUY0n9dQDsPMHm7RNpCqAn/t5KrhbKwUlbdocX5Ghxb+9MrmaO9WbO+KR6
+/xFoQN/2oJryWNk/F5KottB+bX+dEMgjvvAIjE807pxnngzVzNfGroA6wd4q82qFoaR/QzdLGgG
hD37CRwrPQHfRRCqMjU3KMC4YBC7q8+WkwUbdt7D7t/8Ggf/QbDIkv+VajJpipIJ58wZkSTBlALs
Nc40VdihzXQxo6g/zfaYRTUvqRB9H290K8A/XClEHr+J+P3c/sMwk6JAAwy4JS8jA7Cef/Wq1f7q
uQUriQ+iOoOnRfpXlv1fT0femGK1gFL1yKwzq+oBz1SYESJWA+bWEkGvZ7nijsf449mUiVL4MQ9x
d9tXGEfsg54u5cWjuifNxZ1Lbtt2TdMFLhAuAhFmbH1aXepb7MoaFhWfMU6GxKrQhHZhgfEdHSsu
HE2EHuPsYUYrkWueUq6K58iBddz6bOTl5kLLoQQk1vAnj3OatiMr+b4UzllHu89WXRMXRLEy32fi
oQza+syfGJBbSNlojL8HtT5NQY9h32fp7Zx8fzY+ctHkAxjEndV7689P7smMPGxOspwi+7fDj6x8
3y+RQmaITZ+Y08Nxe/B+Ch5M8GNa4zVeXxlaXKP9HoV0bS79e6QMnisO3+rdZWYCa7dsj76VftFu
aBFiKo7ZQqnJGP0FZ6sHBNSV0vMh4jduaRrWY4yZ/Qy/rS5MzpsdbVDOlE+PYBiMUxXa5rAGgOYp
G9tUYN0sCyoaSf/dfexXYWtmvc7E6ZnTcD5yc3TRDthfDjVcOf2K0uoHRNyCKUacFBAZz+4tdY0L
LS4nsOP6JDK3+p/0pDgmrCMCpuQylotcsLe8fSf3BZieK8ya97awilYF56WT1T4+ecdbJLI/JO05
ZuDJVovEKqVYx+jynt5GF/I8Yg3hTbIIf14duzY/rTShj4u8cGVmmPnKp+KOEkG0juftBIVEV/TR
wnIOF58esEUEePXVgUP82DQCv1vs4v4nRlbHOVxzMFUZnx5fXtewcx0TecOGfHDf6qbP6UWemdEC
+NBjkDXZ2C194er5rBMQg9koNeZ5CtAIZYODy1dnaZfBU0eg3E66/snbsyKvDBQ401oi4mR0GN/x
6mWHdO7ZVJZfCy2zuyIvNZKt/YBkNa1q3aLhHG7HLL6oZS29/I6M7DZF823P6bNSjXpga7kMn/nq
x4JQBiZWfFGHMqZKpX3Ge88PyJa3XEVG5eXHypb7mDPDLalYU7TNYCZY4vUqqs4oucQHD+2saZnS
T0Q6GXStsHBOVQfF2nRepYqMajkiQ3Wd6ZuJAETJSbvOGYTCMVXWczPITcj9IPYmcrRRGXnIdtRD
aAWd0mRVdkJEt22IuR9q1bAYYHh9feTiYUsJdLoZR6TJEmawayflVVSsarqhX6ki/TjFMzr61qlK
PcOZMa5czzejFfH8kFF10Mbi6ZDeBWVEdsJZ52LIRbr1wdmIy3ha7vZyyBdDFD+opCahEtVcoP7t
NIWBDG1WW6nCBaPguRb/xAGNCu1M4jeziOSQJgtF2AKfDDvNXYl0ak1sUfFunn2ZUH9W8q73ib5E
bv4nknhUczKTXUrqnfe4+y8ZkgsLL7xrhgF9KHOaS//Tu4W6XZPHnCmqlwQR2X1lLSGVgl6avvUf
aEglp+ykiJ/Dp+WoNFrJJ1TTgPaC56tacq+giNr4Z91fkwakjX5x6LkyBjF0io3snXeuYo9IN4Bk
E6r0g8fZch26GY+IhOSExfFtOvrzYoHZufz10GWMuTbOVvVKzerxfkE/QZ+mKuJKT5By7TkHT+RF
vOg2qdRrJEb8ekwRWRLXdwiR+h4xLAx0CxxKfCrIB8ib1iRqQAioIMY8WIDPoeTsMu9OXAvuZJcp
dTVIt31TmxKk8ldF9Rfp4TjFUHjv2yvhCgnOx3DaEx2rgg7jssgRDgA4IWxvOWa7PhmVgt8k7PFF
adaVIfK0CR7kX9/Dy0/01BdcXAZqUNP0k/colqsh/OXsBoLVPbpIsUCQN5bDkwPK0d7Oe2hH8OiY
DV0KJE8O5ehGkwv8gVzij9bP7Z9yPKs6MB31kX2fdA22VlYWKaJHxpejsZX66hpsUuNBrGH9kA2P
vdkFVg4iESW1pe7efBrT+M6yTmXnOHg8ptWI9DEaUM/gaTGeLLoSDDZp5v+6e36RymhsynCgRPfC
ZbBzF+sCuDuxDWcNHrjDcWbEBGugXKN34j3a8LibNVJ/4AktfxVXnEYezByJXaWl1NDNQDzyss6q
U/LvS021t7Mnx74+dBo+rDhPKBpr2706SpZXEHo11Q1CwQjVXiNMUUA22I3aWk92uARlZNBa8OVq
qcZqf/Y9y5/Tdp/k/twBOOM9wJ5FsApjFlpsasZrTagY5itlgrqup1t9KO1IBC9UX+7ILfIT1ViC
gaMwqPR5yECqMQ6ZC259If8rst7c5oEIDOd7Y/JcoWpg60PHeGQD6rCgL5TgLnS88rhYIj6iqBuJ
fnfdOAaywcaY7dKEto9tbuFhjXf6N3rupSJmyyfyt0ga+hZOskW1HTxT4aGIu9F14RtU9NqvObJx
XH/+ko6T7ZWCkDgiUfOZE/YDcaVXSjQzMczKuLZdVq/Wba41ye3hWJrWnlWZoa5qhrgr2mQMvjJg
VXIBrAlsYdocCws2zIWbiHOcaDCfV0QzK5P4TZNInZY387AT6VV46YCbUxYDRQbZItts6Hk9O0nI
Xq3ubXE+TKX+2L02tzgfgazGUU0J+17Q6N7ge1G0zlcCs/RG4v+lHMzTakL5zwAan6lpErVBBlDB
xecxBwlk77vBmFUz0niw7JKIENoVG5o5f0WN0cJMiNk+KrGJPxJWKTM+LiM/zz6noZ7+yjF7ljd/
ktR8Iwn6rKS8yX4gRf565ns4YRNIpbnGZO2DykHLAgsMKxykC1mDqoD2u5IipKPMI1pMMma+Bn0g
irz7XDisYOKSbhC3JLXYB8MLcEUKnU3YuP19rUQetzASFfXy1wHuYdndoOSdmaaAFhEhkYw9QtE+
4xbk0yrFOqwSzcQiejCpomwJ14WDWM1Auyd+ew0EC4no7HAV+Ynev9tDvWpQab8PF3Jxrz13F2i7
6KhmO84tMk63Cn0cussZb7fcDyX4agR98dDX22kY1iXQFo7GO8mQL17IVQtqv6ChTFLyjpPOoYio
ZxT2ZHBXcY+87E8H/kR9xpESGW0sa4F5WAhZasMmDaFcBMEQCmCGU5QPeLoKAdYwf/ZDV+UyHQIT
Ad22Xx1qh4B47yqnZV884ubMQn6x5nQjHCoc0lLsiMC4uoPylQwdzU0UUg/BYgHpQBLmqaVEvpwi
Hs3VWycQBs28/9+WFRaMqP7xBVEjW/9NTziLXAC+X+7C7Uh8+B7/A3Q2BXc07FW7WF+tWPipkGey
9eSFcWmfgnJbp+udva4J9vRqiXmd3IhULxqn/rmC10BL5fmp3oTO7ocbOzD70CpFP39Q7QEPYlS7
2YlVJAJOaUwIsN2UOC7vx3XCAYM08sQQxwbzF5yI1Br2E1Yv8ZD7L9oy54O8nrJEbyUlHk8eN9XQ
/2NMTAxwlnFXFb47hKgTQJt/zgpFKtzwVh2rCA40MqlaREzhimITPBae7eOLk1vuFyQLVmdvLW9p
Ji9CQPcBXMVbbXgdtpQPsp7ObG2+8vtk5qUTLLgiodmwiNQbzec8GMsOIghVWu7DyYDpsWUmNTZP
ngwyrcNKaREGeQo0Zk3oleSfhPQOY32RLVLlxrPKsDQIAQdFf3Cy0gBDm09/wKsaWBC6iOkk+cLb
KEyUfp1xUdNoWcnDpLK95645RnNH8ScUzldIC3Y1mrqCT/WzRnvaEuKKBW5/TqfASHbNV4Ydltoc
KgLAXAd6n1K2AMhN9bdSTh27VTleGfVe4vgKXcunqaoMdb8mwz+PRbUj9hGON/zzuh3LFnCx1TJy
tftSPB+fNinnkxjsB2qKdo/RDcXBWNfKEfspZHvGR8xly3IHZAwUJPOYhdJKQRLQON73H+/t3dxv
V9eNo8nwzlNpYfSqsAdoy7dITGxITecqqzbMutMy8Ep6zgfLqVWXQkwQ7b7qoNqs6kHgbgo2mG2q
utX8pxVlHALDzIQwU+qQvKR09Yn4IcMk3g+4UeeplVlFufgCVpd/hC9Rs4I8bVj+WErYVQJF7dhg
haianYZCxoXeJGHOSAcqIgujH6X5tMV+Q2HnYFybt1ol+HDAZ6Kgl2GG4fueN30zoE2ujJYNPhJa
Qwqhpgtkoef/7s5ZBiXUgoxfWnc7E5MFOy01owurvjx81SQV6id/bDzMuaWtI7UnBJ6PRzqqL6gO
OTGTNYM+K1qDAC2aAw+DccL5msDIlu3HO0cOmkcyKbgpegNOfBtWPR8GU6p711Da2V55KSF4/mqh
H5yP7OHTU6xpXOUu2z3SPSRNAz7upwOnNSJTrQNJI6kacwvL9BpnCFiYyPJIduIH1CBFENMe6rZZ
8CVeEbzWA2c5GX5bGlX5cB3wV7st50XSS4bu6RIplFZLXWPO1SNuPkNIVj8UNfdSXD7tR9KfqF/+
lB9ppLrH8XIQ13NI5BXIMgKFFOazItxQ9Mn04HFDb/7qtnqjVi6IyGnj6NTOUX8WFQunNuVDJRdq
HOBDURJ61S4k29NNd6G4wxHIpXW9YCcROjF39CU3OkcbNzXSTx5LhSUl67gdCQyD3cjwngJ365tE
WSwwJ/SWmKTtrtbitla2tjP3A38SiJlt3YrjjNJxZ580nYTnIXcaXlcvCJPGFiPCK9zs9EdJVq/+
VAlP1SXaQa45ZAuBVs9Tp/zU+0Y76NQs1skGjQrJIY4WrhgR71IpmpacdF+5eB6XvTbvTORaIj3J
5pK5iGYhRHCRWjREtnTAJuUP/CX6n7UXMlsec+QPOqNf1GL0DOzPQblurGY96gkV2wbJXx7cLwSZ
n0qopWKTY7jXkrC/C+wJzZhW9T3x32fuNmjq/frSCbB/OzUm+CxeCBNjN8aGou26et3eqFh/pBEE
xTLXdS/+mpdn381PzfIpH4sPbMN3q9EkGqB0G1r5EgXm3Iv7LBlilC74or0Rl0QAP95S/MEJRI9E
/3RXGGOYWseFJcZGucPUwcQQDXzJI11S3rY5+KnQN1iapzBR8/syEhCeaod3NZjjdd5jdZOMyDwB
ZIqI6BcJCjgJLBZ0JLqKKhSZt5XN9KlLUyLsgVz9j+nN6lKZd/7a74z5xIDEo6RjYk5TUuG6Wc1l
ogl00iFB9vHl7TmihyStyqBUDMvqEU5PQ5nUim0gKqg2LFbuikrCtRiKLpp+a9QOeyGU83/RLV3K
IbMg1eDZGJRR9PUiTq1N9pOA+HwVbBdYZubJ+y+XoVEknXHSpm3DZnkPE9Yxh8ls14ah5xfIK7yn
E9K//8CTsPbnn56UTW47UPCF4kDmRZI6NGqYrQcH5mMdzqJ/rYepxqF1+/YLUGQy//SxOM08AEFl
z74wVTbIUMPGNeZWEfgNXMC6oYOxEMs3NcKFkMXEXuMRWa+lIgTpTf0gCq+aTWmlbIS+QfXBn7tB
1QdRit8pYtzxY51s42+UOwSaIEnyVm175RmfHJW3WvG8y/JyXt5lUceawevyWtfABsVo2fXs08+C
Qt26zUKpP3H3GaCwxhNkL4//4fTlAkI68+cW5o0OWbnlo4ee5Bf7S+IC+YJHjvkYjXWuElTX+AS0
BwV54/BrD1qlvCOn6Wa4Mwz1UQCen/yBwxPAbvGl6wdChZD4lwC2uxtFGDqrOu3jhmLBwkEFN9hm
XituXDnm5jejnzWhqoNZxxaSR+623GBmhzap6vfMW4AwwUW+9XIcZJTltuLlCNtwf4773jIA0Y9a
qOyRUvYpc06814G0MoMpJXFP3Xc5gJ/6x2JKWKa411IttBX5AWZZrnkTaSfThb7MqcT0MHTUB6MC
t30dGYLOxi0++f0L4jh/EKJfafT+BWCkrLQQuDax3p2dgQ/ufmDJjaWTBf7Y3jYVgyckhA/b2f84
BnYdkHrygecrhH6eYGC6sPucw0rHiEioguW5gmKRoRlcGclNzG2Fv0Bf9Ut/bKwUqOL0Vw6I9UHg
eRq5y/zHzCjl7GewbldeeHeMe/iyqg1lFBTlzsKTlYCF8WFdpyi8bnaW3lQN84fuk+3IFJLDLiPY
UW7ZET2pzG2A6P8yLNsrZzEsCxXjjepJTHzD9JVpWfl+jDv1wl1GC2eREFDnRcEsCI7s+gl84XhN
FkwbJiMSiv46ZmdKO/zD2rxlHt6dvMToYcuiy1NvZ85AnxnhIXZKPfGtC/X3G6WkqZNkqOEqmM3x
EIFVsF1OQXPCMx4EhHFk35RsIlytz5MBLwocU2qKwYg0hZWkG3ZYoDNDniq3iJSNU2yMlUczzQyB
KbPyuivjH4+CuxwWvG5r2pjVrA06DOqFzy8ha9fzHFoTepFJRnhqtjGywyAoxyFtFs7dEi5FvpDk
4+5t2r/rav+bIb4b4+HW91oGQbVOAoCyghw28aWsPapXlJthb2ZTfxk8sfrJcTwMZ68MenZBL6R1
SX05zG2I5NcADYrx/kq9FrBTQw8XDIposJ/qkKNUJi2QhSpqPt9X0sSyLotpgIOeSGX7VlBXnKsr
v5ctuVxUKgOBl1qjZ6xewDb7tiY2kGxcxe2KZhOKenQ24Tp+heDkbK+vdE+iauSJrd/nsmuiHe9S
rpT218N6oodozAueU2hJVXD+99b3at7WL6ai3+WyDM25i5JATpuXAiWmokMt+/u6vOamWTVvSb+4
ksL7RpWTSVTkSGfkjFz2XkZFjzK3NTrJDhfX1PT79TYcR46ZwkL3UfAAGbR25jX1Bqes8Bv/4iKh
gkAs5MzqVDGYcTv/etKmdiXthBBne9h43Gkc/fiBdyQCc0Bsdqv9HS8JnetgJ6RztIU63PiRwULV
cYan+MSh8bPGvSnXu5o/W9OqG9N6sCI5N4eMyN9y30mXc57oZKzXqo9Nl8Hd2qbRqopqEVPaBE/N
HnSvQbsaFrV8ag1zGG5/Ndk6niO3ltH6t+x0o4k+vOm1rAodIN3ffmWKKqdN9AeeXPy6AF9lZgY6
48UXc70UonYbvyKPW7+MBK5YWV5FLo1R27Nxxp41Tc21DeHc6oMJ61G0F+oUnYg9ZGYR+XDDJ/lz
OmdJFBd8T3ZYk5JpO+llgB/IJ9nQkgxAE0MGZ1MYAgDj0nuc41tfdsEzVANfNNi6aA8uQ8dwHkHr
pfoIPRGmKRvD/uaRlRz4rvf44LnggZF48sQHF/CoA9gfdGCb09mjTEtRrxrn1vva/tBayfl9mhdG
eUg79s4OKNdnx0flrqZ95PZsm5bwkg5mZsOVpKsy1gqsILvgxW9wB0se0LAfwJuIk9UN4Q7kLG9a
yNJFimfM0k3CnCJbin3SnxbSSjTCmsybBZ38Fg2sOwIS7hh4s6Ohh5az+1t9MNRDKCFi0kPXGE9X
k3uvYr0ln7uttmFFxVUpnrWHFef3NHJRot4u4RoMm9Lg/uF44JfvOd4GxgHPF9QaOrrW6CROvQTd
zKVj2lVuxBAGMdhkW0iUcQyL92PMW8p48gZ/OEMpkDw43kFgJ6WDTVoWEfFIzeg98trWvUAMKpMy
Okec4oyk6f5LUDzWrq6O2ooOal+8L4PuP9IrtOMRwVtkJBEOFgN8J0TSQ9ezgS9mSwZhCWVrVD3r
hgEV+kPCwPYDt9EDzpNT5kHffrWygp0Ez5BcXFrVUwZ7Iq/t9/JFPSQIdBXPpmQZ2PxLX1EC4W1u
CMIZIzlUAyIz7KzifSLRe22AJUIMZkLOE9qXQzkEk/hkFQBr7r/cY5LzoyLqqaK3jK4DQnDYE4cl
yPAqohjRA2hXkm72wau1N+OmjvkBHt9Gd8Jr82ylYjZncliXz8sZ6AyZyjURaxqXKb0FUT5d6kR2
FX91MgJPJ4eS3CE7QZSWLalM9WfPqdvH9WsW5q93jeu3DNGAIWQXYf9ATH62SRedgJ4XESO+1Ks/
RIpE1dqEw904yRboYMTbDFJeTJkNxIs08oBdbL2uWm1hn8TDwYsO4sEdJTDMVLOEdv9ys4Qm++kM
NOZN90d5pH6TtcZnIDBufKgwSThrN27x54FKyqFDnO1RD7At4n675BMW9AnTJf/nAajTFj+W/kbj
4jrpti4C+jA1fSasTD6Y0OauYZtfDqd7KRWWu1WTCDP9FO2pivOKugpT42JZ4Wod3/4mURND4nUA
csw+7IdMZO6EWf8o4bmgIwQ1cDTBiQ9nZp7Gyf96a2KflGfM5IURXP1YrZ+xKsUbrUB82n1GwRT+
ZVYTGZBA06WZZLmecUa2mMUCPyf1uQjLkuHvy2spm7iFYM3inO8/ggE0uBq9My3HcB0M9B0VBZmb
nq1GUuiOltvnF3xXJz+UzFyX0FPwohG6zqQuWTocXD0N5UPrRtFC+XZGXEqnomiEeaWIk20SV6R4
t0Tropipo63KQWjIAAf+PpV+ounQIsyzgSCnqrUNB1gcMuB+EoB4RV0BizMC5YdzqraJoCUGJSVz
v5nmgUmWY69xKoDUNRU0zsNqxJSozc/v2X12RDYi5B67Io7HLtzU3HGBh3qeYleeVFln96LAny3c
JJsDEUPT6R141a8TxQSuv6y2/F0Yb6urvhuKghFWsRUpGzHu3y27y43LR2JpB+Nd/ysfg5IrLXrr
2WlzQoapnjF1qtFbf5jehYw7POKsrvDAhQ3hiTGLGFvf51r37ZnURrrypJjDlNhlleIfMczpVE8Q
qLyMee9d0wVqH7HoVXBqkXvHEC2tRRUSxLO9tvdkeFovz0K0VVM1h6ZfynelRETxFRuAjdEjUS+w
2eb7XZLCxvIfbP/OGGqU50l6YEYuQLVJh3Zj3jVBVCI1GEfspMj1BZKdzL/BJSg7xLtt3wNM/KPC
AVZlvIv4gJDFVQCdf2Qj97zrCE7a6ldDvAW/NXzjinNWquhofb2hU8ilRc00xWoFMRnyRbRtsMOv
czwvj+jH/Q7n6/TElvDliI+7jKe5AvSXAVOk7wZiszOCmhU5NlOMmOLtNhBg6gDrYw06XAzmzAWA
cXvO6oALk4QWJlG0eL0GxmJ21fXvJfndIIOmNgbXOEGSJebtbLVv0ndvTh8dNVo1llyvZ29vqtu5
TTOmgGzyImRfIve/I8g5FmCFP+pz0j4oxLL+v4fVVS5zQn57mOikhRoNBdMkay8FrF0NCcAYFFuV
xdNVydxLjoHWHBpF2hMVx+Z8+aFb6lPvPfvO2FiYItQgN5kGahfMUAd6bvH3bdyilcNf/BGTMFJA
K6Gdculowx3pe7C9N1TTKN2Ixv6W3Xx7R3+4YwNChPn5lk3zOj21KAtTz1x5hHwUceo8D63vTT+w
IgLk9K+xWqeLXQ/Lt/lgEpGo59klEAEpWuP8+7JrVNTt5m0x20jVjSBpJ5wNRoa5tjB6fLtVl06V
3rqu7/WmC4L9yJ/DPrzIbl+icijMPtTL0iZ3sFnP/9UDbN31py9mfNPJ8G8APSY5OtpVKWcHw5Vs
VuWi/6VOaBxk/lXpcwUB+5OlEbGAnbN0SZxdU8Xvua+ZVHehqYKuy1ABWHWdGTCJ6RAm2/CX6EXu
hAxedHESQOUT/0DvOql2Kv8P55uqkAtAQJuWybpUtfFDU0qdl+igfL/xwzjFhmIsBi2zgrw5VTlT
oqigad2OU2Q1udr7E3oh+smNyl16z5NRPuxqcicpP+QlsjK16Q3MrCgFe7694ldyD4mu//6bexgE
HkeheDv6uR6vgJ6xXKUlrnFticy0WRnCaL5Av1Q6pswke72H3Bd8/v3iNmHSL8nTbflHN36htoUC
HIYRQjClzAbDRSNhBwhHWcNWzYAECY1wGtOmNYG5oxQJByuf9syMrsGgqtY6CuCqvUx+qyomggPe
sWXYV5fZpWcJUAuUKHOLThoCskLMszWhC3WfxhSmMYyqrDxe6tf5MQ8A+eJfgy15EICWXWG3+Gzx
yKbbmnN+5CBamzccFDka2hi9l1mZWeJicMaCUqAPIdyzs1GEXSqdvMq/nijkmVIg8X2SoptOO0hD
X3AMZMQxocdoW5y3G+P7nedgf61xOV8jnsIdjBYaT1URlj14p2gKW4q3K/WVZLP1UQQ48MUEgvIr
vuD2wfx9b/Izl8iELAyOLKv/SQXcTuW/5G0TYDZcyeuEuzZL4pL6mXPyG8t3QiC3T6gHk/ZfF6QW
E9LsY/F2+FImmhMYPth20QR4k7A8BCIGsZFpV4vdzapuGrl8QGpboKW5HAGPW9itIBUzCwrCPvvz
5L59DqbjMTSvlwpS5LF3Sza53w1fXywhHSgAFtBnuCLUy6BK6WavsCoduoILk5uqvhRbnNW41+3h
yMJy/PqCaYv5PHyctdmakIBTM+Bh2r8Yt6LyyqrLjM42IISK5Sk3CqGrcz/nq/AE5asg8zrgPvJb
jCkwdeFqHweOJCYOfDhl/GrQgZUYx3D8ZQZGVYrVuNZ0486/9Z40k4o8NPOKL8zN6ims9fVnhFrg
FSxo1xeHJ6VqeHCVgbKM6/a2k0wFSkE4AvHovuFWlLYxGAWd/HTy+5tiTnnsTfCRqSCyHpIgpCpu
OAlkrNXY5waZYaHFnDnGm6cteEAbZ19Wm9NkKA482eFeQtAfdWukaHyInN8bGQod3plwDiHQzTYF
ezlTDVHmIiQb1si1FYH9BhwdAyPCKa7y9Gs3R2arOuzMit3wRARqfJ7q9W9XYz7ikerwS7e8chDo
7y/c4LYiFRm28CVqSPEjCJsHMlynSH77gRbTr62UmmhX/63sRG8qeyN32V+pLIn0L8C/6/LU4o6V
u2aQmFweN8Gn7CHGl+UCLK7go5GS6Qm0kaXbyAXpJbC/Rsh3geQGFSTh07wVXHf77T3wodMYdZd6
qocjxNNwGdD6Cz0Y1ZNzDlJXiuEt0t6GoVGT/Yt5VJtHTjDsQWFErsSyfT4IqDEGqkpJ7iTSs8iS
4O0zM+dOWzSgrE3mLa2FBjD/PN2TciXiVqye5bKnG60PEg9LlzyrG8PKi4iKpZx2l5G04Gs2UxiH
XejFQCXWqelK2JYDWkWNxUazNlAMf513qvEYZG+Y6WheeIOfQxUNSCu/YP4TEBUgOkIUvLWbPFkC
QR2FFP0PHrDoRYNGy9aKjQ3DjYIyyGB5ld4orE7Yx2vl3GgPBOb8rm+Cu7jhMsaX1+3buEfoeIIQ
AbPD4jleReMRaIETU/rMKJSR9QWX5ClvgatQ7dtAwJ4PxWeX7vToRcgczrF5X5zx1YXT6PQ6Cxyn
iePCqDUC+nSrA2Jej17T/MuEvC3vr38bFa07LpfXlXaFon/qc9FIyhbMifSutdispHGqxNeM7YTj
/eiqhcP946iKTa4Jbi7qgx4Yq9ZUjgkmiaGNZCkLMIgM8LnlqKki6G1N+twE1hdDU/e/0FTKyZNF
349nmK/Wl3bIUODXoaRsj9Web+Yd9Hc11QkBLa/XplSWwhCzb1vjKGCyT0H8L9r0oIYB3N3B24Rx
ZcduX79P4+/wIFu8/9nopXqGWr9r8k53QUmJ8W+fzdPPc0y2rn1tw9rF+Q0jIPcmXMopAGs09mhp
BRquGoAc7wkQnxthsJ0BgR3CkABZbXCqGkFp+Ury8yIUjA5sdCQtpb1oVANQifWkXBpgT6kF2xbj
g7SZdi4ACzai+++/Nr/4qcB4jFacB+9kflYEUQn59Yh/W0uvBJ7/MiwIXOCSzy3oABf1fm3cFJXO
SAQLxatRRO4Ov/zFZtX843dwT9stffJCmk5bEicHgvgt9DbBJs2fa9FB1y7wD3OkyjMQeNKxdlLc
FoWO6Wf16hTrT3ZpMUH+vuIQEGKQ45klHWz/z6vDz0diIst24KofuqQLIFh5SUd8WvjTYgx+kk+s
UeQoRC7ymGtjKWvi96jN7vuBz3vqqcOodKzVUdSDufqKxyBjRiWuRpNHNmWyqSvxKTtu/rj2AKE7
G2+CjVr1quot8WDkYt+v2tF7cJi9KEGauIHdSgEVFr7dSQ089IiD8YJaWhDeV93xcayYp36cyrrv
S8azbsl1tW8l4xxvJju6MvNTm0AiZITViCqVSIZfKML9rcpLKXAS8GdjQUb+n9caQlV27yJDGY0j
Ii1gK2K52g2VgEkjrixKomXSiS65mU4kDtRAssUAbaucR+Uo/O2H6967cNQHL/927nencdErHLTN
jXZKuL6GfKBXYYCT2FVx0g5D/o0qiWtYZWIykiyTSamdBhYmE2wbbTDG6d1CI6fRroNXvz+dHb8J
cRUALmwIWhN1msYXANNQrDfnxTWw30JB6KRbELmt8DitL/ItvPMzZjZrvXGgC5EMM2hvq4Od6n7b
NHJuz3nAtKz9FLwe42fmtbOU+YA8MHsNu60/91Q3qB7DDKTOUB5MBS+YmPjdkXIbxWlhhpSTi5U0
YoTqlFudL9gWmlmbOMpnhhqdNtKrjnl1NKZIWSs4CM4+EVRV5y3iwI7uj6fyellFKSfyvXq7HPjV
oYGHiE/a6Qm1kX2Vsk+BVLMh2aqhRsfLh5+sVYXpBcXcRbU1DCHQWJcYuvyA+Fv5HGQnkErB1tF3
67x5+sZINFm7QOCwRbFlFOXF5UbCpc6CQFc3QIZgcmLRFsJYQsJiiNw/ASNm3L+nSlhhh0k7EJee
3CpOEgLi5qVNd+pXff9l+GLRcGUFYEDdbSBPzlUazsu1j5nGt1iKcjOMCEsoaLQIbAmpl0lu5Lgj
s3Q5ju05PNsOdESP6Ljn840+34FdWF5tIt3BhHT4YomuCPzz6WdA6LrQ6ULZ/rd+hsLKkNqLvsQh
JD4FQarPcgHX4c0qDX+7Pkr2yx6fH5SqqXUKM65c9FoDUxPHZcYuek86jrNU6ByIsHXh92rbeLOf
8IL++XVkLHi/lOCKOSSMd8sEImfbiCiauMu8WNCauhaFL0yJ10p/d2MnvNZZukiHognYyKaB604f
q92IQQMlLV/9B9tbXs2FVfOaGbbHW02t74l/cnKttuueqxTcgbTsA/cneC/ofjpm5xBoQfFQvsPg
lpRO/lAFiuBhEkieAi5hlEuoRJQnGFjdk3S0mKiD+/IiL+vRfY0lG+kkn1Yd+WFILRgj/9DyQ8qS
nxKGQkB5Gnqq6kkqJuftUxOdycHhliiQiglLRPM2+3G5IwPwS1Yg4n685nDg0hO/zAtYRJu3XVrC
dKoIfUspeAZgkMzLYL8PvI1mjR1nMKrQBVMtkfyLrKY8s1wZbQRJWNUJxk/yRiGaTCTJU3Aq8EvP
V0hOiUX1CpzZnkwVYwuwamLbXKI03Eub+oTa9zN21vpE7qBStQXeaBpsX24ObAa4nRGPw84st3MV
Rfyf9GeWF12ADUQRloVFUEOgmfu207ryben5ttsZAxMzoFBM9eEdG8BMFsVI6AmijSsotRF7Cp7w
kQ/yE4N8sFc+dGGD19tDJpRrYMkbJCkXrV94ZtUpWkvYlIxGDAM5xln71HagN8H9U3W0gyGz4e8P
pLVLKiRf47ybLBzBLBhhP5NNzCIwU02mRNbJJy0MVh67cuQ48T0s8vmZFd3qkq9hl2kF4XEG0nbV
nLXDHbFN8YbJsWmt+WEhj7FyhqLLqr6y8Lp9VB7IrLizOQ2NT3Eq8YoE2uISGXmdY+aNipd4P7Ub
rJDwnGk39UEMTIzUdlbRBOTwTg4tt5vf7IgM8WA4zmMFI1VenHdx3ez/2reFc4+QLFvMuAIBr9xZ
i5OhoB8Bhlv1p/99Hnr45dYRBYdnknHHzWQOWNyXeBWhMABfc0ZuFQrRKk4FW/+UyDZpUnicR52K
1TZ6paZO4TYJbH3LPkFticBRy9YR2HmLhFrUk+BqIVk2MDycOCY1LEZQ5gtXDpX7UCt6HGXr9Kr0
CX5xbXSmF9CRmvPDWBWSO3H2F/sF+F27u/7ZLlQ3H+dMb40CUtWuUNlM9qrI+0pODgBSdRr3L7pG
v4XrxySYiG/r+OSRdCjAuMPoxo2WN72zUAChI1oHuFKk6JAqFUppE+jKzzPuTJOYnAZ91LyIC+zP
ReV1jIs4BvBP6Ly9+n5dXpzeG2auaNTjQQVhAPJKygDB8Wzq3mcs/YF+EOBoqHDFQG7SA99ex7sF
ciCjXJ+5EG6VVfYohRLzZqGGY60AycgppJqrVdx/wxR4UJlv+Rqhlu+1TchAelxflvC2T7BY9C8n
kmCkcXxO1tPS6WItsvy2EdXr173gDJAN1oH3lCtOObKnf3QsXAHwt41dVnkT5VXWneX7hrNdxd/C
3ohl5kbET9HWdJKTtfMoLy9uD1zOCRXBZ2ak1YdotLHLgc9xRmIqAnVVnA/muFzV41B91J969ZQl
pPGKyzlw8x9Lq0L9/KdFa/Gd4KIiqoay0PwacqLsRefCRZq0oE58LkFvkKw2P7yhoup1s9YOjh8D
pL44mnK1bkd69xyi4uKD4FaTTlYXIYNvMBq3xLSGSofiAXNKQVfhdsMFboYf9Z+R2A3zliwWxqIN
nOdoqpXZ6iVRJOcSatGbbVY8K9eylSQnip/H3S18hYQ0h1I5TBOZPQqM3IVd4gIjibXX8uuQF6rg
/wxK+Dntx1ppNp40BKiU6/svzM2UmJEtEKIyNNtwWdl7rDpHtLSQxAZ8wE49nOt8mL1prDQb9uVg
gB5S9p/m4XZdXsIN30e3foL124UcmooKV7OEuT3ecXjc+hlO91M3Bjj4ekICD7nUTGXtToYz1bBu
RQ2hjRf2nDMp3OgiNljsPP6ajhg4A5NeBInTKaCvc8NE4wjmo2Lc3VpGhY/Kv3xYaFb6f9WpdbzU
hSZQ3+kSt2y8rph64iEPBIpUS/0+6ti5LvqDdcB3FmrRVO0G/FYVzc1LushDWq8MQKezDviFd7f5
3ISPFa3XWRo96wN1GyCN5v1yktTmfm3SaIMXlDSe206yHEgHHMVhRk+E/DDZkapiYGABreLJYrpY
TrSAAK+ArbdFTZqHeHHEBRRp+ZVj75EwOW9PNOWp5c+CFOG2YMZiflINPGAik+7kRSsPniTrOLgC
tVYf6U72/8GRpFsMihLUNgikdYDdTs+FQB1/GTGuNuK4yDXRDRaV4UDgyUZUDneSiJp0bHOVLBuz
brQaOnxz+ffPgfDiN6Gejf3XK4wbj2VjuPDKwlByKhegqVv9NHU3s0KbWx6UH0g632eteL01xa5R
Du9oWqOvP7o83ThANKXvos/5KGg4+vkaRRe3TeyBoB60rj2tx2Kt7akcOunr1fDsBotGr+TrFaDi
iQA5l4gYP761zfGz2NFDc9NqsIhhgy+dNYl4q5uNN0bvLvdcb/DopzDtP/v/Ues9s8uJQWuwrCRZ
jNUahpDcg00QMtpTS5fMmFH5faJWRNsjyWW1fic5uvK7tMO+k9d0HfoPWbU5rzcOyAytUqwb3z1w
PN72gSAntMsFmh3mtKzGZxSG/9GqNgsFre3cCwdlVTdgpsV8jCOeW7NVhHLEOAyUDcZ2X6/alg5f
1vi2+ehp4zMHdePB2qiPqpL40HMOUzRTtNe3s//qGDLTf5vXuJLPhgOYVKaCqs+d2VJ8i9PyPs1a
kMHrRxOqSpTDJsasznMTibSLdUrmbUOIftApL0qYGQSFyBbUTgKpwI8GkfwjUrnN6Y0jnIo43+XP
ks5LgAqX3tHYeZynJf7EFOtloGZZwL2Bd2K/iesCKQFXJuxaXKEkA8sl8GjG0uXdQi6c4gesU+mR
P0UQLiSD+xPkBiN66PsZ9OlV3huEHQFDYYkO2VBGIO3Usza4+NYgL7y0pJJKMVV/kwl9MsL9pU41
jsNFJGLrCaxLaGgEIP9pFWIq8dgiWBKBTjrRN5q1ZBnWTsyBB9wK6s0tCh0cobcNw5Obslhz787C
tzlCN8p/TMgWL4j+Mn2xx+Jh/8iiSTMit8ZDJMKl3wqQUynNv17ag+lrw47/L3uDjxmdj6uzmv2N
zbKSQQyOE5bd4oDqWEL5SlmSj+BGWbB99kqJjpPm/69tMqeg2wwNYNcYOH9DRQ3sq8+GNa18ZB6/
VgLkymLoLbHFe2nSSz+OcVBpzVobT4Dj41el/U0LxDCoAgGfh3gy827rMuWCQegnaegw5TIg5Cue
K41mHCtv+TXwnYedl46IO/xPrQ/3n8Habxql5aEuKvMvR015Wu03XUGrt7FQQaNN13JgIzPEaa2+
1/FxX65TAdvCBxQ+fnAvhgM7A391Bn0cOgUlZELQGU+J1d9VsX94QfyChh7Fqt2DyHXm2RPEmNsu
awI5B+PFKYNeSBBOPMnNF7/MLeWANIaOTZ8/ZOXJDbZ4Qi8RMwMsQIBfy8HWh+29XTNRUTJfanhA
MZNu0lJLZVUdflF6OQuBGadcM5p2X1fvdi0lFV7D/G7/zeZYxAdMSdkMWiujcjZaovUFY0rqEksd
+02C9ry6LDCe6RFQ20cDBLC0iByXmGs3ckmRJtcjXni4HL84iXyi1+2yZLOhjfk+VmfIv2hRZouZ
TqrHlYdx5k1cbg6PcDPfklsbs31Nxqt1rEYnGGgYwmTnlv9+L76MxtzuQ9B2kTYQqj7WaAHeaWyy
lMGLXFwFKuYMFGs5V0GWCGOSB+FRjvmP1UY4bietQTa42TUz5ahrdZDF0CpLwRwR2hE6LC/ebcwf
IF2v4oIHnQIRtWMIvvWSvdqCzWzMp60B5kqvIkA8ssqwlrXfT97KXrh8exJUJbq3O6HXURby72Xr
dk0kZfBHgGNsbDczvLBjnnIZBldiS0z4RNC9wwa1zboNsmxN6ooBvqkwjmKfWkzy7NtkfQQ2YDAq
mrqRN6lZVK3IsBUch+xyYYLgPCge4cgZzE8HdKdyQ60HOJSTrz22EM501T5dhKll+D8Nic8drw6M
sWUglIuvH1ZOEWVHQRqUQutIAQJvPjg5EdZDHSQF5K7/zL7FRmo9FgAox+8MSEMfCTYVWPE/fYJM
/XTI74KfD0ltT3sD6owsGI1SEWv1to0sB7gjVhJ5oeNSgk0VMXxvJQgO7Xo4hZA7Zp4OwHIJrjUk
438Lf2bwJud3CAbsK6wUWLhf0Yq5PEDBK7V0/xRI+lSiAM0M9Bq0pn/YZZLdSn/a8hGR1PcWXVGa
XAvS7I3sBdCZL4mtv4sinN81VKLAt8L5M3HArUstk6Z0si8/sOVrahllRY7UQMEnyg/pr3bntYBH
KqaU8xm1R+8AOKZ11rdW3KCiKFmV6Ms2PxgVo8QT6XdLoR5Z20EXfV8C9Y07gbT6dFhOQS5yyVUv
TASIV8uD3YVhUbXtmJawk6RKC71gY696qAXsdPHrJC373qqj0j5jelqBQCyWIh0h9L0OLGmqXbXO
4PiS7T+1UDo1kmHT4j82WTpzt5wlMSVM+eRoItLBuvf5SlSdn4vYkIVtgAqfEmpPy40irql7/llw
/nBwiiYKlJVPELZ5ZsF8h8hM7P1MUQYZM/VgkkY9bcxxGPZcKPjysbGpJMEMcNGZuMP1K5NrZJKH
qY+DYdvOBD91KPlDxbd+eVDUyalotAFadEr/g6DhlqdrNqrabTWkwvaDtRkGIIa5S5vU811tIMiP
ODLx0TAqhQuiB1jQL/thTsSJrszY0vMJJSPshBQbealhfRqIdvdswmHnwceyaY/vTV8LPhHdOCfY
fuAUkEVbET0TJf8kCjhXI0CgaTIcxeDPGK/2C3ZOF48g6JLnAaeYp3lSvGJrfYmgUUxQkvh3ch1z
aZJGPKicBgvbJTtjqa5suIoLxE2zVQVhB6RZdbcgE00WpBOdO14U+svDTGSHJEhSszvczaXsHfo1
0Vw0AniUFXdfjDo2CAZZg4boApHr5SjJlpmpB2i6WhGhb1I/sjYKuonggk5Fe9W7yAe+AmRM8zcV
m5sCjn/Tshg8y60eqmH8CoJ9F4Rc3/zZOKh7lNwcNGCk93HTw+Df9tpf1e0BVtLoqffMQ/bsAUgw
VzoCgt7wqQ4YpeKq9tqTqdn25wazJ5umXcdetzNDQX/zEUtiFlJNoGMMzWBITHDSdFvApv399IOq
1aM80HE5808WwxhxNqIqbLrJi8cf6H0aY0lgIuPyt2IMpCKscnU/uNaIRckN72K8Pl292Le5HpA9
2rncfeRs4gFM4BrfXQRw/A59F7dIVzEcBUGV927EKdqP1ya+wnphZhWUsy45tm3LhKJSE4i34rFV
vQ/sDCmFcX1HihUc+xuRGt6sF8gqsGuZhPMSzGIUDeqFs12jNqwX8po1dOy/d9TDkrEIOi2wOL20
wwQodn+xFBiFxwqXrQI772Ti5plwM0j5wZH9uScVBEgWgExnP73JVP5Zv6R5INgiEy0OZZ86CI9+
1W081CJG89oMe0oc9SiLvs64WK+QTaBFxXQizhNU2+dekgqeF186dEGyf5/paO3JFQQBkOFPt4oD
U21ek8sTO+11jgnO0jcy4MUyOiB+ynYV76bYANV0lfuN99yvPD6/fpRuW6hIbBJK7Y7QIiyVzTHn
Zt+Y3SgxGRsqhB+jYX9egPlfk9sKkUhSwgxRRgyC4zA8I/+T0kOtxslGAHiL+QY86mA6+ZqClmwn
0TsNDvSLLcl3DkAvPHxfZHz9iUs537jtoQxfj2yJX/wDaPFqLxbsqmHy0DDSBoZaISuRpzIR73I7
UkP1HFbUkgjRSB/G423Au7D5+Db8MYWls+zvO4Qp9QcoY/5Jg40cfO3qZK9rBr5fLdn8CA88Jk1V
JjSH5UTCZfqhN+g41RcxbU7xrGFqV3kuHbFE47bYNUEXZ1bmhOum3dv9cAsqh2FC/Q2jpRO7UfWl
Q/4hvdiTMuis53BdX8WZNv3pzR/OnJ8ClLlfpQ5096kh0tIKibXJWDbejBmcEfCx/UdXi1bdPW62
bHJxE5TL3m2joHwlWy8C2iIFpnmGKTdpxJ7rYP3xedeyZQv7zD4RQVgDyUkyG1m2RjEKC4uCL9O1
xh3nsz205cuvmrvWPXqLI8yHXgXWheiyivklI5fpo9nBSvjP/c52ueRwMz8K9vvOLSE3oLY4PcAG
NpOUqG47nzd5+K6CYB+RP2lkfmq66j2qq8y35ilG3h/RLR6qLGGb8d1XmO+cJS0Su7Idoyq8v0f2
dWfraxRtJutpuPuhuHR0bOVPdJk8DgQjHpMhBkGXaGPQ9SzJi05OvzGh24bDc2bM7L1GdF5R9sXH
5utAXcydswyRJkytYu6BBJlA0z0NTFEQdG08cvD3AftyH/MNsE6s2N8XEp7zUUL5EyivBMuSOEEb
z/tKfja84ymhQDncbl/pWwXfeteIu3/6q3gpgORe/OMFZnoEQLjdczQSJ2YOPkUaWGEKV30gZdwH
JurkauP4EjK6OwD9OdJ4s0p+XRzzvr9HRb0qH+QvucZw8EW/wD4loUiBmsnP3IqywiAPlw8226fZ
2zVyJ0876Nt0gE4Z2JGGSgLfyjR4bmaSl6l34P28l2xAuyjwd0oYSdmznO29VXDoieAfv4YKteu/
9+Wfov78kRtOX0s3Px7O4VSt5LjRHBQEc56MhSJ/QfIw5j6v/FEw35sSREfi6DW53Hs3BIUCaUfe
WD2cXkGmg8My2k7la3Nvm/pPX5onp9HLMUe2RPqO+3CIckSumRY4+VstjyiAJU94ak4VEWif3fuH
ZnXG7JrzerWzHuErfMjj+PTndBGx/kr4Yo8VweCpDjjoe0J6gw+OsYQAVQOFqpLMpcfoUFzGuSJ6
HqC/HQhd0rQYoi/dLmzjdUW9+Xda5ATxcnP475KnAnah3Q3hL3us4IKoWlhpzEyawyKZZCCpSuWk
2uJScogHcomnT175ZZbq9O+zgr/2lA3Z2d06ikMitgV1xXzoytvrUvzP4q18kNd7UkEzXmafTfdZ
RsvtJSGSOheZ5b0XTaa4+ALQhMHtNNIB1YH+Mh6tUYM4Kihs3xCCW/sjOyPsC1BARFA2Tq8fZmjs
4Lmogg+8BB1GqHOzF3gmnPaM2UKruR7Fre1A/1blAItvwbjIoNn+Q1ZYhDO4BEZFwLosujMTxw3O
/7KoyNBkmTbqZ/Vz0i7Kg3ts6oas2qzs3aE8edh4xrdAqbQprf8Odt6Keh4YWnsqTsveQBm1XpjP
CT+neAdO3E0qN5bmIS3sPqwBc+kTUeNdSTow+ciL4C1dpyfznWdvuBVzcQmugumoXDE0DrhpZ9RS
RAJKCUuipXZlu99K4LqifcFhXvDS0Z2PEJ848eiDr52923klymaKvVJMTWaBpMPWMBB+lDH7DXPK
DNGIUo7jlILr5Zy1xb/45+JaUbdC6CN8bAjeAetxhl7pF01pO03Xuw2DaFMYtbyElZggEqQeteuu
sC+V5aq9al41l697qI5qgsZ2DzglwyAoAJqlKwtUjn3N5xppYQr1s7dc7bVTlgYi2o1dKwiMFK+l
/aB3YV0Xt/HCB9RYJZQHF3pg8MiqS5A0U/0/Vh+KzsxPuKQkT+V/WmdLzzR0EVA5YHwmyHCsrtvW
TucokvLDYbXr+Uyo3UCdBCaJHwMyl4+2k8rNm0j1syBW3d6kNz31sc60EsdwMT3ExljhCrYDLOwE
gz5Ih31HnCa5L7aJg0LdLyqyhCpoC1/SBSJx5BCTIZicRuBbRV+oOpbyhxf9/73z8r8cu13rcAHo
+CGamRsTRoFNv4aMcGRBVLm8NukJAWv9Ki4OGmPVcuFo9uxkLW716ZWjOXHkf37tEJ3Bz4gC+RLm
sJkttj2y49FaxfqVIRYAMwEs4P9kjOcAhnUvNEdaGS7Xgfd1eSfFv3icQbuimzWOxIqk1vDcX+tS
bhOMG/xvvrAMN5j/78qwqUtF2Ty7PvExza4pluG4B8Glce3sEwuC2+g5lD/x28USoJkyFPGzyPvy
GysdqhAcisU9Mx5y31qE9n/F1O/vKm6/iBsKdM8UAbLrECykHatnDH8kbtpyhMhghejvMJGkhOEm
/STi6cIkBgDKvfnaIR21Dz9FOjc6A/hcrPQ8TwwvNG/6eC0jtrBexb9HC3ncl8uGkDTrhYinbHuX
+hehP86o92M4wub8pvlo67DuY6zFd3NHkAGzP72AoiUp8oNIqzhjvFCqAEAe15G2AZVAKfKBrVho
1GE7LebMLR/8wVj3cBwnZPlQgoK/O78jXO4xRROvw162OcVQyox0BrpkgQDXbvN0WKEIxAYkTi0u
eRN7+Hv3OgXL7JUE7nrLZuOVWJYJLBFdXkJD1jcAAIaqds///36AJKr4tJoG+QQospldsLEYvGl3
WIVdUyauZt0kx2oNQnCF7I6tSEVXT4CoW/Q4nbJFM6auVZSHqEFTS6Ka+PTUMfvBzgnv8VJMfacU
Ijl5hLp/OyHGhIg3i3Ab2ONQqLlsdHmdgIDPgWn/hC4PWttg/K8VzCzZCpU1kkkoOGuiCLVTQy6A
KKFjvXWUHe62mwjLLIVU4W4ihla9XePBnoZgUmf4/MDRk7rVHgWPVsXTl0ftodxKg8ZJ8jZW1JiP
UtK7vtSUC8Vo/EHatQTW48crLo6si+oFJ2c33Y+03E1wplpT2QPPctNCD1tt9ZoAjO+Ea1+ny5G/
0CFqZOLyGotvaYBxg4ciHODFzdor7JQuM2+4C+dDwbzCc/YjZooC3pbOcKgArtRkmwDqmzTcJWmd
8kzR2QYsOxEIk9DyLghgBRbnSNanQ9lBr3Qf3wMUzYLwjDO0TamafQBHkooCkDiQUFOc8dZtL13o
ZrW3JS3uXa3wdl7GTP1z4Su4LPHZUcr7UOme9mY1CyX1C6lv4CiJZvC1rDW6O1C46/0EppoYHYB9
fzyN+iDe+aE+stF4jK+hGwL/UZ3y7xfo6retAtwWxjA07zC76VvErgDoUnnG0Cn7AOGSCW0Si/yI
KTODR2z1/BrRaota4CuBST4iO6anaDQv513qczXFV/Bd97Hlwh4w4lCOdqi24A/qYe936wfk9W9D
1ou/thodjtDuQOZL+kpIDpSTNFcBX2hhzXbOiL5gXGhWXLRiizkA9LWUsgew0GqSh+hkSE3ilN42
z4cvCBeTWUvO7reS/Xah9ZQF+m12Ycu4SND+Lz706vLyNHA4hTMyAUj5HK3rgdL8IVxNWMzxkrgc
bqcK6eCVqSsgoo9yE+3LNsjX8079+t26E1fawzhRVnQTxAsHxCfSON28XbNgXFsAKFZ39jiq9uq4
hV94i8xSTSo9G2vtKq5xdVnZaNhgh3GgflQqd7P6yc/zpcZ082fULZaIi79h7r55wTFVEBzwqyw3
26erYntzhfCjsAdIl1MV2bU79Xn460qMUIjNhV//k6nH0SaDKrJwY2NE/CUgO2OWyiJ0k5llGm1x
m7DEuKbqmXVOVIwkNipAKopVC/89PNGkm9DAShUpQzMANmTFNr+4/oR8HIlDUADeMxrMCxXnc/x2
pSdriurY1saunRNx6IzHO7S4QKe8egz7M4kFIaAt/ELgaUSdIzqTXAubQzYI7gNjrchXLHOubwJM
kVzRPCxJc0gpZae1VI6zFYZel2nA0fKLAPEjZxFc3UkGK3N+9Oqy3ryAtj8N4EJ/E1iplGP4WvUY
8HZLnAVI6uvYDecBoRZrxeL6y/7eD1diWxf/0jH1mmzDrKCmQFbZZQL+LEGP63cD/d7rFbIlfY8e
FhByF9Cg8ESnJwe3iHac5Rlrd5jM6ah2s6mSBIu0dUgtkiYX2h7tdbg1Cbhvi62m+o8qTsZo4ock
/3zyPhBzBnI9COWwkRZDgbfiHaxiDQRyJdO05ZnmFfFn1x92Ui0xvBQlTQtrN0if69Rok3mokbyd
ibfDkFrulmdVKRJs7FWnyoz5kzNRcPmBYojjZ8BIBr1B26N8fq86HKpAVFKJ5alL9DqI449zKUCv
cfwnlFjKIUmaV7wtl8zPnF3N245hMf5zV1K509GfUniattek86z/egrxv5Q991pUYlkFnbWpl9GJ
PZtEAwXiNPcaAWwCkhZFjKM/wxJ4tEzcpyrAYgyDk4ph/sWEiiakUF32g4qVEH1ACEeSyWhT2Kk7
BKDVi/cq286QMkKg7UVDNfoPejeFpbDqxpaPc0BdXoNJ9E3rDvCK3YA4R5XtozVjy9iesY09+xu+
qYkPhE9uROAvsG9AC02aBzOAeOLjO4YPmJoxftnhkS05JzSnlCgAhclVKJhYwexhtSw20D6y/Xva
L/Yzl9S2HmIyldt9bBk41zu1BbwnlejpjCenuPw5fytOR764agFvcD/YmGAdpjh6Zd2tNGRKOfAH
2dkmD3jShWXbT7Hxc1klUcMv6o7JgyD8/sVe4qnoubbJ5SJ4/X+xqT3icwHF6TsJ1DQ+r+IoQkVu
rTIWxJJOdmKyS5G5X6ZVIooHwTkw59H+0yQe3D9RePU3BVXJ350tmwIM0/y+6h0OQnjlmJNi3UFg
pL7sCwK2C205KgaZz8LavslBlV3iFlmSgmOTf+HAviKydD0fek5YUDNM8hwAP5WSKEIXeBMZlsFd
RpKz3FjPOWq5GG7WfJYQ2Lxfkp4aZllybr57nqCu9JIMl4o2UIV5YzxhqC1t5xUmo/0W9YRq4eCj
iJn+QQtB0ZhLb1emYfSB10Z7CBT9Sm7iiN64rUPJannuKGdt/635WM0ucwAEM0S91PMhv58aOrHy
WRreZqx1I+56GdU1eLyTX85Uj7PNq/p/l0NT5w2A9fEp6UkHDIvIBVV0BbroJjNHTNVDCrnQ11HW
PYzoI/IdVO3C4mHD+YE6D+XFg+1gMNewWsAPq3S3anapo097+8hl/ajuExXWZiLLDcxrcaHVGgxj
JBhEU51QcwnZ0t96UnGE5fECmBcom7XWZJC7kDc6J8m/sG4zIcQ9ijmgh80D7MXYJ/GCBv63ofy3
w6zDBf592G3opn/VS61r/AwfJ2dE61y7WMmoZUimBX2ovzG6X9XzEq3N3Uotow2H44ERE2tkFWeu
kSMEQ9TrrWsubqXTgoaz/ApL0/uNkjl7qG7sNRWHJXjCcM7upGVu6npnh/5KROl/I6XL02vq9oXS
cG/8M3x3hVKAS6S6Tjo1xGmHkFwz3Uqm2dD5aU1EeF3i1GePB4bqEtlO/hCgysLRZHbknPYHZVqQ
6Okkc4chUXgF/h+pfMY4BoNHFvtWZvvqeT0EI+eqAtGOARI9CDffw8nMFe7aQSrwZtGEA5Um62Dj
OmlhJxhYOJSbZCs6MBHXYlEcXUcX8QDmPDmBnR3OI5q8OjgpmRJn2CFnALLAxvxORFuC47kiZWfK
LYuz0urvfo8NfJrVPn+c2OGja12w4ARR50T/R+yw8mHN84NdrfNUsMsWcUlISSAYXRxm2+C41wxm
vHA8fROE+uaquvoXi7S9f4cx3dtvtx6hjnC90X7ALYaoyV1OjwV8bhzOXN3iSR6IH8dV+JTRCTUv
rwOgM7feqQclzpB+uYkGXMsHOrLRm+KfMf3NJJleVbGD+Pauu4Kw2+zC8blqAmbhLzRZO8DyRzWY
sqcFu3VvqKCEnNvw4hnNKHSUklC5ve56COqyY/YCaXKh2Q5Qj4qOY34GbUvhtKLUYXp7zgZzGm59
zvqIMluAYL04lbe9EbYRZIsAKNJhSGtIVqu5j26EpzTuK2poRSIA8SsRhb6KZcDZ9ajBkmEq2Upl
z1TK60r3oxlevz4i4Qv+UEO18MKIwbmSa1raULz6S1YxNPW5ezLwtvbYkXBhg0yqXre/V0BdQqFE
h45nNe549gwvY9BG1jqx7+L6JPtr95ADpv1+lP3TOhiLf7ZL/chJ+90zbo1oXo/g9sWdM++QJMPQ
RJr7MxXXZoMfbcJA8i8vNs2NH3ndOhT4j2jRJEwymDO7thmbS5Ny0CXH0+ABi06fNyI28PBoFbVu
X5/GUo3QSkEghGXibhFnzU/2T4CU9te/4/h9MM2BfgUGYEhWbGeWX27ZLexVe6Wtlqe8RWL3uTaB
HVvqHJZ8RIDOwPwoTOfIJM8Y8dtPxaRHWjfo6hwVSNqDCmCrdGonlGtDggGv1YcRMS1vFzGUtvW3
ciDiDLIjT3KJgqEdkwF6fhc1jkUEvGa+2SP2z6ElwgLzWavKgmYLCa9nJIO1Y8LR0ZJgOCKWQRcU
QzD/dm03/WKlWHZPAfS63cLLi6Fvi5WyXcifT5gJeziSiLkxAavm2r39OHYWw3Ko20+49R/t2HDx
yjU1UNw5sQJxr0CpHouSyCySxWLKaEYGIkK7OPXy4uCs7eZ0SzU7DISqRSfIFdLSGHl9xL2Bi1dJ
0ZhaVpC82Z6Br//3/5bwHDkmOxROPFwM6yisSbRMPMJRKiD1UkOM2B/xNFVayZBu6fdBtLN4xLIp
oNgKPcZAHUAcQPbhAdGxFt49RTS3wqvAyLMiCLufYQ4NafUUaZrTDxNv6hA2zRbl49JDh4DvuzaK
7A0f8rdRAb7GISUCyIB35AYl8mdLk1t/BAa6jG9VqasmxdcIxVL+ZY25j1shnCOMc18uhv8neHlv
ULYsmfs8/NytZyOcfxzIL5GlIF6hAeV/d52RBO1F5ZUxQBwcdrokAkPCX+9wAkkSgsAhXX+yDZQg
JP7k4IgCohrUPo5NEd8PGP3b8Yw0wN+zy5ME/xWEn/fpxdYPPTwSgKKV7saBlpJcWgS7VP16A2bU
HqhDBLUV8wphutxvqFQ1s6qvNpEIx751k5N5ZtUWCKC3J1tgZfIhjMAMESaTBY3y1GSsnFBbYbQO
z3SF8dZOZSY3W3V8b61VzcY4a9AGxR6vLJPeR2z8s+ugn3O5WzvmYMNDjmp0LhIuhm8kaWaHPiGr
JDdhZBMYwEH814jPVopO6H8xmRiQ3Fm6aSPJGAPmEVX6QnFdR+8PXGFRdxsAXvJEM797ahpQiXzY
Iu9rvTaTKYw7SnRKBWaHTkQOTULbrrHRm0huF0gybp0nG/QaTf+5HOcmtgB1d7PEovmVuq7MYA1R
vUmkxyZTWntom6RmzyPeMdJmS9e+YoMS11I6EHm/eWMqjZlDpTxi1I6UXTZ1z6ll39cXsurckmFs
3qlpF62W9yFXrBpg9kIC/p+S3n1LHm0ztOxI1keygzafuRb8hAlZN5cJMlpN8Oxjbyudy/Rh1nRG
Bn1GPzbZEBH/aofVay6JvVDkegGh13YbY7l1ckruGa/VJR1HHe0ThkQqdMBHIbWSPwTVAPz2GCa7
hKZNlmvBLJcNYu1DUzFko9zjZgRJJEWEXwzypHliu+wZlL0rNRABJpxyGZlUK8HeltWXuyHJ1z0S
QJQQvEh8EK4nP3lrFH+8zucG7VLuqelb9mk+oAkiPBolkAh4mBsbewWiJ4lyb5BVadxHA4O03v/b
iYNwTs2AOagym8yDVtS4wcTrL8qTPdWTNaYJCGUkBgXihVFOIS2wbb94BWSB4sRyL6YW6Tf7E/Kb
RPxiMeHlnEMIN0Vo3rYEfLYe1w4N1JhVUwdM4oXfou889wC8iUVwj3qIuYzeqDYBCVIyMNghErHS
IWu8EAGI+xCQpkglGZI+1XyfKaRg9m6lNfrOk1OTs01QItAW2NR1tOhEe3dYpThJ952uR0WdpPUm
Mpa3ZvV70/O4NFhhjy/N2rOxxNut5RdmcRax7iKqd5MXQ9znJ/iP7HFt5DGreoC49naC5Qhnj9PZ
8SbY9tu65jVZysRJcOQUpQ+thTrokDwHB4GnPAySKW/ZQID87+5N5NbLQVp7lYZFHqDZBg50q+5u
3XcPPGWIs7aFWFBxHiJaxnWAUwks10rlrhh5n84m/6z2nWMbiedM238bmTtoz/YFBl/uMyhPwjCe
CCWaHnGTyWp7uK1xiGxQamgp0WrRgoUvtAeZ9+uGHlw43fT69sF+DMj6ff90gjirB2x9NXmvvJgV
c83tD1ZVJBpBmTo0lnqixZqyMo9OYlgSRGnnM12uGporoja5bHk/bIwjWe63lmtgJL8mP3qBS2Sj
a3CtPAi8V3Mxmqu6tapNXp8lyxOdJQhLQ9j6+hC9U7NA/FrO0DsNFnK2NcFo2ocPpUx8HlitnDYq
0NpHzMDfWq9T+WPLctzaUB0sIWvE0gQy7lltzlGT8syn1ApH8LjO1okBxr4AGS0p8X0U9BQOYnLU
jSaPxIaXdTjc9j+yTuZ3/1eI55cu2lw8Z4pQjyaOQXxhsv7lnW7HgVfUODFSgNm2MGE4kSzVM73b
JTmGZPSTyKlr5XEY8qmo7H9kNTji8ixTui286UTaz99kps1Al6M9K5KMVHH9klTxZdsGaxfZ/lUP
S24xPqOj1dn79kibDcHkAd6lcUX+JFClIutSDiRrXG+GJ1MLvxEDT5AYK1icKsWKN3a/POWMDh54
xiipkVi2KnCal60Mg7atp+ValHLXW2RCSjfk2vmvzvFN40elDK2daMf7H/KyS+i1QsApnxJtz8D4
GHMTRYUvj9MigDwOCPJsrE3LS7bgqrV4ti0fj4x9Dxa5XfQslPIcKhUsShEbwDy1rMe2NINq1cOd
wUwFgwqSWjyFWi8+vZ8k7Do/koiwUUGvimxEqSIclf9eqXq9812w1evCH/QsvZ447AAOpZTXYcd/
/CVErQIpQUUPn0HPhisAeaPO1N9dOaCcHdWoJZANRyavMb+1MC/jWN1pw0j8ykyC91J8XwHhwCHf
Acc1iOBbgjT7QhSzxHc+OlpJvoMyrvd6XlhTfu3geI9fv8xw4ozfPQs0GDEyFXO1naUfYmdx/Rj2
Qitf2cc4cRIzi0c1SjAU+3bJgx2FME5HHVQJzWzyH/1dN8EoRk5pJvj3/cHxt27LbEzG94y++WmC
SHawdOeazsQ4eiEeG85wcHMXwLdj9xCb+JauGas185Hr0jvZRGDbonEL/Lz+epnE1TA17Y+inpSb
pMPz4iCNo2yhMofKYVS/u2J3zEAKfjahdXDyQ0mLQm5+sej6358fNqxZnD+5JzXdEvY44hyKO0Nb
OhlXwJ9yVvbPFHGMxOcGcCH7INZz4ESUKAWWOQwDSEpUxwwqmAGg57/Lrrj7S9/MJ5QQZSWcquZ4
VDFTxc2+3dLIfMIVgp5iir8JuxDw96lRzQTPdZv6I/etxDBAQJ2VbSUd52sQedFgXIIUFTMB9Zm4
Lq5u9cquJO1wUeO1dJwepjVCAbu+BnuloqlMKwPpXfMVobTD2eAFQVi4pIMbm6Q1tILjTVmxFjR/
/w+7dxW4voBKwCDpvetOaGw/3fN992vwvYtlJ3sn2SSAu1j229hlb5/t/yxrmPonVgqS5Zm9k/o+
8BsB9+F0FsTglDw8s7eQMT91r4xeXbS2f0LdHEjnWahiwByQyrEW1IjBJKGi7CaLGk+U3D//WMis
aBfPx8KzRSdmPW3ajI+dPJ+INzsxFlTbFone2/2Uo/7b5JCMSL5dCOIYIpU3181CU82XEcu4BQcN
iQ/Hr1P3QpRGhj/2SVzg3bMiFuTJ/ihPsQXyX76vJsH1tIHNEIcChPSnqvRM77lv9VcC5tL/yoyK
arisolYnI9pUIW2WwI4efTqtX0HhnaPBpktZ/8mw8mZ+7wp0xFbTWT9asygXSv7ijb75JpWDuZ/C
XCy0MRRnydmgodKsKCEc094tFFW13PABFKHdZH6HhZABrdjjxV6ccDJfy01c5BX4LCKT1Kyw/zVx
GwLPgni8ytYfAWodWdZDYzfrGSFF3KwsD03bfGfGWevRHmSA/H4jnc9xw9XlZOctZdy7fxUCo1LI
3r1g6oC3eKVeaDDSgwTZZcmwMRvxlCf3WEz+5r+TFYAmiyMHrgKfswrE3lTPik0p5tZMh1mJxTbp
shVmtC61I4Tr4hMRiW9kJVS0j+d4wdINfdMFq0VDMt0C9nMyTpQQcf11KZm5l2hFnJYkc69Q3xyg
+W6CsGDfLnYLSSJclmNLzs5GphgHnFVZmmsCurd/3YeehcgV4PrbH+CZmzHPsFD8JJFz0qF2BYnl
Nyswt2jMl8HfAI+S6ZCYDOlzf3/sk/uDPz4rHr6aVDlXD+2gtEpAldNUa9bSjxtymRmmomqGscqh
9A3vIDVfYAmOJ3xBjOH3k4pGjdiyxUjTYKj600ZxMEljQqzuDCCuLy3bvp1GqaVOdCZ7jZETy/oZ
6de/lbPEH4snvXEyh/p26BXKdUDp/YaKHQrOHiDMJME0D6mG8u2AsHX950k/8VRheZ2lWuVsa1P7
YzqdOhveYDBlN42xrmEY/Cj1jjqZimYmvIPEsDMtu9nAQhKigQAmkgWb26lgdJbCw1tpXK0fF37w
LuX6xQ9d+Zx70WfIOAv91U+MBo12joHrFB6O/XHLNQohcJ07dBlvpbD+RQ1usMcSz3lOSfCB4XZv
2tBzKsPF19BlLMCtJORHxngw4CU8QToHK//uA5++v1tPoUpHFjeN3GuqVlAmiu8mRW8PStzQXoxj
EyUb+qcGBlrC/4WNjDPUpYHRsGhABnibnMDfj/z1OZhTyfqmABP+NjdllU5IKTVVAN0WdCZdse03
C/jLw2oKDcaHxAfzwk4MZC5zN6xY1Mfj89ZXwYnjYk/y+SayaclbU0kiGlt7uqcMPZ4UHxezWOfK
gax73UsrbsAnYzT6i+htRKyoZ1WyEjW36Pg5LSAR+YcyRahl1nV/Nay87Dja1NPgh+/8DeG8elBG
LbjzsLdis0aqdWaxfURl1rbO8y53C1C/W7orBrBSX3IuXlXrBN7eLQxEpL0oqAc1zigFu29P4Qx+
ByD5oU0/Z0CjVD/s9/mmDml49a+wMRwxjskfQwYmRFbMqRabVcmG3uSXh2T3EyWKuLYHsXE50i/3
vvhisH28/ZsT8xA+JDLWnCNxoYKMb8KWA/9RJO3hYo3DR1Lm0mcVBAh0fO4cE77yeTdnkvH4Xd7+
YC3CTck7iUa6zQLt+IQ6SxtW+AUGDovQHUZQr1L7Z/WNQEI+u1KiEY76cvrSXjRoPflXDa2iLNtB
ULCy4VNUmpmru/Agyl8Bn5BMLN/ttCfFWfC0+9aokkR9H3mLdwOCUOBaTvYlU4YU0pFaGkEGXoCT
pTSzoCww0cPR9LOerqye4VyDXZr9hYcikbVQ6swrGX90JcQyKEJuh5mLh3AJH5rora1LJY3/+gDb
BTMOmRV3c5cu2wZoRxWk9UeQ5SzFqXIlmqUG4uCrVybPNwFjnAS5iffqmLK/6P4EQfa6O1XQauHJ
ubor43Ek26TdGIJySTFLXGzQBYWmd2MqzbQlX6VnegmRqi0k9hsfcUMjWzstHjeZIq8KBNHq2MWL
4dzaNCJ1LEKvTpRRi8NPHByuX+HPrsTAv1FMjRc8QPEH6Dtlt+i63C/U7pHfb7ETxLut7EUMJH2o
Jmvl2zSPQF/hoE1GQXuE+nw/6J5GInBhC1mKzgCCdLPL9F7QhNq7/du9sSnd45MyUZXOH2S3z9OC
hWuZEvYeSvG7xN6z8EevjlcpCxOpB2BOr3T5rxBcaimnRmTuzjfw5yncvQ58isTdJwD9aI/ZIxml
0LEbkVfSfIw8lweQCXTo8sMwS9l/yySNdRQgwjHjtutcvEb7XHtg6/bcAj8v7euFUJn75GiNX6vk
BC+4mEZDbxHrU3lDt866sf1KAHWHl6aQfa8uabmSALYiyG9d492GZUtN7hrtxVImCWgktYpspUmg
BDf+5v8dVGzUFUGEsNp86kpnOgcMeb2GF01mg0A3R5gyCkV7I1dTF3NjCEFqYYMInh2CoQRwNL4r
6dzS9UTQVAnX7iqZUJ0qu1QyyHKlCgCu/fIcXXF8A0/zeQwHHQothNMBqFzj5BXulq16gUjjUqrH
1cRVg0dfLXADnjC1UBWOuIX3RFKom1Dahk84Qx/wT4676DtsNxyqWpEvNv3NvvfyZQyYugfOAAIs
8jzBsdlnIE/anqm1d0asnTb6uRA/lhI9xacmPi2y/sO3xmGsyKuEPDFvEpOnH31K2HaAhLLhz7MV
Z1r22QLp7j153m75nciZPjJfsN3kn0SpjvRYN+WNnWVXb8A1w3T8cCGnY4SPjLhvPGeinvLr47Ih
wAwVf3wxQ0uYBtasE8fDTqlNBAeXVLiqlLbTFYda/G9IBYuXiDU3+qsI04I0ema4x7RhXrpZgyKD
anjP+qMWk/COlk3dw+qMtBJC5EAIe/uWmxoxZxlImHvv1rLIstcLUOb4f3lIyoxuJ+z2CAV5keWw
/nn3Tq/U3N9F/rWu5q9s9z2INwFAaieZy3l2V2hH2ocdb/EjMI6Eeg6L3VoxpAvkWJgAEg145Xz8
luSh8g8bZRil3SH0Qo+V+wtjo1V9nhrj5B8YxKE9NvafoUg2amGza2XexMc0MJg1gx6vX1c8qEFW
cEaIKOpPUEqXhSQvKEBOWbI6lofCAB5z7Xz0ORDFcpBN49CHMRy6HERnMKV+IYRPmtbKaK/6vKXV
HRUdag0pXUki3jeSiTTUBi1R630njgkYq0HB4X8+Z63d24Y58fpVhFmYMUoVPAJIgl91cybk5SEF
CGsAl7xJqJkEvDAucxhR8H0Aqjdv7dzoduRJtWcQkdOi4+kzaY0FHwcCYRkeJbMJiBmbpLgWw8CO
e+VcSvTWLv0jh7vc4Jugp9D4uccLLT5lNTZ5xLgvG0+CIOSgwStA7pGzrvfNvDQTlSEdcqVyQb/E
9n5CKUbaCrTRUGOriv5/p8tHfgt0yT5K7kdtEiYB4pH007e9ELEuIP4PBs+UUE81oiMiUucN3HJ3
sGTHpR+z/on3M/t3//xBD85MIu5ySOzxmv4EmmymMjtuZCuOKOpBlr2lq+PTsrzE4WBSmcJBWYG6
NTTQa+PeLxbIKVJZ2FR3Rupkz523CTjrDG2Ll43NMPxdDMzGZCp7Q4DHGbS9vWBtNxOzQ0Zvbys8
9O3YABAY8bmqwx5q5MxNrFTdM6GJNT4WhQ48HU084K8ZmvzzBgWhH7R77mQdgzvbuhRuMmei5nF9
xiKq7JRCkJVzQzZCwSNhc6dZLBZ36ywmmEa6UY5bdZAqQIlwZr+i2tGr63IfzJd5rkO7SlKnwIW1
YCj0mM4kzWHaiuUGikS71LPh4wMgb6C6i6otVG0UKw40AlutTYGerkJN9fZ53zVc8ve+gQncPUBu
YAtPBTL9ReOnal69cez+RrFCIojcnOlQB3DOlYARbygtf+fIQQU6WfKtvZygCiDCFwOCXb//Nzcr
XScNTk3jjXFBYK3QCexSujJ2kUf1mRXqSfnpHaH6I/1VCNT40xjdv9CP7O8PiB8OX61W3Eqh1vRI
Zb9aLsF2Rnp/GIYF3nbaagoNeTo4K1tXznamlq/potA4xUHfgi2wfSJugM8cXnPetEIlm14K44+f
UFQCON4Uh45gw+a4CrsBOVMdCHYP+JEufiPKV5euX1SXp5nGLOtK684q/+f2dmV/c0Pex9hjry8i
aUM6WP3CCCWzo0nU82zw65HNheGHeIxAEgs7MmE1ZcbF5wPBEaPEJPtMlvRL0ibpx4l2ZDeuIb9k
9qHw/exSkgP9961Jd9cN/x6IbUmWZRkCH6nV9lijiHEdL217VoC/czq+cylG62zwbAbUgxD2IG/D
dQ3ZyBCflEOt3B5zfb06RulQMr8JQ3i9UjTSxJ6x9MPraibZUWj83hWOS/SJVjsXtMEeJ6KKJBPg
gdUdtLyXzGSSdDj2/3ugfHn7OtXYTh2+5B5oDZiYFxDDqNT6qFOzG3rwMDzdQLj4RrBSV0q74kVZ
Mc8sEQWRLb/7nrJsun344gXxwMq2TaaeDDX8Iru9UFdw1SKkV09AUACSGsmQFVWznrOzTf4eZxsD
9EcTMpWXydpEa5/sRQUDitRjcjoVkjJJgwje1YJeRTlpA+ATtvY3UDxJHUfexkTW8X73XnmYOwC8
/VJCpuJBx9wBMgKr4/FlPeAQj/rXPiKSP+BU20LcvW2tp2PnFZNzyOSHm+Ex/1ZQahUpDncsGptz
xwKmF+5hpqhy5Ag/SHJqUH2BzOdqL6ao2PqlOXXDH5QrtCRTZwCRS4Bfs8RkCDJv+HnXIa9qch/a
7kP/muBRUotZc8bodDTbx5N9dlL6agITQds1n+dj3In+vMblAtyUAvJqaPNbG1Hjg+6+d92W22qY
onBo4njBKKS2KWTLhqKJ+rHAs25yloSHNjUweH888E8KLXG7Qnb6rQtpHicW4a0refyz/jTuxomO
7CEHk7nbFj/etxnc4uWMQVj4BPqA0lbh0eJZg+cny5TEESpSqGOTVY1Az+ufYF1mV45OnOud3ssn
Y+hNuj1u/UGFqrEq7yS5uVTQLL2ZI8zLmfMKkY2BwWy4PICEOfG5X/KROMbI9dJJ8/APZsaAN19N
jcKmymcw+hzQ5b/bZCXEV7VeLKhxguLBHe563WZb04OpRY/WCClh7mSbA2A/fNL3M/9eMsNk6cge
Yv+0/4pxQD74RkSLugq1S3Q5HQ573NAZ+TjxoWBklqLuReK0lUrLpT8maU3zBm45mvkriW+3w52l
HQaxQUw4NqQxIwWNPOXfr6UPSo+EngZJ/V3zWPF/RNJ+v8VoWAgGqzAwyTURDOLQrwNlrIjDOGeW
ZZcuOIgqk7GiUpMPwdmL2gEBgMNw82CIFzCC19DxfVneF15lGgiMJRUswNdF//mTcVEHsm+NT7A6
f4w0T3K2ZtLRzLZJwWxlXy951/WLhzSAyy+Wnhi6atN+xu1i5mT3jEr8P/HQyqr/ZSAsSqEFTjry
t7TP+IHF1gcHhpDC94GxOkqAHI4+s+YybBo+B73t7xH+ezwSmf2Kb169V1OObnYLi6y3MsCnTaoe
ivU4nMrVq5bfFfg5VsYHOw+joogEY/YhGdFrYGCkIs1oKrUWFsMmWdo/o9jNwtRh9Tz0vD8YvHk6
1Ba7SBYodmquWo7C7x9PsEYYqeN7SOcZ5hWsgjEHD441Ilt0lkEePpkjVQTx2+W+n4WIK03zvlMk
20cae2zayLYyCwDT1B4KzLRbgFaAl0xlRRjGWlUg1sgYyYne+ic42KikLMeEhjOlg+7TpqOBeKhk
2OhItcvfLRRi/AlgmeHCqVpWmqGOn2Saw1OeWW8+3BFM68evoVGaXMV5DXISs0PYqVsOZyg/b9fs
G26t1D0yIFDV4KmI1VVup+MtYJcdraBs2o3uk/Tz28DMOC/0Df1EeoKXpTSXVdQV9gdsO/9CGIqe
xC7NtbPYB8RAuTea8Rpov+/vROzPa2ThzwKafx7+z2tlJ8RHbhUfn6Z40/pxUL/6GBhyByONtCQH
yNJ8krjYbZJowjrrTIO2jY0NGYiiMY5Q3NxGXqMDgE4u+f0KM3jkNPrazzP4ofZ8BVLFGzdVmMi2
WIHDVsctS+p6jevLvul9OBCuxDcxum2Wt0Vl+SYCxiTvi9V0IYeQM59OXZYy9FgJJ1tQZJHF1EoV
hsQ3Y8t/udmk4VuYEWTVAN1MaksdHnIcgg05NEMNBs8bfKvvzs1OPEyBKWdDmadpum8CnoPkuDyt
Mq4ODlICykOPas3R43ILS4ulttwEBAXYv97GiCrZx83G4DFehDIamMvSw2nmLr7vRpjLt8iCC1fq
CqVMueBsI5vNWLXGXh67394Mwiho5neWCgHT6rUhB5qU3x8Axc1VJ1B6nT/8aG5IS8I6xgFsyHE+
MjouiQwMEL6YaLEfvIwTBaXgSz3s7uj3R+Av0s7J9H+zef2ctbD/opdec8XevCgQOX73egNRLQDc
xtY06Nlnfqk7p5Qs/L1HyKoqe487kN933gqqSMXENGBF85kfRYATyBAf5eimhT098VZL6LDn4yx0
mONXeLbOPG8anccmJSYOxV0hJ++BgKnHtXq5Etrxn9/h24gTAI7qSi/cEsrfOE4fJgB9dCv0ZA8x
4ERwaPDRs/fFO5y6ue5jtvqWdH7iNlpSp5XSnYNqhLw8OPXCDFq94HSoF6yOvoUrplgM6wC/RkfP
XsrXCzVxKSPtHDBI3l1kxOVs+hR1UvrUVGQmAjXHgqA12UVznuW9+gx9ttIzZaswT6YLlcwo0brf
G21oBpacHcJjCcHra5IERp6kKsnr1JQM5tc0/3oo+VStYirIHh+F5oAzFtvTM5RE+TJjQdhVs7yB
h3vbga73pmllRt+2c0htiiUEU1vY1mztGhKRFB1N1ZtwFtWJ82D5aqR+1SqZY+O9efvN1n7JwXd+
J1THFpUV5fNNjLKEKtIPaUgOPR2Lv7V3RgP80hW+HhL/EhtjzGJM39Sn3le24Q3Obx2VMV3XGBs1
+q24O6JH5qz1uPC5X4jaShMmlVlrFiD07mQanprZr/7crHMliOs9BWirvNohx8LZ0uRD+IaD7sdU
nYa+zhyuhxL4JM8OqSSqXZ6dhng4n7hRU25BVmplFfNGY/S0Ai515SMTacVP0n6xd1yT5UO1qmqk
TwhxXfp+Dbnw6aj5Tk/LY/3ERGi29x4b5Jex+p7tK2XMKnt+mCvGeGS7/CAfuUXRJDSfPd0HIQK/
U1wGlEU/3yMd1D+NhePTxTnfFPU1sW6D0B+UyEzz71RlX6dhnkfDkSkQR5m9FI1rS+Iw6c1GLC75
t/fXUYZT/iRnJG6NytG7DIaOYWm0mhMnbzZ5I3mgIGMflZ3r5Z0FIORH+xxB2HDl3kRExex34NhM
PnM4H+2M/48XxCr8R/at5qlatvTa0VjefgU5kws2MCQenYu9CDz7NV3QP48dozywud8A3F4gjdhs
EHMQVyQtpjcxIgCWnYnnpPBZaGAcENrc+uFL7j0QWCyHTH/xe6t4lU029OfgyJyqErag0fyxmhnj
PFNjG60Oqjn8VfVY/BcfwG3x77BaDHpth0oQQPeARFa4O4bvw9N/aqmAI+Nf8wAWpJf/+yLjNOzi
BfmjgCfifBQQOSYIWzNfd8fque94yL2H6EEu4mPUu5Ewt5WuZvuyDS+fVn/SxiPfSHJoE4ssdyMP
cK9AhX4z2SikI2IKBRrcQUTqhrwpla1ww3acUFQ+5M05nIce7uta8abNdKEq11XwFTl93l9oDm/d
PTBqQ1N8EBVZbculTGB8oTJjkzwPN9UZqI3c3cgN74Sv4im6Atm+RmV9clKvQc0bfB6+CxDeBpdY
4dzu7fVcPw9JqsnOVDHsK/5RCn2MWaepSz6adjInu1jBF2apvsS7XVQ69KQmxMrsjBeUCkKivwpK
dqCHIzOxznI043d5i55nKfHkaf5XGeXkeYzIyBv1Qdx0Huc2qgIqUA/usugwwCGPVZVV0TrrsIIw
F4/lmZW6c29qRW254CabGFZ50ahISwKL8qfj8kPeqC5pXZGY5V6MJcX58n7YCgO8Ej3U/P2PfZMG
QZgE8Mhn3i7MUPFpZINTo/bOeNoeSMMoIGOAVgM/zrdjViv6DLCYoNsJD7xnZOJ0MfRRotw12N/n
b4ZmbcDYP0I0bFd90n/fJXW2FR9023m+K/BPW0j+3KO72YB9OobkyQ2u1RE0HrLe0jUpUVMqtmZU
EymVUB+gwN2OR3IYsSVtiJ69oUpYTHHjBdcNmrR8oWB1EX/YnjMhJvgoL69Eq0/c2vv8+2n2wUcv
iYNy4pras6MqVeq/CMZWLJlPwEfKsi0jGjAPO7n9cSUCDbWD1xTlBmiVO63gCWJq96gbQYoZx7jN
kJOW26RkLhuqnRTOa+hfQGqj4lnO117exgPjFY0z4j/X88eOhMz3uSkXwz7yFHV4mC6w1BjCq6Tz
ja/F7IBOYE29nXsvOha9QIIc8E15dlh+rnzbu3ls4O9OAn896SUAEz465OeXxRmIGsw+Mas+qhwm
7l6pnmur8JyxTxuh4BMp2QCP6RXOExTqY7nZ3fHGhQmG+CH5VaJtBmLQOUynyAg4Hg9BbyX9THU9
AB0NmB1D6813wjX/A9AZungJjOm5X4fY/TbIBtgqwvSiyA1/RVrxJGoQFx4/aUIL6UFBSokBGNfH
DqUfN39mqNjKiSJHeX6Tp4wEfi29jPxkYP5Vdn+3bXSvyC5VeqVfvcKhNbp1E3K3/bGLVwatsbEx
hqgTchdekZF9+s3qE4/oiH/f3oxqSf/0jQ0X0RC/QAjUWmJ+ZOscGud4IdKNcxpAE0i9YcmglIkr
C1alO1aOak9ECnWJfaPbbt4QwaYXEwpehmQ72X0layeGdVh1WUPEZmXVewKkP2yNXt0HcWa3YqpN
VtatcjP6rLSLUq/JIG6DGmFQuon/3tGshi0KVKnuGBSEYU1Rh2DOOocaWKflvJjBm7TfUkGJhX1x
fyWi7PF+SE678vi/5GruIN3Hpy4iDd1yF5vRlfx9b0iku/iUq5DpCrloyqS71NOdzx4JzV5gDEuU
FP7tBIDd4kW3591lLziWf4VIkQSYCcc3Yxj5/BGHNCgsPHXKoWmIe86AvZ7rkCcJqdsffye6vyBE
OtLt6P5I8WiFo47xdzNQAHCcCnvNjJ7JN6SSIJFe/tcjBI2F9F9ELZOQgEji4ibLq69C2IET8CUn
4o6aG+Q56zvMvI4Cno+FPnyherb303T5Y7eptTBBGu0hsAf2eF9faGQHxQR28oMve+IQevH/ZSWG
8VoAdjf85pli97VZpjD1jmTCtYG4q9VYc1blCgmXPIfIWMeQY90u/9Lm5kerVbVWdqS4Q6k/XXhk
0d3i1LH74nKj0C6DoVaNY/LMNcvatwk6wg9SQYa3eXgm9t0wWonujL/d0d/miire1R+VQxLUBacB
4nz0n1j+/VkkvEVGi1WUIP8SxsjTlv18yUiRTQ15EOHYOaMCGFpmJoHtQvu2jyGwqIqWIYUHbYdi
ocaZLdp023IB70r68dHqUra50Kc0+YxSujLNwYO4r9PnDEivHLbtVTLEN5C7Lqd+GjHFT6dDsXTp
hlp5GGaka2MVGleZqO+6gOj63K8YAqfpMve/OHG/SNgiy4v7ENyLKRwqaddgtfg8mXokxlWz2Hmg
ufrll0Tmbko5i/IbyqhaKQFCPkZa3mVWcfv/OhF0VJMTT5gUHyIV79A+bbPFOd/vTygicBaFFlSI
icHJiztHRVcPxBEMy60XTxIt34OAW1X4snZAEpX8HzT0RmmyrQjQ1z1kmJBQbFXpgD119sp3A/tb
yV6mtY8gUYargkxmgl7UWWY3WoN81hNYG2Cp2Jfbp4PpjgCVr4l/SAlpdAjurYxwRb9f4AwZ0y52
H0m93Ma0dJoRswM6tUSoOQSO54gKe1bheuj+tAU53QdoEmLIl+/1d3WvtGK+94SVKHYgdMDn4TFc
drH1j4puxLvF/enTTU5Uf+1hQWcxozAwTwCJAfP4ZbzsQLETWngLJe0GOU31xVCxJ2WuOZ+EjlKV
8aadpcIoYU2unK2ObsZ7CHuHPAwSCLb2LBBwdgFNU0KZ8fjGwUprv+M6/wwAUPurVvIFS9GYodwI
Bm24xu7nkEQQAiMkro21L+dXrKPOZxY0WWCvDrK5NHgJt4u1Fzp+fW5Ain8fmRylYdFGIXrXiuMT
3EmmoWfZr9M4LKNwnwbzqapcvRk0XYVbIR5RcSxNjkGN78jusE+1Ma125KvwkHqfl7oXDu4acQXF
786d8UdjaZIetwmMrhLfGCF2P9o8BsbGfLlj9cc8tLD8PbxAhqfYsUPmClw+humA4/5hbCZ05qEa
ub33DX+YNcNoWXR1BxmlhBpsJ9WR7sV7UCViZM59DQc9b7i+Z9xRiOXxaTGVTNpk+xQKKGBByz0S
vfIqZdlux3niX9uI/U4OBRuf+WBwu5Db6XfJ1wUaBQ/Msbh9AWxFLlVypg5SP3aqRvEcoiUkl5gX
3bkj0eyiffAldJKYgdxR5iZqZ4UaWQMMpbBJnZgzdWKqiAzccP5PGcU/SVLK0/Qkw2RyxemsNwt/
XTAU8u9shQkGEv6VcvQOB5fEYsq2UyIIvAc4XdJx6KABQggFheyP0bmXYTk0k4QoTiOpnxViU1A6
Zoskv9Rs9QdakJuqnSncI+xaztf5EeHwREbMfm89+bfFYJGg232RchIzHsXmTYpS0/vElM3cglJQ
S+rSiOXd+lQuJo5D9CQ1Kfh3JH+SnrRItOwd0VTejR6p4XTUCvqNBnmraeZKPRA+ag58F65V+zCC
E/+M6feN+waVJgG82Sy23o0a/Gx+rrfAJh03rzv9aUCKQh6EAQQ/CJVBZVxtpgMPlQU1LBLgWXnT
hxl7eyt2NZ+cbj28VfAxgMpMLuwnDYDCWxToRPWeIkqjlsMnQgqgwKQk3AMxzPHlUKM750KuU+XW
tK8Xr2Ss2LWi+7+27uKtbyAitHNP7P1x8h+5uWaDMc/YT34HRKJ4hzUbvi0zehi0PGfRL7wA4QOU
y5ipX7p/8hiKqO6qhpgPZj5k/HqddhNlgsPZ3PKuE+2yr4qKwV09D9upSda7Gfkj5TeEVmBa6asg
SyEeyAS4U2YP/uzLo0caceoGP90TWiTBneylU07ML7EbXKeNFYimI+Mnkly7yXBcxGyzcDHondg1
emsOnPZGmQEm78jT2S/bOwWfRdU5y66UALGC3siKfSDtY56UBqh0eWEwBc7yXgQBXz6dXUJ8Yz00
NxsJbddkRRS4kpZfUFTOnvp+Kseb2M9zv8jB/5Ud8NEu2eRiHS+UR6YxlWpucmhGQvDEnuoAR3X8
WPTj9PjgomA8O4xrpd6f+OkSCGhWfI9F1DEEotrCBICaOqPSmUvaJXYm/wYswcTh7OV38tmZGTNO
6Y4gMQ1qvNG1hIK0ONp+Ty/u3gwKu3YRMCyBMxrVT/avHxTmwSBS1mt1AiZPoRYF62q2yY3vCD7X
TwxJcFNIInmfIM4VIME9AiSyQO2nEkbVShKw+hYkVtakWutf+GtCmr2is5XNUktE1toF7iMdOohH
faHdj6i9N9B3m7VYmCIyxfIjHE5LO8UC9F5lZ1U+zetTXAEBqlUl4L0vhZvbYFfqWs0lPPGzYKcP
c8ezfg555HpMgP18kxrw3i7yeAM0TQ8LaAXbsxqGJL1WdqXUWZ5Hd5gJyuDkZwE7/AnOPtjKPqPV
VWPoiHGILw5/Dd001ttJ8+rci/dvUiHok1hstPb8eTZL40oxq40AXeb4GZUmeVChPG5jVi0flbRY
p3QO6boy4VlLj0ZnRWUa4LT0gAXUYlhlDfZOUuP5foLPdI478Gs+ANfNK8i1bCmzV7eoyMTCsMYR
3vjKij1lt8oFC/ts/mWhW1nAvisHMvTBpouTq/NYkcNvfWRjWZ8h3lIqgAgCwMtt3mTmFJD3WR/i
i1AEScNo0rcnYCN3DRbWEzUG48fOwEpXLFx9WKZNs/7qP8qJ+S+JZmY5FfzGjoPp8sqxAeAhQtpH
rmS9ggc+JLiey3oMTFLYKOrQCsmckGYDQqZG9uINrD74G5J+yDSHz8a5ut6tArIjKW5XwoIKji28
8+Ft8iQywKb8qTiV7QaELJY+ESaL3+GbVKFmRtgXfF177cSqWy8gLxpHghRMV5a2YB7KqjNXpqK9
DYBNdk0iV+Gjutu8k46Z+Si246CAG1fV743dosCCaQ12PtzFiAhq1SRth6daELXzp4haWgL17A+f
RiV5X7uWj/vHbLUrMMrY/sLmk0hRI/xihzZFfwFs6e+yHI/nKz0okFG7vlalKyapS26UVcv+fG8D
bR0okgAGn11DIGb/3LWIN9SFmJmsKSWRcCwRZKOt+xEva6iEWRcT1RJuNzvRpC9AEWpAN7jtDIbX
PMVl+3PJN5ONhePMhnef/N7SzeXZ1a3cV4eaAWSssgBsJSwbQkrhbJdtmaAh92WnalhDSuDkNBSa
HemfhJZ4aXhxK+Od20dnAzilw8GcRFKV6uKpzT9Rc930y/gUOvqDTq8SirC5VfNiEXX4Yyx6e0Gz
z5znN/c6UgjbcIru/G5hxn1hJoHP7IPvJSEHVMrqGWwV5NitNLdrTBsFxraoHZ+QBRgFi0tb5EAl
QW5FJqa8gxisFabUnyUDIjNcuIoviECkKZJKf5IpVPuxvuPcbgL+rXQvNKazFhQ4B2/vnSK/eBOa
DY9YCvcbCrb5QVzl368J889rIIEWDwCy28vkH4W4BY1rMPweUwthPTObVfFMmUWsI32N7QC/UqRN
w0iv/uX6WOm2qDsHg9PO9dL1ZFgCkWkpcb1jdpDLYe7zP5LrBNMvnLZbrUfqYueTZKFtFCXpaolw
AZT7uvmPsLhxNNJTNzNMZlZ7bVhwM7LckaohI0p1WiEou3BGFFKpr/dmei3tMDYxYEqq+Lf/cf8X
iLqiWOVYfDoKeOBhOFBZFN0+rImtP4TjSbZHPFDLkJDIwR2kVKfLqUwlWRdlAPRF/yBIcNl+d8xm
SO4Yg8DluonAZ9o4Yi6IEPV02zEl/lxb9iudfsESpkYZZ92DqoQUAczJ73kgR5ojCokrKAErCOfm
zhuvryWXHCVr+KTuDSNpwqZCTlbv5GzVKzWrQ5lMw598d8k+Aqf/XbusLCXVvfHqSlYESv0lu58N
dTgNGIj27qe3Vmbw7H8tG6soHGqKjrnBTgWdXOVvi/P6gKQPZOI8MzZThXrakK4/QixlipALiFtt
olM9apJ8XaILByEOGOf3Wh1+gSXcFSaWoA/iQ3x1c4w+3VnwIRoIAozfuOiWVnb+d4WIe4GRcvsh
xKKJlZ7bYznDmXZLWVrkxrCcd6NDdyuLDGvyoT1cA93PJVHHHxRA4nRGePq2VFKxQIHJNAW4SMrh
LrMqHvqGxkdAI1QyDzd4gR8q4uFIV/cEZkNygJP0NLI0blVWhoFM6rGuKCwpQqh/VMBwOyG92lL+
ZvUtQv6E36qg+0p7VyGXvHSzdvMbsJmmDUjk1nt30/9GPTmL9oO3KMBCB2gPw+HeAL/NmL/pxmQ+
XDYYAmlkM9MuKjLCPaPeuKx8AYnOFDJu6idpb2SjyO/fo6a1/6Ccqbawk1lJ5XEly0X4A7DtK+fB
0KIRmJNIgBmQ2rs/BUp3isuUJvsp/fPBD4lOXc+wGtkXjlu0wel9vaR8WmRYlzeZxQupapHJ9DSN
dENJL7nTL+Nc9kyiUy1hwH7L3AKuaaA84DR+HYTUSQAjd2mlaLSJ8jaxqRfNiw87NOBVGibcNEfZ
uDfOvylMJxuQTECGUddSHZmtkOASEfW9tQ/1oyDNfPPhGIqlIRsX4YFs8UEiGm0etu+puTP3Wpko
8J1BZIrVWC0Iqr8djm1I4Y06JcNAXC7+Xgi8QqhC4gVuXbDclT/7rEjHzUo1ca96tdwEmzvqixyN
IoaI79aG3RYjMDFwWA9BH/+f4kS/SPvJ+gicXIEXMybcG9WaV23DLys7ckIejnY3DuE/RQb2ISIN
Se98fR4dntZzVBlY6dKkMQeh5lKRWlh6efrTjhMCC5fHFYLBXPa7mHzeYRYj6BJYig/rzOUnhVlv
vlPRz3OisjqaZHXByxiJBIgOfC8Z9n/K4e/g4MB5Zlf/M3OtiHsQBXQNVKpgj7S0VdzLPAGGriOZ
ltfUj/qWcX3Kch3mqVsscskzoKYB4WIVor4vtNh89NVwahebAYyVjnU43UHZ89nRVpRfUwKcgA0n
1eYH15sNlp6VedU0NrgOJdF0Zoi878duuTfHBd0EF9jkZK8ujMnDWnNmywoMW4R2p5o0MJyA78kX
A11vuiv+SFBM+Xp+TlHTjQBjA6KVzQ8wbhdyj/WESdNjwZbLLsRnpvyDqaUO/w1kBmDqMSR7BJ+1
t4sM723U2/kLuc+GNG2j32BgVTVbIel7pxXDueSXBIQV9Z79EKxaHZEDs8hTV3z6vQCg3jiqfeuT
+vEixdYDUFi1bSkxNOSBzFn39ViB1wxUYkrM2H3bop+NFyUIU642pxgeKFqVnOLmjAre5RAWmbYi
WDwuOz1aODwNrjmC9mMr/R1oqK8axp/H3CaUt2YqL33J8QQvbxm5uNwCGS4OGGbYIZ3GEdtbBiKC
Fl8+uTlyFYIRckXIY37w4PBdIDBebwX1mX7OH3/a1pohlw2R6Tl6lCvJSkiEKY42IgyGQyO+1da2
AOXzX15NMeXw3a+Mb9bEFSc4L05JIPnMEASuP89rOZU6JWLUbN4ygpro+Yos25FLP3cdSNNHy/TS
UP439nmjMB1zCrcm6c15J2oiRc/4movmKp5XmsLeFsX2FCY9VJq30QxjvGKAWjzcbLmwGM+G3oSF
c3NfLXG4OU2kQgyrqluaXCFa5d20pxErKhqri2TN6zb1tRdsDfFpRBx+bRPk0gQxNK37/EWdT2yU
fssBFbvnqcjGGmLHaEq2S0fRx9ahcgoTquby+gp8uBdY90ZtK03nEnfBjnA7GKIwQ8vLE+azxW0t
9Cr3ZLuyop4r0LPJoMj3fvnYv4nKfIKHDB70tDXlNdDWMiaMNn1OpnTDOWT4SH/rvgXQ3MxZlkmQ
UrNi/qG5CylCuPHeEyUI8109vHhKIobN74nU/1gV/xzFmwn8anmjOlNAlamI+DukNbTjlAvhMWEe
41auJ47iCW9iV35j54SPtkVQLUhMpL9/irCvI06WrOhNGlvh6CGope3ozB7qnd4n5iDfUTVUpAJ2
n/lIqr+A0BJ6q7F2C3rxJYjVzmOh3+hLBSdqMBxmpXsJCWXtJuiCfzFJ3KchAq7g4oLA2TvHGAeA
ta3reslSm6F4GoMGqGKlmaqiJxC2P+8XeoWp3247pzgF68eugH+UhymbXKJiRU5WV7Z5pxDX+ANS
Wo68VogUR4unixDIN4HZGUpn6TzyfphCFMH4JEOblezjOCcExqJX/ECvNIWJuuwBq6caiC8neDmo
0GyzP+nlptfcgvXrAAfqgHcHjZXy6NAp0iCg72sHObMUGleCeyEEiJINnj0LsGAC20Ljj+y3arsL
kungGnPQx6i2G4o3gA0Oe0ifRMUDYf9M87rzI3FJ3gKmpIdTZEDNQNHTSPYwRwy/jQDCWPVBCn21
RL/cSy7ZkuwoaxwlBmytlBNntvIa009r2/cvTje1kyZDJTykSuTwswQgthMlM1LC8Yu935Fvqckw
UK8u0WShOXNj0ThavL4iLUDvskXtfeSaky/RhAbHYcn+yfeixGU01+bagclPCU8wh5GP6cQgEREW
CXrGB2RbKwmFcK2od5L4TR/xQBpKoSPVFp7ADeDWDCqPjJvuToitQVpMzW1oGJ9nLrsFB1faYSnr
gPa3QxwgxlmtcqllzGt5pWP/oinVn1lel7KbTkQOVIoGr3kDhOPt4RmHjiV4+DvnZf+YItFj2syr
a+i+9j1MAygw7CPf3qFkZpvFvgAtZpSfk2q9YBKcYyrM5GnjlLB102ySFCMypte9bkwLtIBM28j2
ZBxfgGSiKA9xLLQx1A6W1XPTzUfpOCtopIrrLxvFyMTBxLe7P/C19KcNCKD1/VL1v0FP9KSAl9B3
Wtn67yk+tb4KgWGB9rBAB03mWlDGc2n7Ewa6Xj9uMa/jJvB9ORbFh18UmXDF2THgxDfjsEEMPWIV
4AG//W1QZ7cvx4yq5fVtBwwRH7JAdasjyjm7p5Zo8mDxTQJxMKHvLaq3sux79TvpTcRi2sMqY8Px
qgbTVgDBldwUhJjka0O5kQeewAW9vODbJ7qK8O7rhIAAfVRpIacFA1xhWKdbfTx4sziVlQzvsyiq
ZZuip7iZmc5qaGzWlTcr6rbOWJ/uHmKlp8SSMCysvDE2YLEHXg+qGzol5wiv+beRX3ahG5gF3Ow9
i7DEwZsdduT8mgTAhhKsctKSbTP14xfNtyxmEPfs4sfTA6h/7LI/aZpdcJxJE8Ihoy0RZvdMK+sC
2/M4lV+uP8MVAKQR99rcJoVqq/KAw8iKZiF+IU7+s1pzUcS5GVkm4oou10pMQ0ZNwdUeVIxXIFWN
GLv4APeUcVp1hPo7xCWRbvZYppYX9c8PcPHZBHkBnqdP27IZobdkZA6SChqvYsW5jQFzIYMja0Me
UWMzL8Y+dnUEIjJpks1wmEJ9+IJ5cc6fzHxOB627/x0fJpfoy7s+Gvz56oFqRv1U6k25TUOYjBCP
Z8bNJpRn3IDZnG9oxaH8DBe7AGzyEJjakifK/YXNCd9PCXYMU4q9rxMokTlI5jXmdBiCICTLL+F0
1rW/TTBD6jq9uI0hsj4dSEvwFf4vBWT7oWkJJgHZrF7wiewo33KuW7IYW4CODkeMPXe28wTu+J8Y
0/adxbi2N8R5uagEmgNGCipHXjR2zZMmbbSYZ22IIGrZmCq1km9Zz/Yh8E2eLfEpnp9R7LA4SLxn
UiML3BhWkPpD3F6su+TGvJ1O9xfjFg/Qd6bK4qSbecv/BVsIXrD2KE752kVENNRTuc60o1hihl5a
wHKlgKp1C87Fe1vnNC4pBIPLaHTmKnFQMQiFRxSy4AJaShinY0T13mL/ieg6BRQWkfFu3a69mPHy
IJdaz6qGh0vmtEgru/C12os+Pv8qf/F/kt6HtyMFfhQSywoxSf5wER9F57tgUvRG5iT5DTYwzEkC
hOeS+Tggpu/JYGRr4SMidp1dcJG8eN7nzztYrZsP469EOn1RPTtqo5+2LmLGfaylCL4ikvJt8zES
vVGixES7XVrrB6a4/A/PM15V8U2aFdHbYCuXlh/rfX9BA+FbckBFz0SM86hRrxKfbHUpSFtTZA51
rxSPQiBwtjeWWRPyJMwm00yC7y2duumq3hIq40nB/9hF8WwQ2NElwiUG23Sx4fZNNBgadeWZsDdP
nbkU9GVP6Y6xirNXIJX6GF8rWBJTVjIxNDiR9DFoAyV4uyFiTpbKyVK1kjIZIy1SAf3ca7yTUg+v
A9qHHVGzOJh+nCMmAZHG1/v8Wg3O7aMuGFK8RoT99FOa+IXcAJMd90D3id7YB/0RROglXoTJqeF0
YxdhFzIRVaN8efQRhzXWCE7iQaVEs+4sGT7ahPBXKlg78gv9jSTM+OFYc1aDNJDSRFwsPRwGrByr
andiDbTe/yzgx9jhR1gpxEQwVE6/p2iqcVWTlRXJBC71viXo90MS+Y7dIbELxcoOh5TaG8KFFDgk
nb6WVrrT90kSPrjyDvvZ8UGMgaWU3+H7GM69vSBS8w61MnhbYB26JFozXO87lw5YZvn9lPMNbxbk
yTmQ1uwTMjajhHNqJqicKvZICwxG0nimEC2GLPd2p2RoPBtMq/GWOUgjRdXMUvg7/nf69vrTk1lR
bBeEoTQol7k3/eXwIKg8am6TVuv62u+7WC+as8p7a6pELNccREZ+zapeqpfQEXQUzTcvl4XkEdLG
nWov0OdY6KM1pJQGx4yfSzjsAnbNkN+D5THjwaFroKqyzOeP1WkHIEFlSutnaZzPGPNhUZM7OpGk
xixNPuAJCFO4m1AlxO46Ukb77yZLfmhiigwlksiZnWvMSSMeCcUL88CVFtm8E7EP+Bk0W789ovMl
Vh7QhhpEUfQRwimYc3Sl9J85vCaaMPCZDs2hFO2OPum/IUilh2HsIk/ZKbGG79840LUw0PBm9zBb
uagnOGnJ2SIdB6k5g7NsCu0U7lYdaxZa8iLeDIjdb9CvoqKU95WwUMuwCT9wwO0wFc/i8TBM3/7r
xwuiePOcLrIvDKf+NEIbae2IhWF7MTAZb9sYPF7w3TILKk17A6OyZABOUUTfoWYZ7c+OTehUTlkb
shQ7kFYr9DDZwALXRyWK78HSrgsWc0zX3pkHIW653S70jlbHl7vpQ7Ln5v58lBZPw46ZvVSLyw4Z
e/xImNxNAUg/+kv20M7iE1Pc/+SzEmxRvulsVJ5uAXDSJ19Sr/EncXOHKPC+nzbHQNMUwHGYnC1B
sHexAnU8xFgtgzJgzQXGDhFO9N0JZ7tXwIrq3WpwIwuVV4s0vTF5Vt0QpvDE6lZdWxSO14sk1m/V
M8JZjXTkRPqDpskIXS62ppvE4xABqbEdlKfolH5yAl7J8MG2/l/+VVxc6BnosEAfu9BUXT8890Ws
oQxpRhxrJz4DspLB2MpvEwrm6rOIowCgxZ35/MsdsmQu3xGuPc8Ts/2A7AUP/nICByr6kiVNTn3m
Semd7ij/KROOjxeZs89x00u6qosDkoLa0cKO+fsLZToqC+ZoybLJJ4zG88OKlDk1CwQfr69zeYyx
NsRIvhSVU4qlvbF6XDJIhg5WX8tMUa6VVbKIXV+huqaUHCWi7hhUxrWVmvg7tfC5mr9pQR0rblli
6xrbaYLw9PJtxSCTC6dXdwIERXa7s4hLOdn6+cP8IsHEqDGQg/2xjLdKjAnicxMSAONliW0Wg1sQ
cs782+6nV7/GnnAXfNtnIK/aelV2sBbBzriqeM5iV3Yw+euUUPGTY7NukAgnBPqtd7lfuTZVtOTx
Tk20r6QimjHRub0jnCtEgyPJMtRKMs1vqwI/lYGZyrF9yENapwFHvbY/6PchYJl5BcKBR5ae9ZWU
5vUiKxuy3+fNUP8e59XYn1ohbPWz/gal+qlBr8dnYzF41dqZ4wrGerHGVW9GdpRJEvoaBqjdk+wG
/xM6ShZnKnyk1Q4zzi80MxqJYpyqU9LlXsN7bpb2CFQWClJ0xrZOpCD4xhcutFd7ZBEifeHyR5mk
nObFkUPBKUf4P1+/h9YXkz3R9pjORZDWGBD7qVdSUFV5KYtNHQifQUGW4xQte9YMgjF1i7W/jH2P
xkFBiNyyxj4QFAiTth/W98qhtj4Nbu/j121eLDVnO0RDQmip8/H5nTKocyj2Ge73OHZu7cMF7a+5
VOFmiLGX+CBzuQdcvXI+kgJALzEh3O+08pYk4m7NX72PRReXHEX8/2lzJmwVNfPZDggUJGue5O0D
gTDGPIh8TGa73YhOQ+HA298XsGBbNYdVAu0xcGbFLrYWGyecMKzUTTrjvFGQg76Zxx5GanIeJIof
4+1hP/x28VfI6oo53YdyqV/RYyEDh2WKm8dm6GJsUQnU8bS284rCKfNfpXuJwD24FC/kN7uzAB4I
7ZYawJCvc80MFkXASrpy+X6r2p8orpHATeHllJDy9tA6Tc+QISXvNGdn7KKQKpQKinJ7aak+Kxve
kCmGIaLIy3HeE3tn3qB7itjuE7SiUHQ7ou6Q9H51AdtWF52aNJ4J77HH/uak3ArKqGY2dQcXaAF/
S8sVXWdUfgCv2nr/+P9gAnmjmB/UWbsrsB7kyQE0EMgxjOb5+BZNc2vBTpjGbElt3PJ+YBLzkkUy
LSZtR/x4lqDEAE/Nbto46PT0QdiiYx5Rn4O3yBHkrtUCOD3yqRoKCsNDOHYZBLnyrovCRR5ojjIW
QuUTS5FfDS8NT8rtqprL9OQutURDFRhI1YJf4vhheoiw2F49avuv+vyjPNvELpS3AANAyzauREgr
d6EoYFSj8tr89N3Zn27elFUjgaG1WfKdhKMZbRjbfjYZNraaiFp67IlC9ucaFHfHyXfGw+b7CUGt
UcKlz7RR87CisomgCl1Kl82C0flrwMJbyFqNCHS5urcjtDEHaLfjsdQDMItp6XFk1OmSyhPu1FsC
OW9EqoQqMXFe3oGfU1uZHxNO7Ybjd22lbn3zcRJgTNHB1RtkYTrKjeq9yHvG/W+GvjOKO3ZzpAKT
t9xNZ3esyRBLKluplqXT9qDMpKDXn2MsCmaiHwL5JtV0+UVkcccqs5h+1AYdOTVH6Wk7IrXgZpXI
2DlBDLFPr1vF7CCZ9vliS9vVHoj6KD6DCbtON4EB9tqQPLcbuc0pGrNfZ1Aqf/EYsi+qpsCRyABu
oKZ+C6Qvf2pJ+fgfY2MqHWzemWPN4N8xcthFyjKDgN805XPBCkTlhOuY/q+3LiApcWzzBXiAm3Q3
6L4HVKa69sToQ5MUc7LfC/Mkz63Gng6kVorX9iGu8dkTrOQ8ouXXyKqLj6yZpUrPlkQriBV92GD/
Z0ZWkgI9+WZwvft9FaNEJLUlAUHsKy7sq69X2QEcag+D4k6puNJqy3xTjnQttowofECbawfevgcm
GpSfYsu97bzH6iuCGw6u3Sli/FMNHzIsXb5NkQREJ+LK3GKaciAEa3PMf3mUktAGm0Lfd+ogb8MZ
cKGEFUMjq+M3njAMRjkwXW0ktYmM1IArYQpcEvQrsJmeaU5iTCEkcIUSBkmad6/chpBM2ssvV4Yd
EB2oB3v1RZJHKuh5kbrGfrG9sUn32xxgNvE5HgJ/x3H0Ajjs9EBD4hbLxofJwAkBMDKLAbO3JUkd
sIu++WMPgut65URkuExuhRmTUIW4RXwUhjjZHgpiRqVVUhn5wRhrHv0gJIlT0dzaF5jI9x5zXwim
8FX8T0detSKaZZO4el6lOGqlHR09ZeiuOZhHHOat6HzKFTrCyGUl42w66g9QJIE/lD4SVsELU8AX
TG0CRJJfWAJppc6jzNb++0tqRbpj6OBvLKFG8hpZ/hizDQW5le/PaaYcLFvDn/HHbKAznxG2ap12
HVj8lBWU71S1LYF2P4BIxNFF30oIID62oLJpFcDGwcdR1HR9VhARL3BOHXYo3mA3PlgUatcrgzp+
kzkqPi8BQ4bw9poBZCqDOl1FUIlbr/32h1B4YC3+DBTTQtaXth89eXL+knqKfG38HBiW07XNw8AH
EXczOjZhqa46ub6cYYIDGRwG09sIa0bBqFq513HzjUHgVsIGdByXvXbM+hpsD8FKdlqKNiDAEhHZ
xUbcYZAXN/PaHXixzHFVxocu0l2+MtsfY8dWHoYfqkk1YSnWBda4kCBkfxFwYXYHrZ7ZgC1a+GGA
QOrtMxkPJG9ba+Jm/N5B16cmC5elilDAYvqm0b2pbiaCrQANurRIuaNwza1vuDMYC47RNuZM4cKT
4ni9BzqUhlSmxGAjgr0NncsGqX4QHUVzHp0Gt7O7yICzrAMJH9AIOyc6Ea3XKcBHQHzGfayLwd46
u6y1N4y9nk34WQ+/g+cVnhN77vH8c1/cmJYoogUr/Dz6+LuhPTG1Ing6AGvVtEIgHj0qIqgxjtn3
0pk2lFdBykkHcICnxJPM54UJzX6MLDXvlHbG/1VVtKYpAyB7SN+KlfcblUh+MNf9TNHdLm7tp6Py
9yuPXrYna0k+Qka7zxx6J/zmX379SFjePCtgDT9V5y6KM5S0DVnqvOD9R6zVqVsp463zAvaK7TS1
Ylcc9touue5Rp3jF+QhTfSXO20Qf6WlEvaz7bnD2iJrwnDRmwbjezup2y8AiLIHL4QkeonVXitH5
uL8/qhgE7tu8ZXQ+o8GrC6Fk1bJyG3vlJ2O7Y2hM+3DWdzj5jnygvT5dWyQZb6QsaxJjk2MksPUa
FILd6hoxFvCW8KgSL57/kHspuC9LEyvt/Mq65790+0yg+7RWy2C095Y02T8PLvNahAM5DnGejHyO
lqlYaNvts2P3F88voGy2mOaaKqRf3/85U9LZ3zc7Ns3gtoTyNTCKyFYP3zwQjEXnOwZ/9wXwEn09
M8VzHmECc0fmN3OIzegBEA4cz8T0Z0Bx+7Pjm5ODCKdAm/B6vsFHwSwn/gqmGfduQvMOBkUQHHAr
2FwCPpalPwU4cxo+/LyS2vvCkEj3V4VTfJHka+fkRip7rzVNprE3hbQ3W1Zdy5LF1itQdgdlSOZL
WKF3WvlnoLYI9vz0cbwOQF84sgc++oXP+yw10wUrJ8f6cTRCXgwFGOFkGVx4F39TfJaB7Uxjy3Qk
Rva5Kmrsq8VbYqikhg+F8Y3GmIvwgZ2PLpVlZ5f1zo3jVK+sfA/OH0MXGOKyH+NhpkVHzkF1evv3
YmH+uB34dRaFSJbXdtKlpxGoiVfdHaQVN/5UiO898xxv0jj9PYWuqmjE4oNvCLvDKOt5vo4CokFu
lsOXshp4LHLDZdrcTaJduyORu3j0yv68WY4h0nP+EHHuqGmo8RITIMnnaj79CxAQaLDjTvH6aH1q
wPHjuk4P2vT0YrSdxkgyu9u4UzRzpTqG576PCchhkEyvDOtFE/FESO6lF6XsID9miz3/U+X21Ery
idGxkZSVvwgaAtsjdvY73EbMZD3bFFNVJaE/YF+Gs8glvaOoal5LUyaAs8rFhDYcTbSNiWHYkc9Q
zdvvwbOhimi+L7LDSyxgWhdFeztn0CRYbpSYNmqTHHkG/0SNK/auy/RFTUKF3U3Vdo4EDCyVy7DG
y6drRAtgdA/YSYz+TdkvxyZlw1mriJDYg7hLtVSC54iIq/IIx+Po7D+lfSlVqegyLlM3VbW/WfLn
SrvqA3S/W+u/MCjCVCN+YH07uo88iHqTUW+Q9d4h8tSC/mwXjWvdQP1WTyfEF1IClrQFJq7IHA+t
pN1UqTKZhGysAHMxLu+uWLpDh3A7i/2eqxHdsMEU9eaBYpDD6rAvSLyYfbnTvHWUejVaTWeHAXOz
EDTtMIlSbPI2mdWy0Y8basFfJoeMyS3jrfmjJVB6amwo/17A3jxUDDlgnUZVDdGnm661+93LjHJM
Kyd9kvwChW+h1uR90qb2nnShu8MKYg5SYBbejxeB/IQiHvIRW+2MSUxSevcB7OSVTKA9IgvbXGc7
GpWh3BVKGB6k9ruW2f4UHTT5CY9o9TqqSJY8FedLnoEhhNfFaaUzE9PAOWJ2tnsIaXuiBp+m4hOv
FKRRVDCkkEzkVO5dkuHl1JD5WmodNHiJaR3xkpVo+b+SZp0OXMulzufELJlCaWK3U6utXWWBRVh7
hdk0xgUIFtXHq4/INjQZNYm7j35Zq3Q2DkHZVBMvOjQIfkvyw7xcsiVJw6lem/ez1B0SARN9gXCW
K3krwS41H0QXsXgzODPheNQOZQOMs8cDVfO1hp4zW4ATlYrBKpeDkGUra8YuDDHnWaHZm/C54hAN
lqN+sYqdklYOuLKAj7IbGP1/ZxrLladKZ5htb5UuqE5+gWO7GLlqZjYweMUWhOOSHcbhR/40jmxA
sWyKPWv6UNUzyrN/ONYpOd+w6i9ewVoQTAEr8h6SB2lUqD5ZJ8nlkNEvNhqbTQjeQTqILO9EVCjD
6ugM28qSb4OHeZodbWGcjan89REbf7W4ut/26iMyRpU+8COGT2FzsO2rJkQ1ynrz4w+c4+0vZLTo
VIuGl0RN1qtHdzm+Vc68DyrNnrZLZiM955SqVfQDuqlRkL7+OW9LXJEDIFjkEqdwYGkXnwEfF7nU
LV3baclXsvb1sXwhgrOdeCl/hMd99Q7/5CL7vftaiE2LA7rN3eL7ID+haNLzZLs+lQdjDXzSg38B
kRgXwwXq9kcMTe66qaE87yZrqoE4ghcSB5R6Sa1x86HXL/tagghosazsUlcFTtw6Yo8qlz31pc98
mHE9aL2KXP34/XJV7D/HAgcaS7pG9LycpVwPkEOb7b6FtG48yAs/GUs1241z1NoUlh7e+IRK0L5+
1ELbzk4zJrQ9pxiDjt3vhZ8s0wzI6vJKX9g9WcoyQykCews6JzJs/tJJou/+pyOoesWgHu6F4M7n
sFXGTBc0beL5bmT8plnFefTVrNxMCi2P753puUZ/xhSuTE9L32VB6Ce8Mxuzlk4p00kf3OAUitC0
8orVWSyZQfq9pV9YVVDR+sIgIUtoYIyJ1Y01BpmE4/DIErnfnUJ1DllYYithN/+flXR1nwiAwv9t
8pgfkq8f0jj3zlCb85Olg+J8KeJAHAS+8K66F8RDpQCcfQASAs7UVLX5QmvEOIDGTNkRWxqihLQA
AVzz605nrrL86UE6xnn53oTARo6TsmjQP4WYFpVT2z2Bgn+iQNjiWy6mouq9lqqlh3qjgq300gWO
dcENoC3gPaA7I1rJk1WPnjq8PLRlX/UwM8H/bSLhxJL3k3qs8HlF1XX4e845hDgVCa7U7l6aaZoj
+y9E+HVIz/kkFeSnAiV0Tyc7ZfPDCo62z56CRmHkeJIWX39q4aHzbx5FjlZ60pwa4+NqUKkOsry5
+dP4FYIGxDY5VLRfmdQ6Z2XGqtTHJLunXiRvhbe8bNRXnzxtYLZRB+U33CpVfj463CEMpr+DhxK+
Bxz5W/H6cp+kWrLLn4fKNhi7JVIqDX1Hnf8hFoh4I/0CdF/GB+nJ7D9qojbyCGREkmW5B9VJchrE
YYPnf5LmqCGHg+oKK+KXKSGQFIbzqSXPH8DcwdbRb38n+raGTmlQnuxGogmraFhB5+2ZYjN3knnq
+AnZ19Ykb3BSiF8BtVvYrDotK4Rwtuy1nflVDBFgDpDpvz3LywFI4/oVo8b7SFCOwd5cEHk5zTRi
89N4p2NyRJmeDze/ZmYk5yqgBIhf+tS06sN4tl+9f6t1JliSbx0cfvBhzzxGujedAFWLb1m0P8Kq
to3Z3BUCN01rak9CCY8x+OhZ/H65tBUJAMvALEJkPnXMJT8yKPvWh8IiFk6kyO2cjNxbarsNfFtc
dQc72yxYFSQiuks+w+Cwt2QqFnCx1FyUs+dQWLmMrtWfN2s0CxOOeQbD4YAaPL8dXuruaGueiiVi
75Hg/ySSRZ6VhL1kCp0wGCnKxDXRZP3778rZqU4wXxaMRznu5Xuef/oolXTQYhRNH4K2EOdMLrBo
N/ABZoAgJM6GyU0PY7H1zUzix6lhYAE4lP+uH+OJ2/sbXI/QVX8COnig8SVJNPwGI6/smCKTTNJQ
eO/3Eq7Y6jzyNw8eVHGFsSwZGISNuXTc3e2/v1vI3j0pbLZOVdif5oBHrhIlev4fWUBexzwYq0gt
+V9S6We93kIQzIvNH+o1Jp3YMtyjTPmC6lF1mn3i9kjxahpyt+WYDyv7TMO/CsCY6FX1yl5WL6mf
4HJiB+hpsIwgMFYDmc2912AaG0lOZ3X206sLuVbqjkOcAN1i1//PKP9isoi0hbdWnYCm9/W24FV6
4WR1ZjGJs3oRAREbkbA4dQ4xiWAd2/C0VvqsRB6lWnhbeVFLnHNJY18XtJHF5qiwI+5ibFmyfRdh
zG3pR+h+haDUSfd5PVIxmpBglIASpx8vFlO5pM54+wyda3/xeNDesjoHMl9a4KjRbDwh/wG5WU7z
WBX7/0zsVnh8IUDJzM7LpKIvELE8wvLw/cVWpDm0XzRX/qhgE/LF2ab+BOKe7Cin8Pmi1YuwmvqR
CiRQJDKPu4gtzmqzmIKDQQawjN+rdiI8MFPyGjj9hjksPlZDr16YaCwS7HDG/WmlphJ5c3VRPjAC
9RzVssp6B2n5GyniXFq6hPZEodK5jtoeYCFWbnezBJllFDMmBQOMegbJl+KAtxKXbi0F4ts/u5NL
BNN8UHTnFjfv6oQHazmGp7DX7S2s89PqLI9+L2gp1ERVUHwRMzbGisTMW3dUsdNfyy4SuWjqmcGZ
9ZBNlUGfMhQO8Bk8qt2EgYvl+FDJxpjE59bXlrEWk+oHc53VJsvePX7/5T/ccHyf4F6bO/iuSRej
TC9s7tBpdNu4a0JTyPAF6oJqtwF/bI0T01a0xkt/Ab4IgD+EpNyyFcqSPV8Pg4wzpSu7a0Gzu0tz
4YgzJlATbc/Jf8N3EYcBGy9tHnIKac/TvhJwNqYUbbM19od611hFTAD0DzRypFk7WYBORycYkvJ2
oR5r9FRa0wsafnls6820CNQ6Sosyrj8DiywgIJ1UAKaaGMP+5WMVK5c4mjWESAJVpW2Qc4lhpDLd
/QhvqeJrG10a9HZzMOXj8vwqGfTnUts4VTsXth6V8yVBgDX1OgbnGtwKkd1gPx3Vd3O7ZO2gFjeT
HsjF4yBCESftLmLroeOr8n9EiOuxXdI9BsRUBoC9m/QwY6M55s7nirNWI4bZgJ0BxIV2B8KtHIYC
pp7ol8eS9Z5RvIbu59nIgKdTksgBxOUdGUpZNdT+JX/gc5kGeLyunrhO9z8lEPQ6S6zOfaA6rAP5
kLRpTErk+XQTJ8l3sjKxzEAWX57LKEkJp/g3ZdkX8guf7Ept/r9NfjbhBoHdfiqLXlzaA0r09Z3z
VFqIa+uv6F8AdNCHjGHaTKFOy8bgUqaJJxrlFne7CxWNw6wdmVnIF9pFUCpl0/KvfkQwdbZJyPCX
afDfQ9MYREOHQDAu6xx25Wj5fkgLn573XqVJHsBLRoJ75phECSDJ956brX9649gbAWzgxVyBM1Ni
CMV5PT9dly0zSob3x1KmO2Y7oBvtxTUjrWfVMEKuZvB3arxdaSP0tjGLbi3BWvJXYH9ygjELO9QI
ppVTrTQULh1ti+UXVbx25i2FrZu0z4zw2vP9cDudmndMzu/wUTlCG7I4nEFbEnaksgCA3Wt5N/98
wZjpHCQVwIfpNINFv0f/51jix7v6XOQJ67/PJ0YMpgOfW/Pvpxx2d2AzzWfqQPF8h4egt4+CvkRE
1TKq3Hn0u8Yu0wW8mj3xniHn2av1ZwBYrYR/bJHDjnfI3Ygi7wqmvpiS0+X5sOJTSJ2MEGdoQsMY
8xYQ+iUaNJjAkUA5hFGwdghv6JIAvYMmHiExbniD2YW2wmshAjLdoAKuOWle0biFZo2osFJxZZQF
12n16K/8G1nBgTHhntWy9hl492zDeK2FQNfhqcBxk1wAKw0XB/DYuHXLVxvybpqVNbVDustgMz9J
i5s0O6KSlRx9XGSd5RvdxobHOkPaG+vqW11qEAIyEEunuhuAA3TO+s6rnuhZWln9mltS7FDVKd3G
eRjQB/DV01E/A9f8d+hBiNyx+1/FTsmNMBZeN/3sgZhgrHuDfklXjDmN9bPaFoSHqyBGpA1FB3vo
QP0Z5yip8LbGx09wy0g6ZY8+2mvBxee6rg4B1apMdqlR1JcUksCdiiz1c/GQzCTsyE3/txmvQRND
iaLGxn0B6orAuXBWT20xpS9oWYZkvmXRnUlFscOdcnSs/k7MzTewx+f1d/qI7iud1mVo+Vw8Ux34
/8aaFRD2k2YdTEERBum7zXXMaMF2Mh6UX7VZtUO9gvQI8hJ1DAB9BJXYasI4S4H4GElU0EECLerb
okHL3jRCIOoLhJk2VEe1q2fSRzIlV2vVhPvs4psZ5/CU+fUJXYPUWyY6XN3aQh7SRsHBQAFuadhv
kN8sLPfHZqKgk20Mid2nOJ3rIIw+a/Gsx9LpNbxQv0EUFzxSsUkP9aIFjNF4QAS/xclK/lgdkiev
obtKp7P44BJDEmeZstbq2yucuLBXf6690qT+9Dvsdzsw/BhK3haZ3WaYg4m35JVwW9Y2W7PAkJtg
kp7eZuC/qpcq+WQKY2/81NHi5zlCkUukSFQiuLQ47uszFlbjc6dkCPyWUQGEvSr1M28RIa1ldNvm
Mkp3kEB3FP6691WhQSGKQE3Ixbkb49SXhprwmf0pOpDq4CajKajyAXrtRsFnnkMbRBE4DIxtQEHl
go3iXy4KYH0LdaEFmROgchmLVFkA+1pX74VdE8VmTmHvMsZZ87MkQVH11Ha79jPwFGLf1LYMKf6P
UN8brg9K9CBGwzXaz5jeS7DX2xRD6CH5RXTygGUPVyaCElwIa79f8ybnmomuqUNHqcZsoIwL9Q7c
Iuj3KOu5JzAIbP8Mf3yFKwPvONcyFzP4d1esWRCvNSGq2xXIjyKbuGAHYR+rPf4CTw0Cn1bSmOXZ
af1tB9RgFXkgOBHCTY3KTUig+lqZJffS9bQuLzXNSAdynATU2voUFOugv58LvUvQw5c5V2Qum0I6
qfCRxGotrFKp4au0Zn8s1oyUk23DzaW5/suKxlHXO9H1TZ91sabR8+wqtQV8LI3LNcoHZRJZuciL
ahyElorCFzRwqk6SSv16z6PWZs1ROAaALnWdXYqXo/XiYQo6OCHi1SdiO/naHzb2iRoYkmZnK1UT
q6CK5XdxX+0jXeoJI7B0alZmWg0jg9Mq2nBhoY8Z8EBuHlTYux0SRBI1ftIBTCEh3wYFo1KIzKaz
ZO4O6ZA09QTDcErrP72X5TSAGe/lXrXoZLilt4NdRF7ryPVPXUdC5Q5PoZ6AEaEzq/+7A01MwJSD
buzjO6Z0t9MycofXqqo/DYkWS5QLKZL4KXNJ4W0wQA3m0rmOiLy5jwW8lCZYkstnxsQsAU2DX8hw
yabe8dbMyecupbQ77t/eef6pFli/k0M4stZE+ydhHB0ynGKA+CPvQbJaZpISx9TlJ+wmoTQPn964
clPN9rJaM+r/zrMcPb/Y4n7iSqqcSir9J+ypH/7uB7W/bEhibMWEP8JpJlJQo8rTAJLv/nJNnCWt
RU7YvVnYcfzkZP48AAqex3NNrevMCLq/GmF4qzaMgb5rB151g361cFuOh6CGE5vZYp173208q8QE
6y+DfovHVnmOtPNcdNql8JlS/bYNWmv6cBt9MeipALSq1gF2C57LqhxjERYjd8ahyOliHoqhNE+H
PfgdAgy/7hNsfDrLzPA5vlK0xzQYVf3ci685DkXhR4QJO50QtQn2X3ZdbE8k6rpp8zHUQ5LSUPCV
/aKPfMWKDWKT3pDuqNUNWegMZIFfWYEz3uU08m5UwjLO5AXTROQNKH3cnX5zBE55XIwcQZeemLR9
Y10HGHAOdJCCR/SBsyidUH0tdIrbHPRRL3clhRjfairq0Cp1LwZKMewXmKqXwCCfSkeqn3oPBbHM
rIvOCrJ8NjSGt0rbOAe3UohbdDEYEDuQ8KL2JlDCpYJXll/vaDRn2XRHxY2ZMFA6D1EdgbBUcIds
NiGNBTzHvKZ+f9ap5QRikqe2PTxPmw/6diTNbAa3zEyF1tuJofikziSep8gX9OafRPZv7iPbqDxh
2wvQes7AxZtlsnRCyMvJWuSkIGp29vPKrUsWoXWL++qBpZq2u8yT83v4F9GLbHIAucm55MBuggDH
H1IrTETOz0YBt6DhaaLx9RIc6h7+1vk61WGdXXDcrViofa0MduX6e+Ze4fO0M9EfFh7gbEnetTfk
vsCDX2HjJDzzfszbD+BhaD4mT2/QdAmXUMweu5NAtRplMUunZncUFzFqflT/yoqXNPbZXE6BRz+D
OQv0YJ0bqiF2Bvs0IQx/GX0WSj/o74QLW4lW4AXu0vl/pw2SkyRNrShXCVBDoLLbtANrx9RBi5M/
CPkDUZp6u++ZcxhfmGiNbw+cJR+9Y+a2QfsL/BzFvwJlJyynnlEWpKimVleNZgC8mIlBKOwt+5aE
1ERXwayNqpT9ztRnBtZnXNVeGaHy9nSEve/fOOU1fMd5v5z3BapacIUJFUdTDixtVmZ1i+5BBkZv
ct4SwPfGfy8PkfVpDx530R9NI3o+RgfjI0WFyS0uknA3CTiWgMp24p0ldw40LxxKhfkkz4c5R8Ez
HGOJDxAH4oIOx+pmTHX4MWqBfq2y84ZTEG6c93+jj28o7JweEVcRNrybo3TmpxNXoMcaIm9eTh28
mvsUKTS3gRZ/eFyTLuu+qrpV1xYq+bdnm7H6lb8a+yOwp6wxb+T4rBxRd6ilWBwXzY4yKiQXcSqW
MToUEZnWdJkH576g98HNVekasl2D1dn/k7K30cggM80LQNFq9TFFsnTXkkzkV1V13OOzt0own7Iw
i7aw9MztFEgmhSmcukggn6uiCsbI5haOVHxTZdA5W6ayBC5sI1fSFnVYKaYi2oVCYrVywRv0JnW+
jAGH3nikN5FF+lVwAksxgNBM8ZT0/BPHalm9/s1rtWzSlEHyG5AhiFz0VP4y3uTv+cfdEDPgrxGA
eeDzNaCUBmKiQG8V3DlumUZ62dAv4ljrjYJozhsYhVPNGBCSSBclNvj8mXV/HopkJLc8jkRxb/27
wsAt0SXeJS54hIEW2/V1Bc2D/Pz9gUNT2XkP/xuHf67GkT8YJO7+4Euq8ukvJ39RKGL8iZkpUF0b
cuxZRxHr64i3nMe92YQuTYxyOGX2S/x+GujBES3AwtRFTH6RH8PwPlDqgUrlY4by8LJ/D5KzMC4S
KuXSlfUbctJ8nkr4Qi6YsfG0t6POm0d+rO80QR9xIRzPE6imxdoDjMBeO+r4SKgkqruyQbCMA8Dm
L7e6uuyGeoSjeiRtWdm+Yg8G5DJ0rN9omJsF0WfDl02/JPA2WiMwQsOb7/aNbn7J37GZ2DNGaHNA
hs6S8zHfJ/TNF2rIhknxtNmxahCGTr2h2o2Qns8PPUuGx0EN7jKeGcAoT1Iqtqqe3FGzQAZ3FH16
EyrpSFYq/F9KkssnzYe5ky5AUxozhcfRnFPh3xW7ensmtAVLaSeaKsNn7JrkRKM0O+l7aA+Byv/R
sLpD1HbnHJDZNEl9ahnlhYIkAJPFHVPacIccdf6tUCo+rvzQ7EPrrnelGxXJq2S/ehjQkfXfmk4O
gITP9Y4Do4t/6YB8ZxrF88/9dddY4oOvXsml53gJvJzXoor1zjR+u+DgX44heVMpw/jzBKizMxSd
1o2fYD15Pb3qJXkvTj4Yy/kDsHUpyikT6v4wzXXku4r+NkZsDFMgTuUJqwqkYSR3re4d8PhKqbgp
cBPWvx2pRxhCs6ak923caesW8gYwcv30ya41GfoO8Fb4QyWk0k42YHJh5PlVBf9YhImGnwFV37Bv
nGNMS3KU/BCcFz6YWfr+nF+G1dTndIXU5+hbGBrZ0fHDECOO2KU2zwsFpzteXdwsYJ6gx74yOfGE
y75KR4Wgf3/QR5t4C96641VDE0kZOb2dgTiXNtDjBHXYlb1b4yWSJjLwkFiWeoJ8Efznj8xX1Clz
DK7P98eqFV3uEbYYG2Pn9QxBOuxEgHCgChObpzzXuVPVTrsJiXphJxzaZo9UQH7FNUBfG8RkpJ/I
Kp2xImDIe7TIHcd/+1zPivffnjv2XPsruGWtSdyShFxbIZHz6AXmMrW0EiB+dl9B9t0+sj2mYHCr
55EWQIlJBe6118qf1BT/nBbdQSbMMyVKNEMCvW+uTelw+eNIhi0OUfOQ4VoTPzu+fwplUmMHMfzt
Tqmr7wNagaX/f6I9Lz36crq+002ArtU9+IfSIP/kU0bLAVjyX3bsA7L0CqvuvMSsKPgFuxzfMVQt
OeFW3mba5HTXqGGy97nxyDCVSXaLa3RZNYC7lfLPm3038Ho9lgpcAvKQeuSp9SLgxMFuBQtHCeNX
2i7PcPkELaJ4y7yw/+/KFlxKdOHtwFi54vucLhQdMno9hgZCZTiZbQFWU+NEMufYuYG2yWT+5una
MVbuLp26ynmshPRsI+eSGbAVSG9527whPX7w/bnlZ8C6DZs45LAldBEfdIAZeXkyRQgbVOU53FqK
zZn70DgVEpiSXscOUi0v1j69IWYmIFVkS9Ei5DAE0yg2f3jR2XtTm5WF9KktlldIt4iR2Ap2xWpi
Ky+LS2ihl+PS1OFQU1qd/Gu+DNY4liDWMKh19N3DSxp1GV+Z+LVyFaumvSf5kcGwCMFrys++aWSg
m2SxEiYC78eLDn4Ac3uWQieNXDG1jD2gaHbxWjnCWDUM26HVQa8oME8aU94rH+I3RojqAPkLzVD8
YKneY4IZPazniaXUD/fV4MPBKdGCpLXOY/f66zgdKHdImZVOglxyuPRBZqxZk/iFmwKsSwUio7cM
uDOi4AYR6BL7/9lJVMPn0O//vBFz0iX0zYp2oMte3WF4aBbOmocRUdZINXVpNxkE+KAIIyJEI2pZ
8zV2UqkDBaOHtXQq/vKvNTAKO1aQ7oHPRBcf7HIO6BQXlmr9RSD9yniULDpYYTLs9BOGqcZFnfOC
Li3y8OFxbr2gmRx+htHWLi9wK4g8BtJqYZSwczJAfqxAgixMQbSS/R3YY3oOkBgN0rBrC24+jUFB
fMq55xZ2VrYim6hbsUXQnKQr/YsmXSzbnSQEZ0Ql3+38xjZPeXA0u2jn0NsSr//mKQU3dLbeJ+7n
LyDQnDhRPtdZPqJgshOF4AslMMHpYIqGw36gHXa2Y8yk0KN8YjEpPzaNHn8OdjeW8br1/OCQJO8h
jvychdfuC8bdNXB7dBbu+i+X6/cAXZq4Bl26sZ2oyOzyGofWDXk+11nyYbtnyU3LCoaeKQCJ1CFR
p+33P+kJ0uGeEg60bD6AQ4vVpdBn7edMScqaZ+KCxmh+bLHzdu65dew5cwr+KumOmoZDc1GFKmA1
Oaxx8L2jcEDIj8APv1uzZzP4krhKs0ma9QOyhQ5nGY4wqDr/VSk05yjsKgpZ//GOmr3mhhmAzLlC
bNM+Y+lrGSVVKsU3ohrLKSTT0VEqfHS30jJNybkk1lK/89p2xdq3Y1G37fmPe+7AAxxHUGEpM3G3
YJEzW0ELWh8/REDEd0eC/9UA4n8P6OFfFKUXOz83mibbmZtKQJby8HdDXsfK5//SoWUz8dTuBEug
qVchAe7d2XAWorZpNERDALCm2wSl2tInhFQIJo94EFN+0X/XVEUYK/zeezJ9C9oAgV4hjMK00m4u
du3hgLPuNQhZuW/l8njVStdugrSP1C9ksv6p0gvTKmuVKQecfcK7AUhDXgn61pGZ8+MavKrLGav9
BAwM7ewc09LIU/AsD1PFovkc6JT6QDilq2IhQzZvnqC+lsgQuUuomF79DWeMEvhkceM4JGE1+Jxp
NTIoLXjZm9DglkThkyT1Y5nthY4ArBzbcxy7YdFhNDd2Iubwmh7zt12H8t5bUbjn3PIbgN8SFE8t
JlwARKzQxZ0Y2sbTm9Gdvl76XxCdUZsyUi+9JV7FDQUnGgSGPzouf2tSlETHVipMXfWWs1SasviO
+wkkXXkF28nfsZHSkW6rnkcQe7yXXxT33wenePaMJmakw1UGoxEDEPoLUq5he1WvDJbojomxdBga
INqJ4Mj9Ku7DUaO5rQcih2ODJlGXaIJ2awPfGuXFvk+7DRex0RaoYAFOXmgYV1+njw28hf7ZaMSO
uNH2oLeX+uQoKIHs3vaKT/6cOgWMaoW75MsgygKY+hpdqwwuTEvmuzA0Q/XTOURh59i7fXCL16WR
QyxMi71G/qsHQC9tIfSkAu2RsZHvuMQg8ZIGjNkUF4I8R6ThdgJEg5P8UqmhO99ZtnNhVEdwy1f+
nmdGwO0F9qp+zsnmWT/z1+N3GYOFAD3tua542hqSxggD0EvUGtP1bom3Wo2DLz2SiZC+hoLJgvtl
v3O0fEdmWWE80kM5uO+qUxixItESXX6uXLaqRAhl6lA6BGxlCLa2QdOTdwBDoqvMHiAUv2TwDpjH
FvVt/Nh5wkBgxt2PQG54ZeVGzfTKphD/EPNVSKY1VJ3hyU97IWa5sEMmMvg3rtiJQxm9JjCZvDJ9
cA/+ir9QK+UFp6pnTF01T3MeiU+fZhP9SlyefHOugNo/cuvG8UCBAxQdQ02TLCbvzpaBoitjJvJA
h6H1AJxoH48DFrws9/ddic/jnHUYUj5NTUc95cvhIEpEtXS/O99M8hBJy+G4GTYvOKpbt+iPVlC+
0e/iW1FCBO0rT+gVl3eomT77dGb/xAinFJiaO+tUGI5talUrYn5fF7ljiVk3rGk/3bMc3nwtMGBE
sl3s1TYFgyuv0SVTxA8Yy0HFvXHr38AyB59PHHLXydy+5wq6Ig/dhzkIchOhFzaIBfUK1581+oB4
LF0qKyH6M9Vf7XQ911o4SXIkVRRAIJfLlB/zwkpI+RJEYOnn3IGKwAYEOAiMQNNJGx+h5t3emxfX
pJzt5hFdxt0h4e6JPlrVcmQNfD+E108JQ/WRve0VWscTymdzAUWSxKJhD24V638tnRMvc0VoBQqf
108cmmPwXjNwdu5Bm/eQ7x0lcSQ/ND66n5Cw55BRIjWGU5qS8mkd1atTnRO4sMW3qqmn8MZ3QFqr
5AJ3iVWbbNagsfHoOXOu5YauhXc1LnwzqwVLCQuHoMCOyR1ZSPwH3S5v5WJDUljMz3edrUkrRhjs
uN4J2JCJO2kiyEeZvKp1AlbpfHV+kPLgiBRGALAgx9fg/Y5s137B5fs1VjjQKR8rD7WLaOb0CzoX
Yngb/YaHW8ueqYhTn5P5tcQCCyHqVGfEhsCUMuF6ubt8ELvyH7PKLSlDbJskb32lt1ad0VCPioh1
ZAgtFhCNScEsMmKdi7dZVdkcugO8SrQREYDS+uMbvEhPgO3LXj3OqmMiP4pqbo9j1k/eeBWYn5hy
YtekhpkwN8B1KOg+4lj4+K/1QAwwkjF6uqyeOPU0dsnI0ZLsEUKf+m1wJOCNvkMCDkL2ZYakKVAS
eDCgdPhP3/xFhDs24Rd6Bk+QmaAB60ZXRsmvb+tPMrN2GsUp+HXoG44J6RoTHyyZSh8FkIGGBAYQ
KVYuxrN2h4Z+YtEWUBBH8SUB5Y8MzRi3C4OzUaAYJUwmR3U9Ty9QQHgTThpl+bndRQx99J/or44M
7pJtjILvbRky3XRG30pBzg2QH+Z+aJye4P6OdGHvrw5mrvhUIkkECQS+BaXftx7PxTo/GvKG7+wJ
uCV9ppTXa2aE7hV9sKBkjHIYbcQgH9LYvRonrc6ljU24+bqk4rTQ+uxmgCtKig4gR4G+jucxX93g
wUpRQc5t5psG6u3W9W1o5taLPhd0G7/Ov6oB8YSPdFDVkJpSH/SidtxDPNX+XbyRUK5k8SMzVDNe
L/1lYjju9CUD5j6pvc9WMTBiu83AwWMrGYFSkTh3cIO9pwB0dmbEr3Oj89DtyF11qPnjWWKTCIuk
WZhFjCD6XMgDgCs7H5i8cWv4JjBrBufx2EHSuEb5mlpMLXSzmI34HcERHJlsWjDhDGisC769/KYX
o8mK/Ad9stW5qfHHw0eU8IEbLyI3KQVul7p46MRhY2Ks/9wdbz45ugS12QbKE3qoUDWLhee6Mv28
7kq4zJpkIU3oLtF1c+urH+2tAeuHMOFu0pjS37QHhtkvuFH4eeTKJTf8uiX8WmZV9GdHrOLEN1Yd
SxUdZO9Ic4nl2NCxxTonVX+6S047uSm4c2vu/IvX9uSdjFY//wAwKhepqK2K366Eru9tvHDPCRZ6
8AhgBodrzW6a5dQZEnlOeovZuakLKAmfJmrWflp/tKp6FK0UneajCWp7p5ZvD0oJ4R29TE/NRZI/
c00fB61kis2xvURhdr+enidvpKujGxdqcNN1ql3wIrr3q2pYfxGi9rs3ryjj2JF7WQnEDX0iqbZM
t9rTLjFGOUA56PxWUWoMdyXjeZs2HeD40bRb3j9uvc8WmQGu4Su4qRuosEQpPPHRE/Kbc2LIc22y
iBIVilCBZJg7hunSnoV9cXQ1GhjGAGlWzcC8vAfap81KNf4+T5n6nd12z9YfCbbml9X73cjswTz5
ffVMRHOpRd0uGspm2fmtyvUSOVUqXtVgBgBbHoau2s+fFDa4PyD+Vhr6blMn1R+wlQbIqCyO2T9E
PREXXwimOJy8lsL0FMF0qlJnGy24mW7uuP9aQgegNTh/UQJZtsJbpi6oN6NqiFv4WkvqCUc6UD7I
Hh4/8BGN5t7Qnpmmo+IDlsiiK7CFXilFsAh74a5Q6AoWny7ZlS5OkZNAPrdXbxIa9hFuZVGKjR+n
s2bUEnv6uAov+z+0iVzMKjz/P4pjtmHmjNyiqCdo0ChRPVMUQyzmQKwGgYENJYDcTXIYoj/nq1MD
riEMUn9hB7ifayFeNKfE79P4AxDQSU2MoGrOjzJKqp3Fe2zSPrjZXqivXsK3RbkhQMpfcPRwKnE2
7uhiKDMTQwz64lzL9G4Qy2whXqLNJIdgaNmceEHCzHMYPoyLbmIwZbuI+v4cc76kZvb7qfF4rpu4
7WbDI7xCglvIokZsx2IS7AtgJfRIwdws+N5R2tP5M412GdEL59RSA1nh/k+9ZJp+Tb/mpcVBXZg7
3aSXihlJcdUSosrKZigD0NK3vV14Zt7oRS5Bhnt7KVSHj8g5GLoOF4qS6+hq5Ij5+/tlQqWPQtM5
MAWBNx0h7Fz8o83y4WbZvn4uge29jw9hVtGkWD18HRNsMPEbyKoEngPODGMy0EnTQ8/SESyo9xSi
mvhW1/Dkz34nN/r5stFg29WMSwOWSNF1wvSYW+WgattPD7ffCP2/2jMmrAumIQ64gur4GhtJ+o/j
kpK3skJMgRasYiG5gfrrqyBvWLRmyMvN4YqElraF909dAwjM6L7DyrJXWveTR5dJTR+aKXN7JNKP
hygchB8qRn1qt8OtXyTJEttMxRZ4gP/Q87uYRsPUie3ntUH+XxhVoPxrv1le7e9i/V5Y8cj0na7p
PsJQqxOHTDwZ/ELfhRL9y8LikZEQvw+eAvfW7miE6Pbnu/c3qoBkqeNzSgGMTIyqopo04U9SILlY
yVzHS0UCddU+q3Rotu0zUKWl33r2RCYIS9WFxquWikb/7EcjbES/NkAbCvoWYHpnSmvXV56iySug
v8aGmGNYl9qtmdrt7J7lypslci/C2cLkgORKT2qG3rbXywgpwTQz0XOZ9eff3NryPXeqp1OTdzGR
MbA7dxCBjbGIN6y7QVsHvMlvAmaAkmx3mMQ14y+HU62/M/dJIeZpoVANLkL1Vd4jJTCiyAElEIG7
K5j5xvJQH/am8fZLjRM3BxmBNmDa+cbxgUdmSbXG063hzLlVF8jkzU7JVypBcfY3sltaDGhnpIde
Cl4OEv7ap7daWUGokOETf3gs7cc510/56SbsBrGJ1AHwBdFQrqtzrB9pApBfXhbZW5G3w9PwFAWg
ukBFEy+nG3rQcgO0tdAGoOJSPUh0paocBZf5iIWHtVi5Pln5PBZiCY71Fmj1tI3UoEQv5J0rYwCf
mpTnD9PLc/1H4UlmHmf7w5JM5eb2ratOeM47F4EbwQJizHalf3pNkhS58CGeAlMCLcNLdD5X/Sz8
ExSlRc4gzbFuBfwM1h1QVg3bb0DkbXsmx6aj9AuaNGR8Iw3Pcggef22V3G1sEn3yUETvJKKvvBpQ
ViAut7/eFOgx5TX/hkK+C54sy0CzO1oseC3L3B8TDGGg1+WIN9GY4hM5eeid26JmtJvF3nN9WtpC
l0NvUnSqhYU3vYRsSnnyzp46DtktQhXJK78e2NwUCYBW4257zRFChgUFJSCkbwrpUsp/bXBwK49v
C3DX+L1cq7S/7m9KlWVUo26eTtdwpIsskTLo5aV5k7nDJaM3VXSwczBQZXicK47gGRPMBIlHMcl0
LFJr3p8oY24sjFqsiuuv49x2X6tQ66JtFZJ9oA3XYsD4VsMy3gQwkhciNgioLvTbCNM/1M/Qn3MN
SueRjhbEG8A2R/sAOq5klUJD4Lfev5VDYc6Yes8zxOVXxVf/Y+1lCXAcd4ux4t0MOu/5Xaag5e5q
gKIb6QmouSXWzELAgC79Fy9v0DV+M6tUwlkpKgdyBlMz3q9aleciE5zttu1FfwR4FlI4d9iTcRx+
PD70SG8zgJ4faKIVouEwuehgBY98la2Xz/qyNG8q988urpY91ixHToVUPoqM7y9IFiE7ZQn8cKVS
GvbsiRQ8sljGwWkMuEyyPdM405qKG+KkpNCO3b8RO1fNxNKf/RVYymi9epDBj/1rEM3E+2KUQea7
ejNkA3Fgd5ZqGyZZaOvzu6FSPMgmgr6MfJU7sLrQaGrS3G1BTWlanVdiaOQqdwxaz5br6vfpUTrl
Yv7j6A4tFBXZMD01dg0/4ndo8OFo6HyKr+05lpcvBwJLIhq0WYAFuRCoRebULGwG9OE0ReueDfx1
j3oXqHP0ptjD48MTwrwwSsWyjPevg2Wx5leSALkiwMd5n3gNYlXbQr6u0IobbdAHhKi8HhzW2+OV
U7sWkmyUJ0ACRRP3cUfJB36058cEe6hE8gzE3IJh4o9gY2zDZ7YsRuMOnNQPZv+Z046tul2kgBwl
7z59+0zOl92aZOP4xADP2YHwiaikCtF06fv+dYf9gsHHLVXnPnoilHeA2Ivg0laY5UBeRsFkbMhK
ccUVgIXZVcY3lHcnPpXq8MVO9J/1iRc7enyL07VunW1JkBUKl0kNxgz/Ojt6jC0iyybJrxtQoG66
DB3o062GSiV2GH2sdH67aHPs0qTfA0zBJlkUHVGkvf5Z0A7k7TpQBlESJEccUYvNHQEE06M45USs
W+UWt2G4J9daoAw3ECO0HvnlWyhO6ucoI+4waF4YPgyfAUmZgjFQsCG+yQhKCHit9/BclJrc+98l
Mhcn5PGdBWeOPBeRGzvYGw+uBYKCXll2WY6nDGukHrkS9yicVV+uIY2gpZEeClm8GclC2vAg7rVQ
KDsudwcKKnCnX91SdYz+SURuu3Tx0YDOatqHPVcMoISm08RVDdk/H7zBjsTRn3y/FMfXo/F4Sasf
YFn4NgWte6NxJVfjVfwYiTg6+AL52BLgcfcCae/DCyeoGYe6yv07vPgw/xGF8WL2YaUlchXdJ7dO
9sSGp4BOF22aNJjlT22gFJLYIu8VC4Q3AC+gRSO8fFIex2xK8XXfYMhuua66lJdP5jTwwwLfPfaH
FRx6MOwl82VjHxvrSg5X6Dp0tAWALFNRBMR50RBnbcXw9pzKNB4TG9LoaB5nC5cv2hG++bWQaGOl
uIkBD5F1gNUX7+m8uOxX4SQgKOWOPy65Pr3VYzn2YsJHnld3rPwW8BnUFFdUO78SQO30Wm/s6S/O
6ZApt8+yi2UA6bOwHEDNKFMy2Pap+/OsKTn4USEITVaBootG8d06mRXuXKGxg6JMggrKNG6/1k7L
tzzVNrWJwnuPypL6yU0k+wEyHTIcLmOP8cFfPjGO6lL4XjsGvagMtzt0bL3JkGjknJz17HKcbDhO
qi3RhcXQVtgh7ikcRuH8/bB0qXLk20MzS3CQ+ZslTeSkqFZcqvDKoTZW3g3AXSrUjdtdmKZn5jm8
VMRKPsRz+4Wzv5/wz7ccCdeHPAqftcfM/P09K5E2SepBD3grKSDLWDrSnd2sGP9iVyA8BgwkSxN8
+xh0ZtYk9XDGYoUDVjICXKMGyx8UFY7SHolO2ChzCVMS/32hdzD9CTgZho5+KhVkEu/Z0B02kX9c
tS4PzD6uVzrrK/Yor0ek1VOywRvyxZTKXxQX/DizOHrj/IXWw6Yna9rPwXZ9veHP0ANhX77dWAei
xKZexjCaTShIxtsEEWzWpCjQGDuC3MRagriF7JgN4pkq4WuEdCVwE/Rvgajz+ptEImGHWFv4XZlT
DDPBvuB3N0dNuvEIgoTUMYLeWqmv26sXmMNvbo3ZmUan59o1qi51xK8xO3/AhC1wRooNEpdH7rh4
rlMXxGDHEKlI6N5ETAdkzUUvxfb/D25O5ndZCw0zxX8Ar50wNniRSAwT82eLw6cBL2cM16R0b72l
g2N45zPnrgj4gL/RJWsvhaqDCnwSRz/3XjC7qWunv9/HCPrpNRhOLHmAOsQzip9y/jXv4IRy/JKc
GvdzByMdOtxBCjC8zkJapjcQpXGs8L7Qwkr+uph3k1Ih5vXlkY8EQw7maiMiVQNdec3lKhBuidcE
KByvECH2/4iKpM++frHmD9+VVXHZGpDcDEpqv5Z2/da8zTg2BDDMtGe4v3T/aoDC5uiie8DmfQL6
mdTNTTWLefQPsim03SpQcP6RdcU/agNHNN9xJD3uMrzvdp+OW2PmiwgL4VP2jwWMIaDMhusmPQbe
GSqpWPzVnvhFWtprT+Tbx6URRsiJXyp4V4Zf3vm9WgOm0MHKu34tELnbgDU/qmIlexzFi1dzpZZQ
LtSlFAvaVJvHYU58rEAMnrELlIROPQba/CeTgsxtfkSmfj5x2SgduZpbfkcr4zY1Nvskmkaj8DVU
3FgZLgykmudzVy+rQ5WCQ0BcKa7WthzNwJLS8ZBvEma8HTFy7ofMCZaiycFqvzQRrSO2iGOlnI/r
I+6TVk6mtDl67F+SGgfKMViXhkXW9cljRxTOmrVdkGz2zwV3L8dW5a0mBQapnBko9X80YFwjBhrF
ymJnGC29vDEhFaDhl4gtsQksm0pvCcnnMDZMhHfc+3JPsGZSkMX57vJZgoJS4yxDYR2dSGQs4VXQ
xaAr81Sy7Nrot3jvOc0W1OjyVX+yurrYQ1FhaiJr5dbj50/fy+N8l9CEpZtMdBo6Z73E2chPzuUy
WRTyPN9MzJvhIzotrevxx+c+gBsT9zLowUIRD7MpeCEbPP/+S4IhaNIcLeqT93W9dQhe7ga7hoLf
zGuPBz4D84b2U2nMiQNHcFCzaVBM07Od5oc5Aak0hDuPLquNSAypWwxh2vdAr+U2oGO2JqanJeGt
CI60dqHScW7riV4me+2C46IVk+dJRJY2f4vUMl7rdnXyIKhaNfwHTW5mAQKgSF7uZW02WvOithAh
f5QwMeOSI2axe/HQcP0SwzeJEjPeGDgcSLbKIlMLB1Wf8AQxFTBR5ROh4IVTPKhBki5b0YGFmauT
YI5LfwZb6weUyJFZjFn5oCcAKdohhEJ+2eCVLnw1uhpkBCrMHU4skqzdOyypeCSCi2BCJZ3ETma9
POGbUI79OVgaaQiKJfRXWVcgrKYpkLjEIoVgyw73/nTcBl/VDFhryMvCn5Zt4uOw8aEKhVvbMp93
D3rn3EuihDERewCImeXPRUJdoF/ZOFuPrpNbjYRPaSgPjGOatkk7vQyaMy5yFHfbDrFD6qmhHUmF
Gk+W7yfyb6lO5XVymJ0KFyn7Kf5Cl0ZD2C9en6zdecOWNDyvzxrQHvsB0ZeuxHNADI6P0iuKTRDb
nbBXZ4SrQHlz+UMqoyIVdtKA+K5zNfugW7L6W1AkN1AvnkOcMC1cYF9cEioyHm/ucVrN+jgeylwO
awV+nP92Y+pnYorbjUIZ07KiKjweGlxJ3M52MZqhWsLzicbp8yNAuT/8McVJ0aQM5Miy1S+CNYAg
ufENU8Crx+wSdoomFsjMIjppOjWcQDvMcSBuYBZ8Ukos9gggGK5f11AwEdyhTv8zlpUN50N4ia/+
T6uhEjOvYl1raB91smhbTh5GQ5aX4HzAdRRoM9wJT6i5vHz2TTt+9A4fZRV6w7HBoUeHJg0ozT7L
CHPsrY0O+q0pUAeD2eBbgy4bigBYIwVS2ftXAqHHhIN/Klu07usDnDjlUy/zGgx9IACYLuXFKdRy
DTf6iZo7w5PhbBrwECRGr1/rWg8m8ubVo7zfjFIj9E0iQLs4jV/MNyLzATUo3eS5jTaHF+QkwOoc
yRPJAeenh4OiFyDl2j35B4RMl9S8J0rx7343wOWWDUZXanw+Jpq3L7BePdL24xuEj0oyoh9b90FX
mT3UT0LqXpJfo6dSTmtT3XWWvEvHfIuE/VDmI5LKoJtREcNUisa58gsPXXdZ+36RA9KdDSmnvR2w
emk16moBpHNHOtjpwj3f17FFnrq9IaLmpADZJBOIjCyZlL1KxXmzmJRgNEK5J1RZ4g+7plWaeMfT
P0x0aE/5IUiUpKPZqWY0Vzf6umbuslUxwg8NzO/4Mb5WQO6t9tJC4c9XKmvTHVBusMjF2xDDz8PL
Ld6HgLtt0iceTQGwQUVEJM7YvdbAV9eR+b1CJCaB2ObEbTbhpK7fr2/S6oZpU2llIhlLU8Kk4Kjn
LRnbWo8mcybd1jvFaAIUQW0mxOhhED0Jl2OiXEV97libMdNULj1CF/wwmCuOf+U/7EQOAGE23Uf+
S7BLIMdO6C6nM+5GmP8WMnkfpE+orb/MUEGxNr3sQ8qeIdSGwp8PJy56mY0jcrcGECuKhy8dp5Ht
LheV1uXShk/5cwWVkeZ9KXkJb/STxl42LthnkMCFC3SmQNBCthPiFnmePdmK1OWJnRfKV/smcXPe
WUAqEp8W7XMnA99McdGbyojZudcCk5i9EOF+jnJNY2bFuIq3wS9Y2Z8PVl4mqOn5Uu8mA2Dczbhr
6Hs7DFgyblqDXp5kuudjFa5Me6XsQQ2BgL2x8Wt4S0wOdmYMnqU+AIoY8gEgwNvG8frwb5ygbBIL
sgGvan0mcu2YUhjobo6beuanFe+lQVI/EJxhtUmlYes4gQ7J80qUkcNIMzHDRld3oOTeCRQpIzEu
WlWY4vHBkSQnxs6cDqFB3g5S+U6fSsBzl+86Ah78aVoViXlbGPDcFPmsjbSd1RH70jFfXRFJTfRp
o3/3TfRSf5MXL/d//YL6oPZ75w9e+lH+4OeBguC/XpoTrgK0BH4/s2xLjX3fhe1nvY5m5DIF7+pj
JMqWiTZyQkTx6LH4ErjmnWQIxLgIsBV0zV/FrBqE47yBIKFv75yOZMvUgCbRV/PG0Fyh9kwfG6w6
rlZbNVmCXl6qAkYQBaAvLyG8ABX3VYdLBcPR5609AG/lCsRc23ZiUI96wUmBKpLqTkEnUjIck2j+
YBKlZpa3Wm0or0gwn2neRnZzc+S1JCTVhYsZfW/jjw5/zb+6PtN2iATnWle5oRVksr9+osK4pB/u
mCX+mMhLNGBSctQVYrH+cC5abiU7S1zx+ENL+Sr9y6DdlPGNKvixFWn/UfB3oGviWcUyWDgE3YtF
hb4syXNwKGOC2YtascrLH3jUCyJCv1ghE+CfkWdVrTyBdjhK8p6RZGEemDeo/5vtLYBYiRi0QpAu
0Aj2LmvuslcIQE4ovO6xnWdJuN9BrEUVFjpwDzS7WvAAD8o59LeGUepPbFGI6zayA4pxifcw1Dbf
l5APVCavE1isdZNzhnAgIEjy29Uv4kuUzsmSBOQ+HD3cVZwVSM9R3hMn6Yc6SzqpQidkD+u+TnHk
ARCjNgMOyce5lgIWrwgEPdbqQdn1ro5doUiBBj2eKo7kB00LldOPAgjZPevEUo7rzEKWqijzePh8
cvh7MLJqTs7NVK9WZ9xXX8Q4x6q/niCTElEICf/uopX4lybVSCHADqAcAsJSo15h35zzI5qn4abN
CtJ5mgc+OirziaoDEFGVdj5GU73oeJJ2brycKeRovSyEsk5U4980yngi4GcxE27VlK3S1MByKyTL
1uMozhtIhA0bUBJi+x0xhpepGwmylsxh6fbKq3oxoMg21JSsf0z6WxNHA/cspRdJtg1meZXloeD2
tyb9HU7OFZ7o/N5cD5g2JBOJgARbn46HKEvd1S9/FtHUhLi+C4kdhGz9a54HcBYi/75WvqHPBlfu
mv+HL8BBQRQg2M8weIpVeiRWntQ6apiieSVx1yiZQDyyD7Tdukkgyy4pjaYMTgv+GRX7D0nwpL4I
Y7BqTEbikVr0TzhJ74ivtAvwNgMbF7OPODB5Uk+o2E/5d+4TYDmqhJFhEYrCnrxUtDP9h7R1yP2y
8EWWF28WS1ld2nt0KkmEDmLO5vRi9rGSJHKWbiQdhTFaEUP31U5HKAP66rezWFOJjahDzEwNM22u
mjYgZaiqL0VChEHxK9naBwLPB3JUsqy5q4JZjN2lxZC64ELpY2GX9UcDQ1QKEwSzn4jpJT/dLbor
D/4wgIMxVzNDx9p5HfMbJYeB6iZdCuM8Da+gcjnjlFK7pyiqBvNV2ul+67iesoJ62J2cOn87NNIp
VSJWvsajOV42ksXZcSEkwwdaffk0O/QFRYJUhHptWBSSgOxf/IOq0qhrlsGVRHG+vQ/NyhiT3kfo
bkUsDhTbWuXqNRTrIkgJeJJd5PMXBtNjiz0RHX39AuGypTO9jTDx1rK5qc19rfgv30pTWtGK0Slp
yUcuWQALIkDIAf5/Kkh0AzDQs9r1SGkOC+nYf3lFjx7pgaFAVdrrSBqhDd2iBozfUu1KuryLWXIo
WIXdaYiN26WCCflLVhrU6jyIBrbcE/qloE0O3muXCYoUMIvLC8X23lI8G9IpoX34X7MRsEFHVQY5
Qz4dXZTGgBncIPhWPHmOi4k2ZiqKKuNT94h7hKv/0fi5hkS3zPUlb9cpq5SvXAliL/IFAKiZR3fV
fa1H29Kg5JQmiONczpK0GeOH5up//01DTXiaBtfoMeey411EhGUqHYFegFxmJTCydl2ScONVFlYD
32l42JbqSeZfgnufZrBYe7xsD68Zuhk96E9d29wYGNm9Ns5QjMHNFO2LwP4xYvQQNLystMgemTNZ
npGEnmxiLwTW2Q6p7nTxA9Ht44vBUSfYnViMG1ggMCjDRX0UzrgV7+Y9R7MN3w69boBvEc2/8eGd
m5n+JcHsR9aZm4u7++CWca8VZ34c+5xFGEm0AdwS+RddQqJ/bBZr9CUxbaSXTxnbguuzWHlwBGdz
N+QOv9fSrrIuSMK7Cye9mfcBI2ARy2fON7Ijg1/19Q310ij7ToCfzYm5FswKbakvJ6TTOoI+oA+U
Xv3OwSPHdwyCV2If8c867VFGr2dwcFVLbTnHFbJ9QOnytsJ8WjpGLWtihefHyl+03Uq3J3bdkuKf
xHNVS5PM3NRFhPGEqJq0BuJXpjtU5kztbYhvMCmz544HwHVCPkZDQX7y/AVi08Uu/1JOnQTn4mC1
qdO31fQDXWpTru6E6NG5YCnd3bwNHG1uppcRzkhurpuaFMww31RJMus7Rs/lBU0iawvSv06RYs7D
8FWC1ee4+cfiObdh6I9ZTbx8IE7B6HWy5scrQjrN0ZTjGhz97hpoKGBkVz47wIGS1w+BlV1FoxBR
DXX1pAHQrUIz8lYi2IbwazMnB/b1lHneTOc5yC3UFIT7WSGq3v6w0ybOaUDfR/o3WQuF2POpYWqK
AUgajmDxEFxQuDFunASrVZL8gF/7FEgQM58A4PoAu95buUkzt4e+qDZVMxEbCigS2rihYe+vxbvz
46nPVAUhWYOESX5Id8jVlc+FLSCyuD/KaaDSUj7vQMJktkKSaX3IrQ7DdihdnKlI87WBInpzlt/r
YNVT51jJCp/9uqWl9jl8wPWqv90ra6bpEOBZFlgztPtuNsq8SmL3xsZzLGLvhoMWoH/Yhg4u8qUD
rDjxnLuiF2bMkoGRT+JEhn4PGYvMnzKqYn7yNeDSUfotogBxDt0gC6s7cdM4e02W/XivNctOwSlA
4Y/d+Fq1uLEbflOi8PyyGMbyj3gaGDZkNHKHeA0oTkOK0/XuQxguDkbNWVc1cDYAF78VvGBT8Sb/
A1WB8x3CrJRgc0BBlmNsHfOxXYK22kOuOYI0Kora0YV+Li1v8+svCDsksWp18HrkPi3Azbbzaa26
FLngm/OdgRAZAxKoz8q9xFFO8Awt1nyuew7ApxPj+gYeuI63kusQdNQwkXsbOHdvcUTS83CJI5Rx
WQfD2PxdE7SNaGz3ou8mzH3Wm+GK0LL9P3Ar8h9cYf22cf/YxMfUFm+J1bPyMiO0wCtNyj4/Klws
bu/2QvRqfcWwwKZXeQusZvJfJJS67wqfv++bf6ysvsh317RefVMf4SuCwUcqFrSVGjk0uVTZi0aO
uiY8h61lHZtxM1JjcM2gOYs7g+Z4wfpGzJTXaJatYPofSlOP02w8UC/2Jh/Cw3J8mqrFP+c0D09Q
0x7qmKUbFDts1w5sX2lcFYjFPwMVWVhDMpOEcNa5pUnqiv4p+n/19BDKxzcnp2VLxmst48elmeax
CpblDmVH0RS0fP/pcnwgkaVXjtgKMG6FiL8oid5dmLVcuzItEikWMjioDREanUALs6H0z+L6ZVut
n3Co9qoZ/xvlS52IXk3qHtr1ViUVoeDxdiV7SV+PILz/LvKM/TylPrl82hsDIcxggTf/rDhUoRJ0
L2xBg9jGKiNJDLYg8DejjxdQnayPgUUE/wfOy9luNKfyYbdZSNolS6FnxMGWh9bpn6UL0Dsk/UXE
sGWMlBBHNcFIwJVoRUTCjiRLja9EidVNWE+UyZi5hNknSY52W1sLQfJJCkId/zvF0vhlItHGZzz4
E/wXegb1rfUDywRq9P6zySblHZbZP4ZtETtY7ekT7GOk93flxXbjeyspPMX/ZnYwjqKQces/+xYl
F9yDUfpp+SYYfnesV5qSSeaBxNgzsxq70WFzPTLkjfDq0Z2euSpGtKOFvqbN/fnoqmSZqWHidcah
J5+0d1s+8pg/aYLjLeEu9RkiJr9rFm7zyQ7TtNXWyCaPjnPOY0UbVPzJdWY8WJAwbWgUb5+WOc2O
XMfbWQvHvouxFTVgqYprX1FVvRCK4OqYt0cujLO/e4bKckyAXLBhkNWo16QhmCAUZsSp/IVNOoQl
Rw/RfwnxevxhiM3KMTPhTKnFv0yj5l76zYyXia1K3lPM3DG9OzLMSdggcY90l9r2d6AZ3I31sQQH
eOZiEYCqhMejVrzK0h6M/eb+SjJfjH2cSHwYkEqOsvsQQlfNGs+l6uZ4EmyRTcck7y9EX40XCe5O
2rlEboW7R9P3VnraQsd+bq9ZO5hQQ7+W0fJCA/riZWZaCmieZUcJkneqhyDfsfPCRk3tcGJZBn3R
7cTizZGmKTP1gVW6zV/HLt5C56Dcp0SeSD5hyJXAFLdzFRiC24MfQbJT52r3LRQ+0LC8eWWBCVQQ
MOiMsQnFEkqbVm9wicfUvghJkXwWModJpouytQue6g9FUL9lG+xQBLbdfZKMgFx6pIlhb7V30fAR
/qsrkdmwWHnxdeNVyp3lJZ3f6pK2cZq9xRl/TBETBNakdxdjPpAh+rgk3tmNtk01SEiOjZAHo7Bo
ChMfxJPTOD1Lt1YQ1Vv2tPGRQJF2qQhnbX+vCDSeQUmy2iTMyRfKCgZOehp8VZTyP01yx7L68595
HhElyHpnsCMuY1fw4M2koZ7CrbmhQyI92FgG9goz2gvitv10HNayF4s5mAs0zPC+GVmWcY11i8zj
wRPrJCOD7c+kUxjJFKvwpAo7SxaXNXVVnSIUhoTW3Np12lhXR5fbZdm4E5eWmCm+Cbwdwjp0WtLr
nxn50tECBwu0i+WmfKXiiQwhm993PQ+s0Tr2qwTKiv9gjM6ptCqKQtTt6uMAhP6A5HzdcX2gx3vf
BlIfhL2KCtj9c/0vnPfa6ZPhNcvqce0JG8jKkGQRg8OXlljAKTs8MEG5YmK3Ck+n8jdtv2KtgtGv
5uvMKO9a4dbRfGXtS2+7x/saZYntlXPj+oVVQdTKWlvEjtTraO1GNd+bloIh7ip/g1kd+5k/o8vz
HKz/lt6NJmQOrho5qQ+KILOTyMGRG6FP77K3H377Twz1bKLiLCer4Os4FCoORBT7IKhH1o9V6x57
GpswXO/ytuDRIW4jENn2Ql5zVQc/mPut8nj5dMNoDvRBXeEbPGJ/VdLUPJcauVt9WwjvJA0Z2Abw
+LOXmiZZXWZhZ7fY3s5gCDrpS0hCYKcBIUvidCmSdiRdxinYho2o3ITVXMNaPrZMTPd692nEJJc0
Nb5hfRKoynWoG9rrA7i9rBB/W2a2bRRQI1rTArp1fu5y9O6CF+8/ENzG6YAOTWy9PlLRRL0ehRU6
4Z7LLGJM+EZtM9KVvoic5DqGa8hbSkEWOs+dASWeKGpWTOipexVpC/fTqrnpDBHhqypj4RvyIAi7
D/+ednWqGjDu7mS6QBHW31gaz42ecOT2pCTdd5+pxJL4n0Z+MBhUSO9WsA8r1/LgU4pNPCDWtW5n
2tICmmyS8krj0InPJwEU8iFgOKSjP0OYHRVPJD7gOvwJcuCRD71h//p5koGvTceVtrhWvZbFtNsG
sppEk7lhSqWchdfmMqF+SxZ1LDdJIuoRU7GDkeGPr8u7WX9TDoEh1e7IoluDrG9v/zgE7hvC72j/
cMjrTIN7bDJ1nR9lO64/ABIhq21ZgDL3L+Ww/8sqeagzFZm3DHkJzmkpj21AZ2cEchS5Gy6zp1xQ
J++S0xRPNGUAKQA8SPMxHMbYnAb2fIUA7mEWI6MdXhenslAn6MGcwq2oOvoRb9knTdubS2vtkqEj
Hbg1oShOutdv+XxEurp3TPEcN9HIeb1DcnjPAUmNMwi07r7hPdqgQBpugsz/2Vys4VCI8XUyYio8
HoVHArYRRC5CeebM0LdTPL9P18zvD+zf+fIDa4Rh5f54FNzaIcYx+FvzaHzxlYrmV3WJtS6OQaVN
K+9XPUzATlpo0KC96bMyx2Cc3qek7Kf50qgP0oczV3dEDoepy9w8Votigat5dE1IpLFAfMxAPj37
cgwpHJLRYUA8QFXEmkGbeSw+JRy/V27Z4QgcS82c/lv+W42CHAvR0ATX+fXapn0g++junHHuDzXJ
U9Ai65FjJP5X9r9vxu/KvVd2GRZFzz3JwJE/eJ6Z7f6w3cybbncM4GvK6VoR9JbAMVJgZFKBQNfr
X2if6OEiS1/JDqTK5nzu32WkhIaceVOSN0vP+wlEifxQRdnk54+34ZF/qMjfIOb0ERBODplfWC/E
p6djD9eURP5W6zez70DZjz5LuXFI/qZBMdsHcT/6w4kgEsLzvrGzrqQJpPhJgJ0z9X/eYF5FyCvo
83zb0PXMf9Ut5fXbOoVO2S28aess35tQ0FpeA2NpAZWLhSU/dazIYgzrTkJYzjBQ5Xi3lI81J/To
KAazJabaM1QV5ZBiALBTalCs3hZgEnrl9PoAUSyZJpuUAbnpgHXkf6qPXB5oT24kPWT0sPS2WAgy
H6spgBtSxOgYaugfC49/B5RCG9ekFKoFL7D5M6xFuR4FxGQNpHyBoMMPquusvHwW++5nUslcnoss
zlBEqmGwilrAtVMEwLSlKcAY43Pz33C1HNnje9vP4str8UekYdMzL4jId1fXOjNZhvehs+/Jr/q1
CTT4pUIt1MlJU/mkdXxZGOA3UlgXXGvOXZzZzrITWPeh71MuGw6zkZavkA6WAAWyC+KXGWRZoEZa
KDTo2H9iU1yYZB+Vi+Zt5maBr1KtLsHTabUVHGJqQQsh0/iHDQuYQ0Tp6hvpEH4vpa4tIJzgVlRl
ttdraWu63v4rE7W9Dise0yPOhLMA9DBfxBGq/g+p16QU7yKrw/5FPLeaDOc3z6fVQGBavnsGGbNo
2X+ZIpezU2Q9DcqCqzpdYyhRYG+r7qQMRphpgh/opFCkfMqd8XK5GfiKgtOD+P3xpVw4CbUtEDcN
5QV6Anmpz4e+xvLec4gLpINa9ryPb/3yx9tsoLiinxtNMZwz2FnEdqlwDFeaAGBNiMcDDzJJpgNl
m8jmUQ8yqKQ2P4QK1S5W0hbpd5tktv8fXSBdsXvcSd/q6qb5kY/isYpBSQt8aI46FESw2tBEfbGE
+OnQ0qX+I3bagZi8gSxDMSiZElY6twRnb48yN2Xh9DlCscmi/mbP1Pw/dQfCpMXJ1bBO+HTNKqhP
j1LTkZtlckthUjmm+pTz5sQ29BR7hiEGUyL5P0aZwnX0fQC0v0FnbtFO5vgTSyXa51DTRZZ5YCTl
ZdqmOwVaRPdfxleVyOTcZph+SbqrMKwYwCi3mPoMyfeUos5VS0xzd1Jixu+VkdcW/agt4YU/MNt7
iWyHPy4xg9G6hnqQtUJNWgdju4XUZv6YVGrUGJdNyoP3pxo8wheVc3fzvwE1fBbu6Hq2Of9wDmyO
XaYRbC5j/3Le6jpajgDUERQfAJvVrXsOr9XKhpIQZiSmAm49NkUzw+jFsxqPIN3PAtsQuMNKAEB8
Mx5Kz16EdWeUIspVh8Lano5tGPmthxFj34II+f8XIBZI6T6cOBj3JyWRHnZNaHz+/gHWKTly/7N9
ol3pJVDQcxOKHiKdGSsFnK+fCX/Wer8MfCL4coRBmUjL8Xh8VMnsea5bZmB3k9Hj7SglPQfKDfJw
rdMFLITMecnRi+Pyg02X5wM4tjdysSBhylwUgi/clwxaIvWU2xR2rFv3BqdsrdPO/pXJY/hbuzxS
FA85StEHyLh12fIjmR4ukBqxipOD5xw8Aqwzevla6Bnmr7+7Q8PRyPDq68xDiGCRAKrUKGNY8J5f
t3bcz6CM3PcHpgDVPjR6+1EiuFyrKqqZN45m30K/vkQ1no7QdFgQ0Qy10j5JcunMfPnZpezCGF7I
RUgDJ7Y0KpuxFCEeCJuTfciqFKSkvwYL1wP9d12WBLGcBHWMRWquNVkOzMMvMlVA4ZVjH8RbovsW
ywJTGr9fiu1tA5Bl9IZITUH5jV9AdjEB7G9OtuM8UtEJgSk3NSCtIWx23AZZ1quimU7RC05vDicS
aG5p2EWHOG3gpE+MHKmN5IBXu0HIwqLpwOo+xErBxhA/+WilxzA8Px3TaEpFn2G2QUWzGYQZ605c
AMl28txeYvBO1UIwJ29OxUle5BarMUd+54zoRWDgu6+OOKwvqM9yaRaTosAAX/aNmfx4uyihFUOk
D0x3A2woQW6KXQKQVJyxF0K8EWQGAiP2oPfuOW00U3WpivhmJhqep936PqWx4sdE53glOFlrblzf
2sSg2SBALS8pFnCab8ZMge72bsQVrxXClP6XIHRBcHByUFLjPo95XUFN5hDklohViv9cjCHjkDaZ
gtzPsXQNzYD7JVDsUv7grU1wmb9lZ8MdVb5R6vYFPcU6+c6YPHY5CmCCcnJTkY1RLgvRPCssLAgp
7PXFXV7IHXPmwc0a1gvrdbyQMIJX8kAJ4w+OFnZcrUAJ+d/wnBRPBByUKINmbtIC5EJtRpd+xOmc
RdtKLzti0mPirixjiXJhvjwXstf6K6Bmr7czn+MO0qFmvjvBA5Y20vPbA3dXibb+FQu8ueN4MrDl
r05ys0vBPwYLYi/fxnPnNWhOiiEcY+o8wS1ps1g3Ba1uLBiBv1tvk8twQlhi67yTpUBf+MeVAKNE
MDOK14gjtK71NEF7PfMoy8Br9yfhznkloHJu3ABD5Z1WN5lD+NyKQrnhM9upBkiQ2Vb5wxx7wwvv
iGzTCu6eGtNxNnh+4/gkTrXmavQZ6Xi/acqcwcd0rbMnIdmV8qETCWsS6ppNm9ie/9O/ZKJ6IFZr
FKIRKGlzNspji6d1og7nk4YQd2U5URkmFrMNWEBKydwHoxzwP13YStDNrROd7GxpxJ0JwXRJLDW3
D/6O2s1A/XmXLfKNJg912/fKiV2fG/W2SIhCOVd2gMFSFmRspr5RjktkAKr3/Snp4Ra5iiMd8vAG
wylMdOeoObQUdNgofnPRrQZANUMbDXRyhFNAPmkNHjGSs2BQi1YpbQrGnZkVjqsv41NSjC5OmV2H
G9xpYYIv9N28JMYx2K2VLrITQALSq6hhuB1d63dBxPQgepUXExLJT1Af+QmBYbfVQSvdpgL5phhM
ha+Uvhz461Cz5DmJDbxvbR7wlNRN8l6ZzmbEA4AcbAz7aXK7T1gtBwByVv5yWn5OZFlhS5ywt34J
YTIxuxaZwqBN/E4T4qjFe9T2Al4hBlYKDzIun5XrBPnebjwDhj4MKe+cz/JxVtnrTLtVWcaHsElA
hzXEH58JoZ4FmNB6fTVkSd1avFWiawoKcNRTktXcuIag11zYKOxN6N5mIxT08sdJDuwUmR9B16BL
rh4Wmm7gJnL6/PuXTlynwPWkcT418LwmfI6Jgg0Cytyngm2pPNCwZ0XUtf+vOUErN/Vb0qT8Kydy
sruYG91wHx3PISbonDxvHGIEuESutjrGKFJXnTFjJ0F8tSpeU4e60848trarsL3BDQ0xGoYT43PI
oLb4JFj1hjsk+7Z8SKOOd1lvCiSP8IuvtaYE3cajlJmS+1zbMjwgStdOfu0tSFHDJTTcpoplaF+k
HYP2t91AXiMD87Ar2+dUYFK52645kU0SekgBXRqx00yzvGzyx4Yn+mIObFcYv6+yO8K5xObx6aOh
0UPPgUAHGDzqYNJoKBrbBfc78k3pd5MfUgUuy7s9YvnVwNjG6ANjynL7LhRQX8vEnUcZUguAC593
V7ICxSF8o+aeiNhBCz8SFRC1t5Ia6973QzzE2Psf0V5Nxive7dY9+hqYM46cBT1AwBOfLj8pXwhM
yPKDDu619MZDrkBKJhoyzQlsG37mtUdC9/Qir05knmKnDQDbjp+sK4A8k4JCSDyxSccnFHDFe6zt
Xs4PM4v67BtKKuoqbJT46GlEGMps+M8s9157hYLJyndc0i976mlULgXKgJ/gY97gpC0qdBOyXelH
gY+strBlGYgTnD/+YSV5qLUezlsaeBvRxlzDH3I2azy2zqgUkrbqCZwKiE+T1KLjASocR0ZAFfE+
Htr1gHlpjVKMX24zDgddLnuqPguTgWf11kh2r3rIT5eJjEsWMOdHIHCuWQiTQfD3HMfZykJ1Msyq
TNXkkYExMyOpyFM1OcFMdECNcCkpvKHXCseuD26T5iQGWYxqM5gL7onkeSyUZDZkjq1k5bI2pTk5
iebXGrTDLVhWxCGQoRD5a/yo27U0j9QiCJFx8RAn2Qex9YczRh6Pq8wmfZ/c+Upn6Q+CxYM4B1ei
jIa7Kbi+LHu13uklfiedLULLdPJiTLcND/mg5cJVBBK1M+eVa9KGoctxv8RjE97QQmB6BF/Emiqu
caWSUVG8X28jpVh1RhEqBfwYCCUxgaSyQ0bOUAaWlWunuhG0WNjhZr1s5lHlRPn24bOcr/dz3TI/
zIzX649L5t1NxV/SuC0OMPcBx6BIhOxSXzoIUxTF8mBbjgN+V3egs1u6WtK8E8L1UeMOwgp4obtY
Kd2vOaR9ItBDqphct/sUrhXNHePmUn5nAaJ6rwXwJVYDYnTVFFpAKWyhTLza43RnBhDhUc867NHc
E7PdJ98uIcv/KafLrPFwrug61lTEwI2vVQpOGozGWIcl1G7asNC3hiYXHAW2vGN7Zq2MjdpZww1g
Sa7vXRiX/FKeZV++DLu54hJtSXDiHhWaSSGp5GrRarPmAWgEoR/qCvkL0e52TdJIGI4T5EVb2EgM
7GufZ4Q+aIYuNyRYtNtiJfWjhWlo4STvN97L0/PxSkcVrNVWBrTUhSR57CyvgoRolhDeFsnjWKrh
mNVSRaKDrQrcBLg4FZK9ziWEBbIJgTOHA+kpRgRoUVGFCdFeiQVz203X2wLof/pztz8bi2SbNxFY
In5DMkNd6dF1t2k974xGWJKnY0TWTLrGO3yhSlgOeN0/DWscqVI/GyHcMHtLkxe3K5jNbIBfK9ED
ew08mwqyCmjSArQDJ4YXDdcfTW848yRvOKQQSvl1OuCXCdj8NbjKVEJdMrH60Xkm3qcw/2Ds1WYB
FK2MbGEOgBwgpfda+Uhh76XzWnTGmOx881RCvXuJ6WqNCGQjohdg5z8gzn64+nHqmnV2wi6jOSIj
/u1L3y3jHacZO9km6BDDeZVCreCtEoxk7Vdqt04djueSUJVd5ftZVjEB6Fryy1ho9ky7CfDNYdSy
ZUsTC1hNmR8V9TUxgtQpSmEVrlBx5CSpcbouO085aMt4igTKzHZiRCO41cMllv9HjQPdbcseUUgX
XG6Pik4oL2/UjdpfFMg/THd4d6RvZ63OLp9PdEo7ie83AFlZV9wu6p70HMa5yHTIT3WJNUN9P6fv
uBirr5gAjPPsywLDrNGyGChSWE4WA2102wVlIWkbh2691r+J0VWFYdZG69VDA97cUsWaXR7SoTZo
9pIwTvZuH7vajyYdI7pO71AyNcasgJIjYXjmJviSYmWzp92uNwZKa26APkRfnyupF0qF4/BHPqCx
dnMcnKSzzuG1ECGA0muJ/cPhiUGUFn2BkxL3LiKTbTjXE8FbpUl0SHzJdrs24EiQJHeep8fAQe4s
DGTMfmm3iIYBW2LQJjQQHll1BGtXOvkxfDq+rDHYQe2Ky05Noaw6UEhOnvomNGlIgTV8RBNQv9oT
4kwQvwatbAYI5jSx7k6JPythwAP9tYYWwMrsuC/eRHOGcGl+6ZLwAefOQlb+/0bmTXmvlzi7UJt5
M68CV75sTUrdgRUuwfnRZmrg0UtWaMpf6Y/WGoIrDbDREYg4D8vupfGJZLPGiRY577QbSyJr5pEL
qYox1b4rbs6arBTZJDyPZvARQf2IwKxNIspaIWhPZuzJticPiQkfh/l0xD7OTEWZCfpXcK1a66Sd
BDkc4+ftEaS/vtAqUdsR4RP6U45rEZWgS9KHxtqHR0hRE6Q4M+kMarEEVFQrV4x2K2M339p6UfED
NVasHcTTihkAgjBgUexGe6UTDXfisP9uM94QcdPXXerBFdq1sR6kcidW70llN4Aj8bSj5EM20Ug0
A7Reeh3XrLqpUTA/aL46pKuUvMI9A2mcUmACPtz5RztrKZVRDsYrO95xcwkt/N4u8t5AeRngmywg
ox1FXqciRAh8i2EbGGp9n6cUhQvZCCA2DsjpGPHLxokuWL7wabmjPctC8egSz2Bjvli8NHy9o0Zi
dE969YvzXceZo3HsgG7Hjcefa2MUAcy6kk3Rryp1M2D7NwK+7sN/e5orxsFPohamI2W0q80AMbi/
ukmZvixMxuuJXqp0wnHR5W/+/DS2L8LXpherrByoxiPvr1iBgy7m9DBWriNxnGWH0+LllPBHOGdi
dTXT1ji1b4QmqIadJzJYN56i9lxWY02GkiEV9SHsOZcn1BgtR9E8gCrZfcFqxlN2g6bPlHrl1s8h
YJAANnHuHe87rxOe68GPsfyvLCyFm3yiwA9ocF4GRGv1DdaPrgU/sw3PkwJiqXkO4Rncl2uW1n8a
HU8WgS4IT4AZiCmGzoxJL1H/BFBX6R/e9g1GPhU+HJjAwBThTKKhIQuTP27vCgC3Kxf98SU2PKED
nYId8U2IuNkiVSRn8dyMiMHaD9WCFaNEOXxwQKHPG6Ca1ykSZOplrYotaoiKw60Fzp2joRBkx/sy
JgKMQtPWbC6cME6Qml0OXvRD//EJGNDeAZ7wVNUm2/aLF8v6PmPif0Ao/sPtQcbe2lewZfXHJrOO
X8IamC4ejtiB/9NljiAvpZx44OwTo1dXM8csa9czh5tIWbuoKrJD1PSdOXGB4mVROQeketNp9nnp
9KpvIGauj4YDRc0AswgEk6TfAgjsENfQiWEhzds/I3RWdEaxs9jBfQrS1Gr5QqFtGv/b8jsccEO3
keowCk7WebjdcTrv7rTYBsDXq/J0Ku0Ief8/Emkmdt50Iaiv9grK5wfiy135Nd0ydMTRsQ4S3txl
n3g/psnt0bL6Jc2OyhLHVJbwBPLsqlcGI9QOlhmL6/flg7lFu5Cx84A6mSYIJ9NBarkEL2jvLPGf
ObvkUyh0cC0fxQkM+oxwg1BSPkyEd9aDqx0gu7E4tozj6YFydXRSpZqAbSxg+3GraqCUcmGGyXpG
PzOXmZfwlIlYXr0Wuwr/CAO3yd/EFhsPBvhX72L6TJ0Lld2lYA1PjxuI2gpIqmYQf6O/x4Qsxv03
l3qh2vpDJHSDU8FwoudYUDoXedPxBcWZkrV2K4awof/b7wgUEw/LymgGXMoAD099ESQMd4AZ917B
NVnU5riWT6ADRAZ9tRpOWx77hHwXUoiyTsKKYrCfAZToSpBqyA4BZ4bmRlx2Xn7mS/owQ9tE68Ax
uHNtcOeEApBbmjQb7zuY2eu+y51KLT6WsZrccHTcIcQTGpvA2b/Jr8AJYiXgKq3xd5NKoNqUQtqg
e3TSRDJFKaQou0u8exF2cwu9/GtO0aiPSDFCya8o2TtOI0USVBKM6mRBewQ60xCOTG0gmLCaNL7u
dcTHR9c3ZY8hqwNW8T/ik73Jo9u5kUdRaYmh1S+u0tX2OI2Myn/ttbYeaZoEiTAFisLwp7UPMYqm
k8jXKEB/MHhzSEahcoM28xyiIN+Pgq4kcj0/QwsynJocZBpBFzKGYUXUvRh3+kZSQOTgXY0pHFhw
n+Q8HV+5YyZ65tIjgUH9F9ZyjeJ4W5O62KOGDUQEggq5gc2YR+7/cctd32YWvmM25L1XWi9lsd4d
kW02lGcswhgnPr6onRp661O4KtcVk7UxsvhkYdLJnzKWwX0P3BqhWYz18wt7Esr21+mehRPWTo6g
43tVGvTWEvyZVjaJhEAHwnNtDb2IwgjTqdm+Z8cLX+j4//cbzdlnU4GbUgqi6C10mN6UIDSKILqs
JaFou2MIgg5gVRHRcIWXTMWGuSMBwaAbjZZDubcZ4uznsWyRWtiFWcUa3dNGUiTaVHTApzP6Kuow
Y4bNaftoZUmlyvz/AyaJarhlCyhdSml9Dest/I6I3EKCs1iCIi8+1NLTr8wxLxgzECySYEreVuRX
t24GfWgG9PB7LeAVpxOUb9GOilnbMDdI93cmxbEMSE+ztv8zoF9K9aYsKknHe5+puryYJmEGmdXA
dt/AIk1QyhVEvkNpy3gpuZXhhxyKbo4n+MjOFAYT9yo0jah7vpV7hr4cwzLLsgWJNHwWR10e5PWs
QF2tV/9doimX5FneiuEyw8SilTNwwpuhf/ndpHd6b7i+38W32GxvO3LnAzcCsxVEKn9jyO/W9h2I
VJYIJ6dCBOir2nbaYjyaLWALdqVPyJXUpFMfIhFuKjlNiQ9Ct25uWVNDfEL+sU48c2C8DDMIFBbk
dlo57fJP5370wg5EZW0pptmHde6kF5OOyeCdkb2UkCOgCGorHAnq0leZfUkGfHcwl2REhoE/6gyD
fXO+9Jm3789Ks9MfQdWMmykldc/sIoAKYGsnYMgDe3EIqEmZQ2ACq97B7xjLxWN6HX1/nlPIrP5p
xw47nv837x6Zdyoe5EAeGTB10EsUtxooiikhSmosZdjD7p8Urufz8QlhizREeGIGbNhiU0Sl43Nv
gSdDOOwtdGni4CT/FJtlCEUAEFxS4EUqLHqdRAfiK6nwn9vuH80sSQcMt13V6KdqXzCTmXAoYH60
Q8m4uF9Z2AfLQyaLK2ePLWh2xT+5sNVAs/k4Uz1wnlRBM7RhT9MgAwIAR2n29EXWEB44koA0wH82
vyAmdsqP/p5TZMd9HLEVQRXAL+P3HazxxsxYMsSN7caHW9BVFw3ZO0V/xhn1usmivGSE3nxHqbez
h9WL7WzCxqZp/8TypS/4zLCFhaXPSuESg+kpUG720ZNIL2Q6lQyZCqOv9HhtiUFKjQjAbArv1Huk
q0U8aQqs5CaEadKTLVarV5LuppwwrKVQFO5GmJabYOtuSs6+uc2mP4Qn6yH0xq+zPL5GNcNrElH6
vMOuHRxkgd3nEx0bep8I8W6mDEwVtYJNBssnt+3qH7hzIm5i1xB088oi41qWoH5nIRFm19OkA0dk
S8mIlyHplsWM55pBHwPDOfC7WVxK1IIXyyI9AMeM++vogJ+l90ZE12zIfLZsiWT6rrSPDvpRoEXj
p+Yo/lQ+9G0O/Zf2swS2Kr27CpcPpHig2E1+iuB83yxo0JnILexAdoG2Ktk1MA1+PN1ZRCfSJKOT
rt24/sa+Xo4GyKluDG6b8RHfoe5pYfk2Ciok5EYcreSxe3zTFE1g3x5CnC1cGL0cUsEk/QOv6ABd
7DAlBQ073f2Bu5WCv3+aUJjEPtfVgWoteSkFSebZ4gJscEVhtXlFDsMZBCbznBlQCM1cuCnOuee7
uTqqm/Ayt9+ftVy2t2wcl26MOJofo5qwiV279liVjrbllN8Os8BbrGS3S2DgL9V7OTPIpJf1dR6b
J3csBVoA6n1868VgkScyQfva+MbBmB/RDm2IwLVbYn9fq0NiZq90jfgNcoY3suVaqXQv20HBguIB
Kq0wV/MDHQskgVWtTylZvaGbNw0PXLf2lIHM13oEaMIVO7uIP4l+MmHPb1dps8lgimcJXZntsChj
VpxRPEQ6u7ns6nVVgIleZCsa/4gMbFNA2Mx6Iu/RVGMfUoGS+5l30pTaqLFizxw+Q5TX+1CDVE2o
WtGswk+9/YAUocBKIUd2Wxo0FQcmvBSPdnIeswVAKvpgvnWq9rZRq1XyePF3aTNY4BykeYsRGoN/
Im/5/RVCjb+1XxG8PqMaQzS62TErdxAD6YuktXHzc4TeVax/88BgGogN1PXIGOUD3J9q7bYQRcOa
ylMiyy3ZM30BQMngyyD0BBRnzsQtlWllbACdmKpAyEKEgn1ZvEKF+2tlMPELW2+12H55Lu4XWA8R
vMEbei6Ei3KF7tr8LFI8gUrFghlI81iGUJw2XZeIuPXPZW5gl95GNDug6i5v5z025Pyh3WOj2MGx
ssHAjDhgK1gsac2bSDiJwB7yH9BW1Js/m0SkjYycGjP4Qw06+bwFQL6M9JQg4Lbs3pTX06055OpM
Aom7KfvuNdqxzef22POfGl+XHnP5umBjbEMp84cflWxhpSRzmHitGTDS1EYXQCm7p/ES8vFtjCHc
eXG8g0Py+IrD9pFXGcMhutqdWbnQmGePuNuETbt1at2meMftngaLAwtzzGDBDBxKHMivhfstvoET
+F8DM8VL5rYiGhlVLrbmm6pQy2uuVJ8QKPpc9xUJNH+6k+1+anxMgXnDG3NeHHBwWYmsvKhZsMRy
GCs5l5SN66OwM80pBUdUv7F4wYZlLVesXXLVYu6gps+pYyp3O2t8smfb/JEbrVzHw+UdhPlBv7ML
ERngwaQN8aurGANGMrphfFJnWnj7gKc1k2g7LR5c1GBTEfY8YiPLPMd/SmzBlI2QGYFr8RVWFzzP
Z0Nsao78mlVRO/O/mz+eZDAw+qlMRsboOl3EquuLqWz2vNruplSFa30dZ5Of69xAlszxZClBaWTw
s+OaSI9RWnXtqSnvWRWDAv8kQVTaH0c/TacdFk2rcyKE4pX50wh1gZAwgn7L8ohk3DihEsrwUVAu
erNABlNAjRzJ027Ywnhr89cAdl6sVWdpJaiUnWTf2YxdiK2QDLieARW6LhhXSW5mDe3Wq4PO8PXN
m6LBLqalJqPEBwqPvEEVfG0xal5psfXAlLP2hWfZujkC5/uyeFpQDXXNv6TB9i3XqkKR6SvtCWHW
VCjag0bIkkBLJJuS9XK/Wf2fxfriPpSgr+sBc4xuSPBG1npQ8rYzpZDYgq2P5jQJmDZmakQNyLfe
+P5dOWI6nsi7X8NNMYA7ACcZqXUdl1BIBNVc+gfK4w4seJOTXlRl6yTZlHdBhxBX5VyNCoGYeuY1
hd3/C8VxK2nvOLJdp1O4z6qp+a9jKqloKqSlK36ubTPS/OLnsNkoip/93m/7z/0DLt8g0a/U/sfF
FYUuq50TJWkHudwa+C/oP04++gU3AVtdJZ2w30qtfsT2F/FFMe7O4K9bfNDv7t+Y26ig1io67e8f
H7uIgBot8fpe6WnAJb6+QV2VV27vasHqPiK3BfpfzW2DZPxnsdHyRA4qIOxFkReQizkfZ6/Yelbs
5iE7iozrnjvQB+3eAdquJegjBJDWHXegccEF8UX7tk8jAQSCINUrpZdS5Fs+/fYHBACe2NRec9ZY
lHTxUBZAHA1ibJB5jXQLEFhmNqU75CPV6ikAXgvE+aO28DdCvmZ+3l0uEcYYffV+qRv8PDka2XW8
XRKaqlzIEiDy/YFOkVYo2kXKjTH40XuJlhLSDyoHsFIAb/fVTotp+wFn0M62w3BpaGJdKtrKUzrZ
itW5boN1vewVffwRb969K+5huhC3CH13m4t513waWavdcbuHMAl1K8rRArOt4Q5BuPBpK2nF1Gb8
bhjh4peDoNHvMjsByA2+ZJDJz0BHJ2eNzInxmYhKr0uFwbGKaOZ3LRvhNqCrh/fWwe68GgCvlYJE
HHevKlmSF3C+8i8wxoqD8DTymHTdS0PUHSon5XcPyZDsxx6cgG9NZogwHqNIoOexns66ns1uivCl
KPj+lexJOK/WNf7sdauc//HPflgxpsk5yc6ew2t8ijA6Af+Csq0Ez8z3nqmyjSzcXcSOacz0LWqh
U/61h6GkIsIVrWtQ1Fx80cvKHau9+T1qQfsaVJyxiqhsj0Q3WWNlXmPWPEVYUWlFkxOwTg+9eWNw
QUhAD2h+M+P8Kw14Ye5NFoaC/UYs/SydZ0DAFCv6l+TEZXTFL0cTT4zFtdTudSY7HStzfndd2Zh/
Cy9FMldkdtHzoapV7oADn8+s/zneddx9/OVYEZEa9fOSwE21bVtQ//AXVWa1269Q8lxvi7gsIg7I
PvjbFciDKPiyn9S+PR05kKtgCbDw4qxIJlDwrCPCFS5K4KiKJpfFvAvlV8WTjYMtNmRyIJJJoAy4
WgzFikUMHIhhhxsSJYhN8f/pqo+Qe5HfgHnSWReppfrgVgKq1d63W809bQ7FR+uZ+YYMT0bOBCgM
APSoYOeJ4xvTszboKGSpiLCUBUVfcHqnwj7qAwhVG7NSzGacYkbhuQVa0rWijg+e7MakqW9hZaOF
Z0zRGSoGdeWSijGPIoi2hXHkSPoP6GySOwPX4t/N3SNuh9vqOFj0/eylWOBbozJwc71WxlmXkO6U
cg0RMpVOUpcrbx3DZBgwjN0Ptsds6GmCWydAAsCJMviV0WIzCXeeN210eU01jPe3NJhML/16JQrY
p1BfEq50IVTNDDuK7JGv5z1ptJ3hrZmbgyJTbSJoG7mO4VUOxujxOemw0H3Ikm0m4WqTcWcr709d
RwhY3wa+tO0uQD2gQgMCBuoLXy1Drlt5XQhl78Tr6a2GVy5igvIYlF/MKQspH8mjdCgyxRGTUhKD
KOy3N2UTSVcqatWn3G7twL1kwZCYkvZaM/sclBykFJqqIWfQD96/cWjsn4JkRu6Du2P43nLT3KWK
XkwUaCTf8VvIvzAj7WiTMlMREE8SCVLBpCvZJvMMEC3Fj+8LRoPiL4RbmleFK2kpXzwYT0VLwOhE
mBTivkAbYkfoDsFX79fMaG/6ttHs9hmwoUDJsqy6NGZ6n16fGRrB362NiWSc08eYi6/YLqLJ+42K
sm3ehA4z5RcFPDhOgdZ+qcFZVTlqDNBdj8QwmJtA4ogJJPL5krMdyiTjpMAGJyKNs9FLc103jPex
bXj0VxYlUfg0N8/jelRcOBeFUDnwXNqMmqMJUti+1jYYcBoKvOrgoyNck47hDSTzJP/vJpZKD7p0
7jYDsDOZbafqkW0mOXH0YH7MbohjQACfnQrqGPeb/rBOwphy05LKHToPFLoGOQTER7HxUnwlGpuV
VGx+t8+IImuScwroB6QUma6dlMM9l+5f31j6apvyjyWZUjoWSCAHPI0BPniNDqfiOyL6+iSRokIW
1NHINvg41oMf2R23dflJegdGM6t3HdL0ki7P3RXqQOzoaJ6dB7Es4VX1U4cpfdIA9IjppESFF5U9
FNPpIHkGC1N+QS7/CbLWMZ6o/xXOexfo/wpSS567y37S6T0hwy00r5iIcEfNN7jjDIf7vQ6BQw1N
KBRlUOd59c+JJ/MAv4Bbjzq+/AJvQwtilNkJf03jq8SSNF6OuNURwZRvQFvu3k+7kEIjNw7Qe/9N
uAQsYrXUlp1dJT+vanCTA9AeWZmZwwH8s7Jg7Y2nAdQ83qpFQocbFhSE6Er44oxjAPX2BWoY+vIL
euixuckoa6hIWFSxcqZIYdmVnt+/AhLTlZtg9tJ3lkfLKzDY8m6dlujyD4Li80sfpJqQGxEaIykL
GqP7iltmKTrOtcH0UahcBpTHJFri/kc05p7Eu4r16FDlRfp3TOj1v1yc4TsL+ydY28sR8pLjhi2y
H4TsK0j3WEnya3xBPZLqCKxqD1UQV3nzYmPkuIcnfXkH72uwIPAmGw8g67+WV6Bt32yLTS/tb0Wa
qwsJcskNv6YIMXPxLr8NWUF3kU7kBztQbHNZ2Kb1KLzmfzkPSau7zMNH6OL01E8o/oIH26CNJkLf
3EX/3WjfV4aB2j0eRApcSaXbaJKz9KNIVKaE/32mOiRAYnuREJpi/JUgGzixxcfaGQS6pa2Hzdog
ZBf+PmIa8fvaQ1NSliWT4gX0YwVtNJW3qzFDeK+ufRh9x47xaKIrY9EEroh0ofqOQXeGVENcASyJ
tx/xrFPOuDELMKJmn4zLWwRrB60u24w7SSLbJgL//D6yWwjv2IWeRNQ/rneRKGShS5MIBsba//XS
0fXF07gPaiioQ5Gg9fb54lOfkAw5ovU2si/7lCOynXgRYg2ykJ/KNc/HvPbHgJnkUoDWnD8q/MKs
OUMp9a+xCzCl1AyxevReCtflCtSPbvL+eTxViCcaNG85EkLN3CZFYXKCciN2CzC3C/68rNGTs91C
24woBTzqrUF5bDb6nq/8hWDq/SfS7YU6q0sPUJK9nW4JQg7Lxa4D5pjbJ9Ib+eikhg4ujTKLo9GQ
ZLsf5xmbt8Te5WKvuqpgl8vdyNtl3JzLSS0i7WdlVa4NlOnAvMK8FaowHqlURGWqc80eamZChcHi
20nonURXWALYCC9b92B/+RMdU56mQf0yC+4rPU0IxsetalxykCEi6X+Mj5KInbch+e9r/bcwpXz9
N+LbXMrRJrOK41EzO5Yg6WKJquHwblrECqA9Fb/8ygyomAvOwL0SPf/W3wpZ6hAPaVp9otX0ttzO
aCKRqtHLYF2wwIeFv9f7CazsaUvDAYiXfFPK3+xmgp5uQahdIs61H7e9/x0rJc7V3AmQ6g2+e1Pn
kQer1BYYnxTfyd1G3rRzqOfh/y+W2EBL97j+Jtm5uoTfAheW5PCmHmfkareDKX8JWOMwjuCEcC0c
GgNTU/ZuD6O5CC9KefqsCjxyS9AcMH313Y4zVRCf/XqHGYMuhmoldJtcpd+iEMlE8cuVL2W3eTD6
hDXSggYt7tBABYwyl1C7E+S2ymVM87Er1mRQOjnCubrX7nupQvRFMIermFy4MMP247suZtJ2XVfu
c/cVMSYxYNvknMHoE8mqGR1oi/nE2Il416A8yzyLIIYIe5uTKhFUVBO7mkoEv1zuZPhaRw4oMxO/
oG7Js5WtWwwS2x99HsttXH15JNtQ+pg3WFV86QCPylOYKsZyHY9y9bKcqZ3V++ymw2lJUIRVbcj0
TlaDkTftV7tA8HecbrypmalbYHFP+SZogIQHCDg8InkjYt3gubtvv9NSJtD+4WjqA+5skujow3Ae
Z1NoztagVqqM4ciYPLm7qz/wfsFITUDjAY+vWvwN+ymrJVTOTw7MOv+A7pkHasxFm/Lbl5bB40gr
t/zrCQAgdlB3HhKfgtadDo7pCjPrqdo0agb4Nt8POgViIbCRWY0fWF26b2phSzJ2Q86TJ86eo8pi
Wo4MPuMy9tO0pBjG5skyyJVvhEsy4r4Mh3MiwlcDE956YjTnODHWSlRuIS5IdRKXM0WCyLuaNi/w
sCslAfLb495cUFl8n52etxwLDvNHRLXKz7xQlHHhrJvV5f9GH3SqrjEMuPjPnDqchxoSrMHQDXZM
eoddqt4a/qs49FcRw3u2+Hl3DyzAQyMSrUL0EhMIaH4V50B8NBjKZvMWN/aP2rZKTm8r7KKXoI2q
I0O4A3+8B/G08CM3aI5r9hMrjeDGindmxJqoSSlRUR5yVMJdy42XwFhSk/882zTKvEij1yOput6v
Bayw8jseLf7im4lI8dolDb65Q+Jc6kOvpJIvzRZwp/M9WdOQMM9K363PiU9ia8SZiJWGyuu7uioz
Pf3wMsTFxMHCq/+TYvwhh9q+iiikcr0CR2CtbmkzDZYgc4n5bPb9+tlQbSDZzf3Qv1UOfhw4xhNh
mwfwpN6yPGR6+GHElLolH0GAhRm1c7FJJfPja2KBC+GOhv8eMgiq3vo9uIGy3LnG/gNEO/kzNGdD
2D6FZzNCmFekoCYXgBQy0vle2aZ5wh8wjXOWjGGlLOoNQyZCGI/OkavS397cE37aj71HxtuurxpS
Asn3yA2AW0kC6Va+pjz2AUPUZJj7v/UL6FTs6NWG7dgylIzLQ9ApMI+u1KRWMxtCC3OU8qEzAtds
DElQg10PG3GdhBFGfXKcWkrXj9BNGJGX1IHhubJnN6hpR8030b7Y68CgMLdXS2uH35gIX9knr7gn
SoxtUg4aqi1g9O6H/92NiqME888U09fvirJJvXVi2gonnkl2pEXealCPf1HYlqNdgNbj4OJelu8I
hMJfIbEZrJ0oXkn3b7YvoHITpjEFOcJhjSj4ts6j4ZiHZdWP3gpLUm7upB+/QkttcjMSKqF2TO54
zSbARgo84NDtj2z9d+X1DTZS7DaJViqL3V34jOllhbX44i5T8N4TYeggwM5l+A3Obp+RCEYGM7CH
caU4+DEasM/PrNhoKKGlOQGztlCkQTJtk16G91CQht8/BKpIcYyvvQvxREMaXSL7/TXhIHihO+3F
J7WsGVSp/GpB7z6DviP3WsFpnEVWX+sz2XI7N8tOxaM2GV9PSA1py+NAynQO4T0SZOCgMXN1dhbp
x2wkRJI9TxpRuclXccgg+a4KOG6GuMEUO0H2XXjyGGZeHDON/cjMf9AtFE90KJ7WFy6RnBixJyN5
ZEb6KAK/LK6uM/HLBjHeu4ey+u5BlY/+dJK7IhD8W4exzAFDMlvGtn2j7qVpRgNfpeghYDLKteiD
mgi48okqmZr/XIKfjcuLU3wCuYwuGLzl+YlQXOZdf8db/guUDANa5Rud4kCkdWVxhp+T8CnEXjGV
G3jKN/NVjVS3ACaTNJLJRVsq8Ji0Ua1rWQFPCy2RXlyGdfk1RXLu1GnSftHc5D3kSdeS0Mx9ZX7/
ngMH9+hrpNdpBDOCLuJOTr6XewSh4JYIBeRwD3yxn3KG/AXAMNZaFWvMM59RYnTPCHEyY5nTof0p
tE+KH8W1EJ67b+RWZUoyWJAv5+xyX4XqJBcTAdzaTnDQoK3BX92omjdB04u+oFSRgBjJJGsnqvnq
NqgL134tSb5K5/NYTBT6AMZBLnvjDUQMWpAgDkXlc13TJc2FlbdxC8RqVRdASf3dHIA6kxxHw8cP
Io3F3K4O486zFWaLTEsEIl9L+Wh8SaGJPUGkKjfFcZ/kN9L3DaEQyDetzEKzQAkzPWm9tG+AP0mn
B9FrBy9MCgza/hnZq3ZBI1MG8DaSYegVdZpNHoNf7AJ0FKVoZHOowD5NzBY2Pv1Cd2mcdnoeaYCg
hcTkswVR+AxX3YbwnQzQDcxTmovWgFhsqj+cDrPRlJibhea5LSl7g92CBAuGkp7Dracm01CO85yw
C60Oj0zMoD9/dKsbN8nb73TwBseokZ/E4msfrQ4JHCADV6xqmjxkIRHFfURU6x+7+nEvGERK8b8w
5E6iwdqjjZLVPuxPzdxjEWjmBah74O/8POqVUHv2USK2v+sJe6nuTln5TyIDjMp2ezKFANtzVBrd
q5cnR8TbdEyuuE61dYKovAaxL+ryEyGtD+lXwjWykQf+hkESaYFR4xvsF8F7o8ptwUaBF0rYS8Su
FwxhwLAiyjNb4SP/HRE6dHgi010GIRI2rZxQPSf9RQVvPPOfZuMEB1GIGy5AIl0NUqKfppRnl9i3
Oij9EqFw617mAv6O92b96cpco/g8ExotUtVeVBZimmloyzg8CSDT2K+TbHPNgotXiqmHml83PW1m
ROA3mBNAGIMXKUtg9lbjzqJpoZY5mKzmadEGSyWV34wfngbsJWDj4GqLgB6R092DBKfPBo0TblB2
5xoZ7OMbC/pFeKGkYBz5H/7OZ5LjXU2CkKKT432+md0GTbDhtwyQHXMnm3WPGZORPQlXigCxujiI
Aa6FNqqW3QSby2PpILAplbGGHVCvUr3Prnm1N4xNETYhQs+4S4WW6+us8+gKQ7DLjz0+idmMxy/y
U+PpbPv/LjD3USm+kxA9/SueVl6g57sMhVrqXA5sXuQqAQlNATQLPTFx5xirrvieb7s4Rk3Y7WYv
X6BrIgwlgjZtcNhrfy13Sim6It+0ufnSsMX7taWYp95cqGK4ppwms8b+vcSbCQLckjivhTbRVSG3
jz4hy+MkFNX8PAjbRp5aIIg6W+wgIRSrI8cEoZctWbSSYAbNhebYEE1xJZpfAW2/oZfOKVxP+LyY
V9RZ2KkCL1xCWA29pYNj5Xh4QAOgwh8uMBlMqQCe7PA8SJ/L3bNGSTo2nMNP2Hv4zTqW49GujqmZ
a23r0E4eq59uTMLFdMQL4YBlGsgScmv7tsbHsxpNlVpm/Q6JA27kwp7aJyy7necx38O6ZjwGGQvM
ijUYFneHm4aVAu+x82xpR3m8BAb+L/PLdlS2bdX7+lhhAFcnx5c9WJahuNg8AQE9vjQMgDyqnoLS
6zv3lA1fSn8AnUJAnc0F3nFIgowXNVaS/dsWLEtdQoKHS+7wtKPGdzcWI846mwbRd12bo/BL/GMJ
25nLMDm0I5ajIuYlHlEK6xo4Yglb8hyV4hioF35jIU650co0MgwofFwSF9KPs9lfHzLF6IOiwEAc
yAhoVXf6k5YIie6G9NG5JQwlOW6k3/hJiM8YfmLxmh2AHlhIBURIV8VbVZMYLNjmmU+LW/vFWMIZ
1I1t/OiDJ0AjpDOWkRgqKNkIp9UPuJqbDYDJBxYqKV449JSl5f6qzg/mLqIhlAaZJtxwuvVBggm1
XGj4DZZqR936wuvqMzf4lb9tYKBI3UEVIPpqkYDtASb3C9zK/1P+Q0Q2ZXn6eZOpiiTnBLBQAFTr
rpxHolLFC2WkI9GIztpP0Vx539eWDQE15kyjC/g3k79FfHX4t9GHeJzDiYT1fo/nisgSzWXyqmV2
FJb9EAiawZn16N0TwfA8dgDs8ycZvY/Lnx3fKz5u63t/bl1Grwk58+iB46AbfXCF+HeuRykG7VCf
YgSqI/EPNhZ8QzXPUpXfXLH/BfqTBWSeMKj+5cKCNP7zYmUS9NaxpaSrTUixCTUVb2inbqJ/u29W
gQ0nsRnKVQkkfQaSTLJpWuHQXPTzcNSicbWBdwcPcX1M+/vgTjMFq8TnrTUo9bng1dm/ULFTOciy
TTfSiQYTp8I+2BPM4LwRK1qhqjkXPczWpehKDYXhcvmT+eA02iRSaC8FiwrV7aB5unGqzmZNOkle
30oIiR6ETMXrzXaIouTGAMhmdcxP6O6koE/unU1syv2NyjkKnOFrS016YogCrKLjlwY4brKMOI09
JJXpu5JtrH8DF2ZxitwPqWov25MWtWX3j8Y82KFW6NzVBk6No1MlEdTpKspQAUJPUZ1GFcHS837y
BdBK3KPJ552/9tmVscgXqZOAzPOgeJjT3iXta99WcOPPC974T6GFs9tryIrTa7H9LAwoJ54cQPG1
7XHwD/LhLN0Be8ZSEz0EVcrVhUEMWKVr23lG33Svtl0NIVadwm4Bp39lN1oGWJZyg20woxm2unok
A5V22Ploc9BNVmLjf187AHzfrI++WQJ6lt96y8yuGOiP3aQbmxPSenQfmwu9MYepgv08CZ9/d9qm
iYWdPAic3KN+jUq7EUofRcWQk8d0MkLsqYs2Xioo6CglZbRYWODld6w05YOqypt7QQ3Guym1L9Xq
2Vu6/Uc4sEx/SraYk8VtRS5dhar71GVZ+YGpSOZJzbvaKt+36IsJOKIxjVx27bPYcttHhY0oLaAH
tVGHnLmKHFw1IB0KBiEgrPd5xN9UuAmpOFZEbuAKg3i6akP43kBakhNeaD6wZjimUcviMFQmVy1/
kdxXy98qM+ck7jqZXYF2MwiDl64FE+jmcYG9wyLDjUuPXOOeBOFmm/jwx6g74L+05RIOsTByVURX
+bjQ/Dq6O8Yz7b8vrnhPGAsTqA2WTBrj3RNc5cOtp/tWNr+4eYifDO58hZbuPjB0dpGYZ61TlIOj
HM+OMR1XEddea293QuEiz3tqy657xmLF76oa0WdTphxTDQXM2vAbu+7OQbmy4S9zkwFOR/bAySB7
DKZkhCwFPNP/cs+2nI7vCdcJG/nL0qxj4gDG9t7F7Wk6ZElbyHf5SfCwtv3UAtH1D2teeyAPK0PJ
ph6UE6mAUbYAPcB0G1R2ja4vn7mYL25gP026R66PG7JnVSrBVgq7NwlINDZa7draKfXDa3hS4951
fEM6OlbSiP//aMrhNuf6ZMt3QkmhlZIxgt5EHIBryWM5irTm8VJEYB7tOB2EUl221GM7UMQObWWc
8ikNIfYmJF6Xzc10g1tXwtoXFb/VMUY1VpttmDj7ZSiMwr2lKLFQCroEyHuJxMpBggE8VTfL2RSq
tAQVWZq3lbn7cs44fJIZEEyJcqzblXLaTHc0XcnTnH+QNAUkNSQW98/1N4fULY7UwJd1BJJ9Gb/E
qMiADnOQzAfpnhmZtZ/4C1Vx7XUUwXsW6NE75hmnKbzKz/GQo+Q+PIkMccXQPKPVQZXLw7sFGhm6
dz8uQ32PgRjzp/M/WVeGFe7jzEGsvWsiUu/SYDfLtkJWF3GNVFqAGTlP6c+cfRWQELPZLzOA5gjH
cZYYLiWBs9M4IK8AmiHcb1qAW8S4LrcgV8hVt4CDGb8GBuCMvSBLzxg42ADioc2gKn2nOQYMME8S
3CdUZggxVqZaAgPPSXF4DNGBAaiypvwpcgA2WfTtwik0/yQt0g+lg5Rk59z1y9Az/JzSViijHyE5
sHkC86dMfFFfg/eJdwimLrJlPh9TzJaOuJdwexFk9mpsdincJ6+KNFYUlHaDgz3QXGCXIWywFsLC
KoInWSNYQrUZixvLbOIJH7i1AFqyziVz8ZQB9lrQlZDN9UDAw44z7nWKzvigkaGgGidD3oTEurKP
XxDhdGYis1HPoLqmtkflGkAzxIXncCy3aJqMdqUhGgxBgao+LWUKE4LlRaJZSi3xoeOq1hAXWhOP
N7xaf7zwn/ln3WcrZPKjZh90oU39TBQZc67lHfEziJZ6PjvI2yuH2kvw93BwmqJ39e598s/XY1Y1
3jO+gLrRi4guTcA7uhngvElm5ikxfstujQ03tT7FgqXlHleVe/GOyHWE4fsXjGg0obzXxwqtQaZP
s4FTPcTSHFglbXqi3vbL+R//YFgilH5O8dnP6ZdFrehNSvRfIXAK3R5QsXDyArwD9hw5LoY9PGKq
+VJt0Wi/sGS3Q3BMZCyxaV0FgcVyzlOJKhfov5epdyByLdICX8Ss3rsH1e4EUUJfa5ZoH/GaTnq9
JZKVzxqlAuCO/8obTJnOpvjHNjdvyN0HpsduGI91O/zrjZudBiiKaWbJK6L5Btgqq7WrzdL5oBbo
hpPtxelYOKWt8RKBvCpzfuqX05K4DhU1IOLl88irWBJZayi/c3vFeNpVWE+X+lGkyiKGIZ/78AQx
UpoA6ExJQ7kusIZA2+octbzGNkg6gQkVfE3PLMOSxxbQ9de5vc2X10enUjhKIiVrbcKGIN2Kpoji
EmslF5dvEEQxzM9z+5NtB5lqiDdGdVXIJ57H0S8roIqLCfUxBQm7nPXgpi8jfVDriiaEB3erRYkA
FTURVq09VwdWkgegtPqYRg4FMyVhFypM7jayuknc1bBUYh4qJBXcBsVfKcC3Ih99pvPIbbq0RNxn
OsGdB9XThj/xJpO6tZHvAJo9r3oPTDGemYAYl5QzF6qnFrzw1FukAong1EcTM5WsI8Kdh9RkwK0M
GzFyK28FMEkFJ921J3KlMJX0bdVY40y0vHSP1+Qs0P/Hb3isnVpzpJuJ49X9cHAnEc3o/NyuKlJS
YDejfEbCCJBRpdWu5LBlW7k3oTykeslKH8aI9lKWouf2jKilz7TRI+Z4YxKMjMiNOMxznWqqBP3F
SzK714Z/BAfWiCY76m3mELmnADj2WI93PwVFGf1Th9mvD4D2rnXdJ1p9oC+gySmcTUyBGSnZzOHq
VJmK3Tgj2TnF0DXU9ZRaxKEAjZhPzu1z2oW/694w34mjK1srbaSEakjuw1dpNHNqzuLR9c4+PzTx
90hCYEJS6VUDIndM49cztn2mj7JsivBHyz5yLdl86NN0gKuTbXaSFTt5Tt15S66t1mnZt0Ve7PJN
vD8dFbh/XEeCn2RHLFWOntSIMC0GeZSYoITTN/IeYTuM3Sv0KYnQ58v4m5LOjVR1cwF/m3sgwZwG
d9ebsZg/ct/RRJt+QKeR4WyiCW1E/bSWjheV3mKYBdos6A07s/RND9bztoODXSQpeixTvSE9Bbq1
AoU4dbvRxrrz0gG1evrcK2mM0k7//zMYXuuBtjWayB/jpc8iiW1p+EDO8DnxNIhdDrsYWbjyrl2l
YXkHXSvueymp1aPbrzpkTf0zxynvD18pO02WbM52YkHaBMGtW13Fd4KYAcSlrGDRxOieg80VFJEP
p4+Jxb1He0M/AFZdUU5rurXRee2DkDTQKAGu9o1pT3o77PzXf+IQZ/Ilq+LeeFsyTb/hn2PoAFTb
oNxPDgFSzUXtciYE+GhqKimeE0HYmSR0nEDfZFxydM6KCJ0U+F0KZ8EiarKyeafL34U9OgV6YMzo
0fV875TP7BEk/BznLmRVfjd5eBNbWkNa6lacQxacVHkIUrlNhvSmR6dxI8LPwyxchppbNYtgGYa+
3Paq2gncEV/7nJqLhxvX0At8jiLLOjFy4ucdHGTuqL5UzkatOpEbowL8Uhnn3nMZl6lH7ABoU6dk
9LL6pRA9u1FaxJG1GryZ0f8fzHk+UV22NRAzLzBDRWA2bs5gkGdD8uHnrFIQiS22pmXafeKmZ07H
mYtVplmxhoe2KNQJ3RbcjaEt2n+cqoMHCKkLAGNLzp4YZ/sZuDynlO33kIdDz29l0B9FJ2IXjJik
FP46k61F3cEVX9PwIPU1hYDVp1n3Za6ECk6jPaLR5iFTb0uj05/PwXStRTH+v4FSl6BUiOkW5pRa
llUkaGUqvIOjIIaDDJ95ffqdF1RCum1c/kKP1wRfg35oxiosT7mOOOYUE4K2uV53BXlUkGX3zq7j
Tm5TwZsJN47EuzYmX3dUVsb2dkgUmZYPuyqDlkCFYabCCXdTzER3gY+WPM85SLnf341qT244Ltxr
fmXp2oW9aM0BkQZeGh1cKDWGEG0CJFOAgnl3jT6myN4zX7NnD/8eujeiZmaFIktUGzkpkagNNwwK
bqEAKa5yLxXhgwQIWNt1AEcHbJB1vO6GuwIQ/jwPKiyQSYMuwFbI4y8ogg1DbKn86VpuCBI37Xhk
6+TMRDQKI11tP3skVsrEAa4qHafUWvezlcquofZMkArCZ8+1CxrVOs5cdOoPkFVeoSn/AxV10wRT
E9GNbU9J2vujndQCBAv7nA2rHnLBIrSACAWl/cK1EY0fkVGFwQcPktPuUNInJGkPzOWq0a4ZIzoI
la015O+lxc+9aAUbaxMfhsSyu7HMSv1rXAuQ1ugPTLoZHVVWQbzsZ24JiJQeNble4Gucasfs+sxA
dYnCfPsNMiKDH0/dEqqw7bYW/LwwxUXArXtDdU2I+kIGBfPfugi3Y2ivSzBabGhB3IvbRs0kH+iU
hS8Q4yK8EqsHQvvxp5PVN5plPXVrtnsxKc3SZFSu2LSBT+JCC0m+AfeIM0Ha+q/ucW7YZrkKxRl3
aJe2ATwxx4dBlC92SzoBQIZVy3imMeWzsnV1KbozvmW+U8FkhIuSNk1I+pJEqUBTXr8f7sHZcKLV
AjBeYF/mqDOCZcu53Q12YDPV8ZfpO++/hTug52ChZRq8aMW/vKEqGitzg33A2eIU+yayEUzhHBQN
oEhJEn+noBbnZHYvsNOc/9AGVYd4JHFNfB/S4x77C+Ga7ANhIW9kadLAbo4e0qGfTBExx0F/MtMC
KD1+eMjG7AUQp7U4/xizCeablcrrNhyGQ+fMzoX7T7Ix8MVk4YObKNtHsmvdg84D+0kzoLnT3Qvr
oawz6INw+juaANOu+M6EfP2QPTDSaNaHWz+TQMtWCdVTn5cNQ12AkHjx9qsOfhLikakn4XYjOUaB
QoFkcYV5iaa1Gb3/tovX/HdhM9VKqd1ENq9c057V/1qdkISCfwRfCf2LPiu/la/e6HrKZPAseBx3
4TnnESLEhNzz00tdo4ncQiZA8mzA+hej9ItDfhog2diqMiquIdXR8Dh1523m3hyNItURK7BKf8J2
fMPi4T12Afir//X6bFOdNJk78XNU/WPfWX6C1ypBZoEeJWrniO6bQO9iu4sZ5du0PgZRlqoIkALt
zGn0t24dQEC21HV1nZ4+MEyLyFSLDEnJfBej3ZF/wuNAVeCNMniQKJOjNwjbqgr6JdV++ubyc5Et
Tyx9iTwoUwozMzqJ36vRcJjsQsDs8RIwQh/FmZJTUsVTrGQN+uOV4Jw+Ia40hU4VlguhBPgr8Xvg
5fqPN/L1cZca83nXOmff67zx6aHrZsdFBAqaB6gCb1MbbIKCoI0vX58f6plsZz6Aq7T6IN5FStvg
BBJ7EsIzzZTelX5kNiXi87whTzVWZqFDSAG+RyUyAsctbo+AaMPX5XrjhMmESbU8kjQBy5YZ6nIX
NFqobEiW4Od9el6ufPkPlG8BDOqrJ3iSzdCHH+Qt33Gd7z7KQF/1wndIVdE7rxhzM7CwzJ+rP79s
8kxtvzc7pbFIzMHB5NmLnGRrSsDlzeKYeREIfq53b95dV2uYAzenkl40UNcnT4dv+7983Wbsnmjj
P/rdYgaYojLxVTbWpE5yrm1g8LkANCZ+dsII2C90p4uFNYgQc9MkxDf8Devn13kInFUEMiZTf6W6
DprBWltBAOjIUlyr6H+Hqk9eEFifbAp6efLuBUFxqn+2gsL4RFIxlRiI6oVQsb9gKGIvyrwPSDuy
NsC2dKbQCbQaT+7hZ8Lc8soNpCvFT+HUTVrqkfZS6ReLf+mGARgAsfW0hPfp0zio+tZgRUebSHsG
NxWBZnnaEF8lIclLYFIbzUEf1vPu+xlwVw7ivT3K6BXtKVWwYciJlGSGh3PuCxMESqs5dj1RXSw5
Uz5zfhdYCNV9ix7380DzgyRRJvwgMGi/jlWvfN9sKNK69kD+zPfwbD3gXCosDcEwjaV1/0fIKGAy
om2puGuHGu0cXxeZbMsdkRy2OJYw3QrHtU1JXzH4LlEMuLXiN2wCU6Kcz20ZctoQ6KYnVrHo6gtL
uHRmK3y5q6Nv2Q8nK1LXhDCxJ1kbBfh+82P47EyCJFvPOGz5OyW/xlbaAWrJ/zy00lKSEXk6s+FU
YeG7wqBGZv7nwRt6F4ug4uxzsao6pM2388/r9gMV1ZTcHkrkcPzW7uJOXLJ11hIZL6bPZihhjWqZ
yYrd2fzFJJdAem6H0ra8ex8aczETs6ZoLTbtX3GlRQwD51j+1WQ8QqnJgfB4BE7BMkdlpCdgoowY
Iap3+xlEKUTfO2VAC3idTa2mkJ1BJxycEMUlg6UlSpgweBfSrEEqIzfYBaN4U5jr6NGTQFKKWtk/
flEpGBWbYzoQUaWKKA7sysgk8y6r4ETXTi4IE2uLRQaYBurQxSyeSTxzT7hc/N0ddPOsg+Et0FFX
NhbI6lQTDYTO+aMTkPwcQAd0g2+ZhmCq/AB4+bPH7Mp/7On/1OQLSF8oZRkDubTlAr4IoMDPbDZ+
59upb20BLsUHoD1jaRzGtNQOidl3Qyg4m3lZOkV7uFyJ0BH+XZ3Na/fxeADd3iPALhOfUCNX24dx
KMNK/21FmaarlatK1HiQmiKyarkGenLnFjsNoIWMVRa3SX7WMHPgZqmZKpTtUBdQcb+XJJC4A9rF
hf6L98iJMeaAp5NzvLKbwWKWUagSp+plXEwE2/eaoFwKLVtXp8HFYgJ+4e/zuSsc1knVhlcjJf+4
WpebzfirHXaJP/42LV7F1FXuybWtfGi8tO0hwW4ht9MA2wPVMUkVc2SN/8u5xcc4UGkiVjJl+tTE
1MwLRM1FIHOk57BYwTGQngeFM+v8w2rQGxUxvuRmWvRAiEHZ41i0i51NkIV1pbwWT96JKUie9rbQ
wrU27WatwHIyTze+FKjDfoyqg7tOyEqayRRsXZ+clBKCt/RauRWQJmsJUL873q/1ttwl14ZMIn2G
iYPeNkGb+L762Texi4NjXl+o9+kyUkEAkdYYY0Rj4iXCVDUT6lQpEMEaI806YTbGTr5xW9lZPJE8
iK/CZf+5VAvTey0fBDQ48IyKUfUXrMbGqsq+cSoLqPIYagCP90Rg/viXDzW+5wR7ODmtsFY/ks0W
1VsSnt8eQJWycTjqM5TNvQ3XQvjbAqw+f3hhfaziTj1wkNf9lMycFJFLAWPMM3hiQo+MhOhdA4Rd
D+J9kw3erbaL4evFDlB4C4yleSXJG/ABUfFn4soQmqrPF4TtTcGj/Ul665rmDd2gHQnt3j++8HOm
/aubVZhqjuUsoZxmFBeXS6Zf5kcQO2QF/tJI+oRFfVrUGzoT9ZRIkuK8EMRiByh0vfv9FSkAkCQd
W6trz40o+rN320cHtggKVJzz4+//xtAg83bTSU1xfGNRk9VTCh9i1ajijplzUc57LygKk73SdMjg
TTik0t6EXivNimZ7Wwc7CMgKW4hEuj+/elPCJ0OczYhTtL72tqncDSk/imNzYuPuwwbOgn3SF2Pg
FNeFWlIM2tdlYhs6KEM1aLL7t2SjVHJ9RX4USDEAJJFdEWJ2u76kJa1FyXSfT84znVL+cvYMydKP
vojrjVMmjGAqE7QeT98OwaCTIENZLTfcOVrdm/TirGPuUYZZGP17R+oVkiRXMf5qSJv0klBGJfSM
JqydJn37qlK/O17InTr5CN0KAm3EDu2W1eOmdXUtPXlfIHKeaHScuWcrreFHpTKThexvrfYuV/zw
aA4oJtVoBRfxcwZuCFqgt+BlkkpeQfg4vJUsO9YoUSuPkjBrrKWlwxyB2oTo1y3MQocJwYVxcuSU
oF7I1NGQm/dbDdLgb7E9/dvwBIeaQ+3tyDg0bb28QewmOeW6P49KIiYZCkI2cB2RbfQifrbgkij+
WJSlOxb1hJKRvtaRfWQQoculP3Z/QQkfMcVIym/faPx/EBd7Qixv2FZFRYl4LTuEwXUxshbMYaDd
rSuWvKC+wq02LnOCKhUgEQt4nfXXfX0aUWTYlbcLD72wosiDW9sEPrh3kdf4CdD9Y1c9HGg1Fnht
a2OAU/DgftS9moaBwHfWRT4bIaDkzR7WntoXjqNgeu+n39sBVncEicyrSIAv3lNIUZcplekY/BaL
JkjsiSUeWBPcqDN541Fd/v2Ubs3/KZhd5pAu79bCF+QFOGtgSWuh1IY2/KXOqj1j/gcL035Nu1n3
nGJjxhJlwG4z5ArfBC6/FBSUtvQJXzVf92YTdtf/cg5H5Jvkvog4xbhkRqmdO6d5usqk/DdGVW4o
nyRQ8oPANApgc8yQEuNPer7El25wK/z/NfFyRE8hPD5hBNdvj6MiDu5zG7WTL+bKVV0vuzrPcOc4
BWjSfDD39XZ6YM2PfOIu/0z4Q4byqlxl8nyBS9iAK2iGPpVABs93nJEiK+6MQSeB0Js5RcBVeXxT
ivITL6QRyjkJaboTsnL+vYVc269BR7GuB9yIx1BcMjZTqWYsJTgHdB6QCKIb9aX6rpSqQJBvXZSC
EPjyotzxW5BMoiDZ2vPenOG404V730mDJQ6fQgoXcGMX5hU6IRtwQiIGLQBhGH5zyTg2ayeSy5MT
zPdje0NzCYL4JXcyxUA7B1eSW+GH57V4lGTL1aLX8DZMKUp7MCwhBV9qkBlHKNGYv3x00P8jiYN6
S2L7/N2h+9OAVDeqNIKTz+aAnKJ1Y6Qsaeo9x9xasK6OExbg8O0ceaNgYvYkso8e0MK9X+wC/IM1
dthBes7rgd2wrnUjc9PikIRuoCno4WumP07i5gOBqkW8GCXbrVtz2pUYoq6NNNXCXXJMhn01ouPu
JyRh7yDbxAY2uISr2oaJev66+m2tVtczcXehkGm8ErRJqpfcaL7GIpEl2RqVN2eGayVDUiuTG6fC
Ky7Ya+hU2/+L1TSA9Wq+BgQVobr1VmqjY4SZatkgzzL/VdFXTx59jXQcyPBu0/BYH6BfET3nJ5iq
wnIUW/JqITFH+n8KsIQBbnfK1H2sS9nflo4QLxLfDSEdX7rPkvAveXrARqXP2aWaZU2AmSJhE+6T
6ky3mf1GbyPX8yKEqiW1D9KADPklWPWUjmm/1Y5yjko1IEtqBcR2FXHLgxtBIW9Gjq4miQnB4eyJ
DPtkRBADzf2vAQO6L4Z8VIN+MEGY0W3plW67l9S6JIcXEstAyRE+nNKPHEkEX4GbJNgzUvDbyz4S
/f3JGpQ584pkU9XwAVDD2DGPWIhVOA6Y89QjrpJ19jXU88IKp+5JQKgdj8F4MQKPvdQZYs9wxupV
7Yd/KBjDVue78ZM9NOnUkwNJtTxJz7qCvlXFvOyrVXpDfl9zpKwDkUBdRlZz0B4/tNBMG/zeu+S6
TfOBZHejTIiam1IAWQzNsbcFpRL6Q1+GZilIKdRMVhWlSDPo3NgIPQyqpfplA6/hk4Drwp4YSN0e
KFT9cs8mG4QUDMLyMpY10UPwp6iP/zUkf0RGXihtkR/su7UeYi3xpICyx993wOBAi6HZ1dqbAD8D
BlZ5NcZGURwVarFHbfN09VpMIJGeNuPRfh0YFdaiwrZgYvOzA0I4INBpjFinpUkka/ImlO3hNxhU
3FIcD+N4qxAo62IPGG1Oo/ZIgDnU3z1TNGG92NnmieM2D3WLNH5ancg0V0hccoxc2k8wptv77WS5
8bV2NvK421XPr/GzWjXXWxF+t/Xcf1ZXNh0krtD0GLZo7IZD9/RsIxZSLaEhAVDHJoudzNfMwj8d
AVKgBSoruJI6k+TOrWhzRSJIP7OYmCulH5VKIl2ZUDqKV/Nn7bbl5CJLcUVAh97BIoWxBPISY2gc
dYUiLTnm0Xlyzoz/q3OyXogF1NAsEO5qgqls0gS0MHxSiOCYzxMTSPZw0fXNhfYfR2ygZBTMW57C
uEr6tSm4dp1ydi49CCuxRCZATpd1Pq5EfZop48yq9hIbHcVha/+WwAzu8mhYqIeHTsDGJO2aDvpV
dJM4JArD/1lMAH3H2RMKPiTaDhlKQlBdwnrjP8zLNAZ9jhdgmhIUG/FA+jH2iygyLGWphPlyVz5G
wZGKH0gtdaccMwZ1Pn5Y3vka8KhU71zFmlI1j9YDsbZptfK/tH9+Opnp/+LaY7se6K1fMOKcqF93
EujfodPMuBIje1k+DMCdO0jtKR5J8UVHZwQ0jHrFKKy1b1CHj4r8e9uNVuUyu1PmyEs62TGCIXe2
byA27hB7HgnBALy+Y2MJrJBcTh4EsrqndNQ3KgKVflOhGs+qHVxe8OKVK7oYvLWwPdekmKYG6FXe
7KB5qFwCGsr/j+lIdNXJi/FGC524xWs+T8PF995A2uh7ESANWnwaMAV2PWSSY+9amtxwsnoOkNUw
5Cwjse+GjhQgxoHnJf8lWVV09zNPb6JQwQeh6jobKEKG1AWZiVoRL8QZaRnfPVzrsfTDYHqk16n3
vDGSHkKSm3odQDdJbhsqm5X7sA8aEqIy4GcAqI1Ex3uPdWkczV6dvzdx+C/r4CYHxY+CVHu2SUnt
Px5u2Ktnzs3egu5ordVVPu1LS3x91RAiGH8UMdwo24EvLPWTBMf0ji7jbmlSSowmNCxyTaNo43HM
vdKIK/3xGscUav3R+BIYzIBgbwbUU6F4RQO4BgBTFbe9buP8oObZJM823GxPyKTB3TaNb5C1uCkU
MOjH3w3GVi99kiySFsKwUQ+pOLsVUTylJaDIuIF7pH1Wrn4lQ2S6/m/aiTwdKlFTEPIAVfEw0qDV
xIWW3iC7ff0X/F44vVBN2AQHzfntgJmWTFbjtCXyoZIK9Vb1Ib9/EHESGxRGch/zazbXEDqmiwbD
ysSocp0t3nt6BwI3CZSPh8GMp4OAy8i1PhDEgJGQaegTVR+ubuB5WkaOQv2KV1P3EbZwgT8jqFXC
E6wrAfVsn01dy+xTi5RX6iMWPv/sdsSjvpTO5IxGvwYsSfCo3taJeP1tEfKNICPuMJgfEDwJ+5VS
xkx9OwI7tDenRhDE/Xb/lObtiTcCIHxz0/zf7Klt78kVAKZRFhj42PQRhbdPIfRENxQ7M6PK7Z5V
SVJ3+yC9DVeMeykrlqe3bNy62oL4MbUUJrlrwPgEurdN3Xxal48D7t1o4DP6Dh7lngQ/VB64ZgeF
UQ0AjsT2kon7a8pYYefJAlaEutlcgzERFRUDjFeHQXP5ZF0stjrJg4DYEyzWeYg+fZuF4BPA5ajv
wH757N3MK3P0Rhc7NqshhVzwoyNHYByb0I4vvRTEyrY4vZNiPfz4AioA7vLVAjcFQlNnWcE43t+X
m5Jc1JuNhaedofXm+9+0O+nOIptWObWcgWkM8acDlHEoN8YRa5NrR5UAC4iWXGH1Qocv1iR70scJ
oIoHLaeNVLcTHIE/DZwA0nWgGoygiD4JkEzsVgdVvKZ84ZjAumzgfEOpQXi/uswyNrb+aXTzFiZx
Qzly5ketS6+H6MLE7ZYlhXGBF8jUSpicPWZg4ryCM8p8yul7uYbyPgrk2N0At6jGzMbvjMfImLNi
AQYphPWOqCKb/lI9jMvwr9lUJObxFND6w+bVnzGaf6dxo1olRXd7QXjUPZDQbRYWk+wxpehNm0/B
ZlhZ8ahmgmxR4Umj/QhKLeQ0zHPYJGJWzKpIZZr5000fHZKyHmz60ve22LL0qTIbH8K/nhME6gL8
cAwfLSnYjAaWtcIXHXB8L9Tft4I9IVCMtFZdX6wccwlusg7wNjVRh5jrJKNnXef6FoKgImRwuKSj
WZD8nX/OGDBXaBdU1AQ0v/JgVPQ2ftkK0HmOuLMfZJCTRGGh1NJiZwJL9X+di4GJiwcrfQBZ5Krm
jBkbXXVGI2vkcsumHjFnikv/GYqK1luBkKy9BJK1h13o1A2iyesXgd12xXssYXGeyg1o1c8vmcBi
Ro5Lc3d83gpxjttLmz5x5Af5cvBTa29lHdWb0O6ADXBh58/YjEUgTvAzQiLO6S4MKq4znwZYsLoY
22E5pKI5mAJUWTqDpTCqpEC5cPZMUSqw920Jrnwq2OV8oOSJQv21T91LvP5MaTfWPlIlWlfHqj+J
tOnHsgdE3l6a6kZPveOoL7R4933yaITB6ccEdgo3rKErTwnS0V14g4Huca2SGmu8uBDLjCzJRzgt
ZcQkQoZb9nPF9/u5p4Ukd0SM7rswKZY38RrUgcIX5v8XgAl6GYjQQ6TGiAp0gQF55nTzwHer+i9D
pC76vBiDZFlyEP0vPBoeN3Vsf5dXgifdvDUv/H/8PVbrMviFt24d9DYjkFl/Br2XfBy8wv16cd2J
ZUYSlBUO3+oxrPkAz5b416Nh4/lkWyKPaF5X3e0SX0FjlTsK3rPROhAHC3bmfe+GEF9yHDrC91Gc
P65CzfcsJ2oq8896qq12qlXwXdnMrrq1IBgrjFA5b8IcYUP42zSQYXdqAmb5bVne25t+4nz8AYbw
OELDVxaHv0rvzCV1x1J5iIUobPLe9jE5uXdBf27IrYcVIcq7IExEqoOCk+naaQrhamT2ClDLY4Fq
B8V5SsHrB/PfI6fKenbXsT8esMJJZ+mIJoMaX/wmqFOTuEVfeRyumNiatpdgKPpUB43cquOeerb5
XK0AmoQVNexwAOUa3ijLVTnLoUrPPgYKQRBkPJCWaHoX0JSISfbPoVmw/spxrBY0IV56FJRLBlWR
CAFpYjfnNDBvNxpBPBkQBQJzAbsPR6DcoANZ1c+QRc6Ae+wRiV0kWFw9a9M8ecQYWgn3CyXDOB2P
Vu+sj5SFZc3c4YPpzr2qGVtgF5y/aOG0hYbtIMefWurBHA3KYX+pa3L5lzdRTgNHziTPVzwxHd5N
i/99kK55G6QVamxuvL3tM/ckYUsmSFHDvOw+1OWZsHtJE5Wltsd2ogu/jKVfY+hNbe9TuPoIz9iy
+yxDgBW5z8Bq9NOnFIpdc07lPHZ4BEm2LijJ7kcFlVBApF1U7q534LSkZrg19s0bFC5uIydFc87J
YoavEOFIL+CeoDNTAuCnv8jnt6R9/oe1zuvYkV+uqTB2vvQzrNJLmAcBT9bN/vFOj7RTjTaUsU1x
jsrIFynQ5FUdwaxPHxAmCnlTbSFrNRvjKBLVY2u8RKUZYpg/VdwzB8olu37N/f825oX38zWFX01K
+HPkmTgJaKVdvQfe4rmyCcRHXS+tvBMSJ459P9IEk4DuBsFUBGXFra1/Kggdy7MwUaf/V23pD9XC
z6IgGsauIzPLyo8cnsILsyPWkyTzrhBdHzL2oYFuAZj9N3iupB1WYqbPpAsa9n00c1cdPguq8sV5
adUMtm5XhQvL5TfyD5sKsw9rP7CYkXDrGZbyF+zNixUtUb5083ArwxakFv2fgIiPK9swJmHmV5tS
rZPjiqQArhY70h5Vqw6hrqsgVzYoVu+6iWQ1+u+L6K/jMB9HaRitd3zC3+Juct51FQ7wlRmmSnUT
8X4yC/fcsHV0tuCwZXmOaWmcbTJIIk2QNMIJWvAELQ7qZGN5cQumZ6afdHzwEOGx7nv+WOeeAFqJ
JAL6PhvamHZ9oYMPYBOpHG0Lm7RMwSIfT4nxdvMhTBuj1r96ec2B7d4EkUJzofdBzqM10zzCx9ii
rPsVaeVuPBOGZuPQxep12XRoEnAZWMQve/ZwRemAf9Ret3+iLaSWNRH3rysG98itYlRQRu+xJMZG
03Jb+sUojjYyLpOwl2PFxkxjLCASAhsGgFzi3GFogjdwskEGgWqM03JM2/yRPpqJq64nyIpO18fP
jFIYVRcf0+Uf2L3bQOg1f66VmgPThuahxlOqqHB/tTsU806O0/Q3kKv+42XZKYqhIrcRQ9w4Hl49
d2L4WLccrpO7OyAZ8r9aeCw+GBBK2XsGtUmVXarzeQRsRarH359Ed5myKzJpoDBRh8Czb+Cu3TKq
cDmkSd+V84O+0cNKONjY6mZWNObD3W5y3sgP/z/xPsHT9DnRjNehe3Iwz8/frx9XgewqDjWfeZwE
jn6Fw/YyH4UdUUBswF8FAT5aVwDRd7kkUtWXblQNJn6jAd/po90ig50HrG8ZPFAJQozguqATMWK7
QS95Xo6yWRufZJF0sjZ9uEQKYFzygLOiZ4LDV+IjS6KG3arbaSzheHLG6bN9PLhlr4ZirNHFOUKe
5zsZwdYI3Zh3jlOw6OgmqwDnAcVG4VZO+13RJLjKk0LDyn0UtxgIdyoSHtjHSyKVIldaqR3kfZMf
nfuhvGtQOhjPHp0VLjShDaf0qLDRTzEwTluPaLqbULH22CkxPyUhmoCFndlcmN5hHLGEC0LZL8uC
NB5n830OwNkxM8OH5u6NxkQAJC80tHFY7/KEPN1xrZ8ik26dziHpeIRM4vdifJOfkgrCm4ciIacE
qoiirJ0hhutmiy9ChkW+47OOJ3F3G6g8kRb0dKW02/WPkmi0OQzP7U+dMuKJESyszZexcNCazrLW
+vVaprP+n6mNHV4cBvqXpWGTUJR5KbKj+etYiAm6Ou94Xy0aiBTC4xXPA0Icyfaq+Tp2AW/yGDMm
8w8VkcZdJuos8R2XWrISveV4aosOhyky0l4DDB/uJ8Yx8rZ+2Cc7aiaqV+zIWjI8skqMltBq1AH5
lZE2wLR8XAefaWKH/sT72M/WUsvrZEsYfBwO1vfZhl7C6IWcDyoV6LRVdlDANtsLVoFtRXtN1/h5
V/08d+qJQiLbkoKLcC+Z3319kpNlenHFlENA/BcHuNPbPgNrx2J3NrOCx6w8cxuHKoNrLTpdB5fA
2/pV/xUEZkIyCl36Hbp4r7jusR4kHmK8O9JUEYSNINVUe3/NA1y1ifX8up7oK+eAfNhEG5vltdBN
+EvWFRtYxmg+aZMcWxUsUL7vCvFvDosYe/rXgL/2mMZd6fNpWj8pWlrIopf5cRx9gJ6W7MSIJ0xH
yuqoYGlD+x5/d4DUlDaPUGB3ZCeF1zu8PUpjh2Ur5kQlgv6HWI1oJNpySCY/OyGlGTicCVF08BSN
fmme7s4yj3teEoe1bxZj7/iyLeQD7klNK1HYlp3WxJhTFHil0Rs6SQd9MOl+M4OoVZJkPQ3jjR/R
En7tUFd0KBx+MUfqMLdNeq7DgkA+NB9vJB3j3j7YhL4C4Tgeyj8xzZKyInmxVqcotSxqwktkDMQo
w25D7zpeZCFUjnaf2S6tK0e2Y+W+mbymC6lNOgnkhqR253iTaR6wsSPmjHCVfbXiPRTqBGClIroW
a/Mk9Rtnd+daogptbg6ezHVrVpmYX4Iy4k6TcpfSHrdAXWXmbl8cyOL5UGG7nycZqG1xapmhXX90
HIrrB8StadoGnv7YsX0Vph7rCCZcWwlhp6BK3UzO0/icqCT2j8rRRHvJ4TG6G/JNt1RbqnkFWpw3
Vx2N8IG/nn1jflZhOw2uhuTTSNdvds9pOz+7IfNhhlACplnFNtO2kyx5HT9/qpLAcbjFXZlltMY2
kEwMw531JlkIww0MbqE19lFWrcqgRgQr05pGi10/FCTwdzfniF3f6RarO+g1qi146BSM7Og4twW+
IWPjejOWf6Q1sVgmQdOiZsKY3xGDnceFEsaEu7VSajHTJHY2O1OAZrjpWUi889rklemmL/EU5Zcw
oG5iKN/RmNu4OX4XJyNVmgVgvsPwwA0gaJHEjaQgtixib+7Wp5rYHdlxam4JXEZ0DJDDWCpv0wph
CZorgmU/IZmtJZtxKa0M16qbK/BveqOsYGQSratyG5Wp0w5BDGTSyNBfdoAp85Nnz0IcV6RkFOoH
5SAQ6YCvpQv0SCFZa6EV+Y806ieNJLObh0eTdGmpgJcczsfNfFc5BkeOYyarSorCq/kDUrB7aQ/v
VCbNHpLHPK3IZw3UkArprUiFpH71xSyrsrHaTESIFmMoeC4xpp6fARwY5kXBUEbLFt/rlm2Dsezy
5A6pzmSsfvd/2hnu2bYRsB2unqBq+Gv3H9MXbfyVamfN2NBdPuSW5i38pYT+yZnTvn8Qbnp9l8xk
lMroFYtV+r9Y07994TQjQmfduzdHLqTqO9dv+lZBjzMtsmx53vLVEcdgju0k0mVLK8z079qZMtnQ
IuCVc5x9PMJrI9byNmR5932wss1XDaIcmhTG7nbovEWCfSJSE+d0ZPoEjSnhd7iuozUi0Jqdbdji
/eZUMGWMxAFK//SxFip+vS+9pa7rVc3yoV/U/tgi+jsSbDW4qbFYXlxv4UfGwkh0t10/FVP6gyOL
/KrFdWHoyb7NBCckUCWIw5PpX/Di1JnuYO5EWM5S5aOGlUU98s3BypgHC9r5N3wjH0Hnm4mPQ3Dr
4y528Gd5F7Lso1KfPM+iqqvWxpMo358jGSA2zGRWDEeKOChdbyorB9PnDqKEKz8GoNoRG069H5lP
PipkUeyjTE16rTf5TI31Hec2bD6SyhS1O+i9abCZM3uUoZ7eEBnSVQghR8CsNuqIzsWXfVLh0pP4
F0NM7UmTegqI0W7irpYo1PxFkH1Rqsk0L+gcpN/lRaTjIrrrBmlMjomqvOPhgGaLKqWybBlmatJ3
rLBNmnt2Cg+w7hsdNIkz8ArDs7/J+ZC1aHb1z4ZX2KOGjGbhgFldRnhLJc2M4m2EWGsx3IchuDZJ
DOXGqPeGV81grQmEMzQYwxi9YE1dOCyrWx+tcBy+uGgPAhZOlHQqJF2T5mV/ZlPVL3mN5EHAw2Cm
fIiz35cN4JQlg+LIlJ9pcdol2Yx4uRsFfFQdwi/1ScjIcuOn99aoJprC2HlOK88DjWN4pLVSGLaD
giW4bz54mbBc/QcviZqG4D4+s3kfhrqOL86s58QjGa7FiY/baUk9yvjaP0mG5SaPG7X3dTijGAp5
dEs5YEcZWR6vAwUFaEPeg05/ObJ1ZcHtlT6SWfE3c5guFJm3w+ZRTah+jOteKWAE9lxrMfx25y28
5n1Odxvij2S+MzBHgS+nXEUVuL4qw7UutjT4y7YY7C5W3ianihWZaawH9/kVfeO4BXn2DIISONVL
BOeQVSpsZ1uvqtZ1hurfOaJXm3QAkUjv1N7zTrm34O0YVDOcd3gxkCHqSfdK1OozSl3M9gArH+p7
BkWCnKxpB3RnV4zwXAX4ROdFnUxcYdOxK7YcyiQGOj5eFBz0uQCPT8AxYpwR5sSgRFNk0jjnklDB
0oTfwVfMm7U1Pyn3zwPnHfRalbLuV+zkcUQN4C8GbFoiYkaTYXYPRDHPVMwMpTHd2+LfpSXvFtE0
9/0RWAwt0Dt9VG2VSuH4WyovfEAtGf1Ug5nYEAC/ySc9biVhGXvtwNfEXJdjFmp/GP0ctfio7XZC
L6lPmtAwkOrPB1l1OzxsDteSqiduQsQqNxPOE15IBuBofXFi6/nEfrVSixz9QDAXVxDYkcOMJw88
XF2RFwVMftznVTzfQCZAcWRxIZEhKHMbI2zeNWcdp6w3l+lC5Q9dIw56Bv3Ys7JqQ1S3lqC7wS5g
HdKlb47XyTKqChKlo6dTC0tVygSF5VLvA3n9/sO5vNMLPn7pwELZEPhjXaXe2Ysq9eAgnuBCg67d
Y3nUSrhdU59P/xEFrgxrLRWU/1qdVxS43KzOPfCVJdJRN5JYg3q5KUMyM2KKPWi1sXgeBB/6DAif
SRzzGzAQJ/p7TamN9C7KL65HiLbTVq5NY+05NCXpG2qoMeNOLgVij36/a/nE9uqMsYZcB3VKm+qZ
Rci7+WpP8OL5C/GA/Jotc3P18o8NSsYkQKC9Rxf0zWH3+6/+/fYHAAM1W9x5OLQ2TGirSuKiZcTc
IX4sUAbOJgD/3BLrvpZFucYUmuqOQtkRIuv1EdEZPEwdJ4Jwk0xZDU9IggtfRiLdbq1U6qHZK+3M
Qc3jSSyI8vI6xdcPausDYSaY6ANT0rI4tfetFyAjl9T9SUT/yN04NJc2+P0y9fLi5U9o04feQqg0
xo6Vm2f3IcDIMrFrvCyP64aCueW4iL4jrKhtSn9DgdWviHTX+U/OctaX/heHPSqWYBwH6ar3GPKq
Sx/LxpP0hZEP0N3Pj5qSltZVlSlYZkqTYJhn3jdwkxa/4gjI42jYyG5WT5l6F+oO6FqCv5R9ibCL
Fm/NDep/hSo1qb32x1T+DPVS5pjE39d2D8FruFB2RhpBxUb0RzpvWXifXYoHDAzRDAPA56kECbaF
Ogj15iITzdUKqD82fLk1vC5jchKadIF4LANJ1tKKam4i+VpsKNIoVLjE6CHBhK8m0U4Ca+9g4txO
+RWhVskXf+2tC377bgo6SlhDYTDit6U/XG/1jOqsP5pMT0oh5asRhCeqnLq1jj0jvNLg8mdzTeGj
dqbbUXLeqMFhKbcjBwCKyDACl6GW6mNHPddit0JQ30gMDMqHEHCqi4zUN46/l84zBMbc7PNVad+1
5tMEGiSNmaWt0fxqzxhBHYLWpmsZV2ipJtTbcRG23i2+4hPo8M/WeytKJBppEcR9zsQObsvXD0P9
HphOL4pNDH8Hdshodc/yvD2zKl/7jEYwJp1AzKNKIxrMJlDhGbzeKuELCGvtj3bFdN1Oxk/jyJA4
+QdeiSBDRXSElhGjhbik9wVEk2pAlfORlLjbM3Z8OPwfZCSY39hoIDvWsuIoFJq5sK4tS58edLCl
1gnJPm4oN40KaDsr+U/UylO2uRxjUyC3+f0JJqit6gVhHcKqwCQTqkdHVdKxqHHoQwcxFz0g4Vpc
wLdZ6t1UhXaE7DBk/BZthuP5jNo0VqEVPBZwNuvB4QvCqpOFRAg91dtHyV5CUjC7w9CtaQiWb+wd
wV0yJkF08+CRUI5wYuo0fw7aluLF2onT5gyNhYoTY3N+EZGfMW17X4SlR714VLe8LnU7FLVc7pBQ
AYGI/M4S6+ob1jblSfuJp+rAiAvOcLrQhGnAl7fnqmE/3qdAjdci5ipNdNL6QpqY4cmiUSK9uobA
7SheZayQ9TXfz6mSdrOyvIGVW1aAJwRk0dR0AOWUTaEviLYJCyA5nNP0gOj1uUgWkP+i9hB+TNAe
5DvZHo471W4QtKRXdqBnyXIsDd2ico2iSPL48oyrXYtWULex7afRm97Bqdk1kf6W4lLEnR3S2h9S
vTtd1aisNy8swDAJy38tAZQqT26h+q8dqYojWx2eCvWnWbzHGcCp7pk5RJ+3CQTlBiUr81ZsJk22
thblvbqp08X3nST1BpGoYVKIkNOQ6vtWsn4fJyGKjevH2WyLuUzWbbyBMq0u856R7fjpNr1iGcMe
JZjyI9dde/8lwTrD446gD2hQHBLxzIUWOiwhp37LU+RcRiZhyV+0U7kpaoHnRjSY166NHx7UUEb4
nulHzSSzgbt0Xyk8H0nscQIi2/g/rWXs9KkWNZ1TgZBb/3Bzs4p+uMbTBETL3MaB6MZbp6yW9HUF
p4cxxsfiKtpxmlmfaeAqc6Xrc1QrABXwuR+FhgmwZs5NqymCGAgzJ6FNOxnXdrnp4WcljNzX8pck
lWrY5V4CxuzMbuTafcZ7EwCVslrlnW/hjdYv2WWSPfFV/UB9ZscFLDEo5PkyGpXjhLiHVrnZIAcr
ibAk1XY/qUkaFkFTxneMMUSF11nqmNt579cianmDI+KMLMovSPNxZYji00TC/oi4FfXV0GugYZ0x
moqCdPEnIhKllLJwurdGaWf9BcsminuNn1EGzzU+cRFgCNjxooSFWlO4oYGjYDR6IgVRLEoLjcEd
Pg0dCh8EuIIKn0jmkQSlvzxZ3eG3AdYewQNkzfXY+70AfFI6wZY/JNG/5BOom7XfSMJpW+RPnnFn
x1PQmfSx6N6/xJ4wJ8wPI9LGPNDt+4mBCEw/UJkZQB5+HkSk+YrcjwGe3le7trvphp/JzZHl9tFM
rhnDUqvmm9Lje14ZjsRG+5ujbF7nNBtGk7Wx7OkgShhutW1DIyBmL+yOI6EzlkGb33+wzj70o9cb
fCFCM0R4GwlByHW6irST4DqkoLUnQn1AcjOjRB1dMyDJ3BnAZKWLcxTNQXms5XIfahPTklr0cxAc
+tj2/gzOQWDyEyGWHQmqf99V5pJ5ixIo2Qr2xEOE9GjB3IWh0j3PiadPZoruyNi6FYaMeeEIG8we
k1esCFwAJbyKpR9of3i7HyYuhac1NhfXaLR/WCP5t3JcXez9Lf9iYZi8Tvi41ItHa1UIc7pctTHJ
cOH1x+k1zwE4g8h7vXFLsFyI9rQPsXjl3vHo889q7y29xADp0/RgVVOUODdO5lRVzc53gos1ErU2
/UnnGUeRJYuU/tvA93x96IxBmA5Lv4kRR37xQ2CFBDwiyVk7lp3kGMa4OLgRYvZJ1CtPHjk4+cWb
UCkHe1JOpnJXCAkUD7s7h0IOnikb1z2G0T6K9ae8rxu5AqzayJGFZJb593n9NlOXua+rnVETIlPq
8rjuRAoY+lHbZ80+OePWI+BzF685naiv6Z62ptaBZ2TA/y9/CZR32F5DSvh7UEHn8FdM+Gez1IdE
KkF8kzBnKAjKVk69w4Uzg7n0Ng6l8k8TvhG8K1WnsVrz1Ji4vs+cW5jwEiOJ4Ipc59jsTTDubsJ3
owrASXvL/3MRmQ4En6cGT/kNzlRLwyMnBSzpcsQgMMZ6OlWMbDi1xLr7WUJQdL9vMn0eI+hsI90B
ff8ppQLMO8Wh7SBa6WxbXmPdBrzlQ12lAqX7j52uXdVxtBFK1PHVmfi3eYAstwiIdLTztSVt+q7p
a480f52ONl/0Dcd/NW18QZC1ZkvcwGESd/CC8Q8FOLx5+0LAI0rZaRIP3V1LHUgUZejf6CptXCAz
KBA6f4a5h8LTBc9kihoqsQRjE3Nu1MiexlVXVTuYCTn9gTG6cv9bdpZeRn0EisBXL9GsGuRbW6hO
wKAQT7FGKCYMltmYNdGZSOm6PpMOZy19RwZmp8X7MBA2TJ8LwycZXBR/1BoHmMuYDbXbKHEBZWgO
HY2yZTru9rxzc6zQQwi1TKJ+DPJUEmopQRZycnJPw2N4imPNhcuC2ZhbaCijBDdIVY0rnrqJUtDu
SlesHmeDQPKqBXeCwxe2pet5BGe6qsJGWC5BuRA7JV0YfztM1vWUvUGc/3p8/i4ebYLGC0xaNd/X
t8R43/aY32qXa0RepmgAAzHqZP3hjfU9V+tKKsNGIezwmNlyBmeztrpaXMDiYdeyb/skwmdYApE8
tfBKiH6ZO38iNr5LevXQ4XPE3dOp2/uX+H6WAcTk3VPTQz0jjhDQTZXR3hHaRiHY0rP3Yy4otvG8
Awd2+5fkq4pM4IqSFEFbMCEvxQiqx44tWl04nG/8Ni1OzNxBrRwjUs9OR5ocXoxHDC6t5Wg7+FDX
XSXoZGK6S0KZ9Xw/EJ2zajdt6YVI0h1X4255VLtyS41ZJdzKRjGCDTZwlZUCX+KDOdMY89dk5ONZ
+n1r3iqas3GCWQtvr/0zj7t3P3LihAoSODiv5B1J/KatD2Tny6sYMHFj7lkD72Som3H5MPavqqDT
qDFXsWDsUpdhGCJUrbCi3Ee60Ujt/dyL43nIOGhf1FHebIZNmR16IA3037czZrXNH19wowseyTnl
XMsSjPUHQ8IiIbDDW1fKa46w6PsInHNL86M7SNXtXTDJhlXwKmTmjKQRqBXoNtYQ8rbupqyVAUMF
dWl5HOWu0kWwPBqBo7qBUbsQF8kzPfaVqLnxSRIa1/oTF79qQoekbvbi9/fQq3pMxa03JeWDDo//
W4WPouINbj6fb0C1MSsLpRMQNg1wjqVXD+xpVyQjz0vef3OmlMkG487miey7N1ixewQ8aje/8Jfh
YSH8YaX1WJ1IscfBWnERAnUxxNxLBrrpoKvOTQFu6pPfw044TwZt68tF2S/YAbduntBNkGNUcHAM
dd0OYGupSTMyeoKpoDkO7b0qBF0q4TktMK1Q/YxGmMDn3JmtdzdNZAhmMLQ+4HA89Fc5GXp2qWP1
O2nclM1po1jykC9amC4IYW8piCUZRYuAcFwpqZQcZ5lDXB/dK3doCPyXrd9lwr4qnu75DycDjHas
I0NMHsMiZd7QO7ZwdW7ujlJy9knEAZDyST/Q54xEB9bKy7ZOiKtQgqMjJJXRsOAc5iuLCSPARLb9
F/YMH+fWn4XemfF4+zpjxffj10imSRZnPQnAksAE9RrzyIxrNWppLojCd9vTn991WxR0xsHXQZ1+
wbSP2wzpy81VMYuTVyfpThzlNOUgxdyZebEsuhMFmbHGDRlAdY6S3ZOBwyCXEvH+697y9DbFvdXg
dhXVSUA8FUGIBZASyT7a67mIkMfEM7tAUvXqg58oTNCg4CFO5CgEcF8+eZw/sm9xvD75QUXVxVnH
BDhw7TprhvCdqSjczn0us72LcxLvdIq1UMZXBr4lUSOwo176uAhLZdNnYpI30RQDCUQVrZgJAxvt
8pePEuQFTHoAK7Ytr33NWG3WZNvhia69cN4arOysGQx5UO/jMrKioXSUzPEfLQV3YBjJY3b6IZvG
8fPIifQ0CF+tw11w2PYdRR8IfY9wqu/vNnxc7s+3k8aYH/ZoHvZDHqbvyD04M//fCc4QXliO7hBA
FzVz5GJ6EVTa1GiKjMOIQYHacgpq5rKFoudr9A6dTWlo5N4vF3zCY4ZQ3sPxT1Ks2vl7rt5ZCBWY
3tBtVJAsf/6ALMAG52tVAt132c5Fm7D+Eoju9bc4L7t+O2QDJ+ekWbZikF7kexh5IHKhsyxyAKp2
jF9ByiCGHAP5WNcjtFo9Mvx9A16wOo0cWWf6SRh7FgXI53u2cY0uCAGso1tLkJcaa+nNDYrJMlzG
KYIqx6NEutotBB2hXffx1y2vn27iPFqI6RuYPk26c2E7Xa7PMAgxLm7pGMlybwNmLOaxk754Xpav
ki4LEx2Zj6CEyULBP7CsMxF1nYzk+mUnOiWEGImSX+mXklW+njt8vZMgm606bYmKg+IPcqi+zocT
ktSRdxhsoKutKCgZfvcktOPxyNMq7WD91UBadKTaSfum70eqUHjGh/vUPY2T3PhzbYERYW2g/tLI
1mpPybQ1kudhy8r+7zSIobhUJSo8lI6Z9dZw2o9IxxASJd4D4o/lFUmDWLDHY6BMdt7ovShMw+fV
Bxhe328FpMtyhZTjgIeXjXRu53ZkFF2mBmcaadfU0A5X/zRz2dV88oG2p9QsxTUqMUw9jP2lalU7
M23sUxzJXlceAnpjviKSWuGi086MF7gXqnGyFUbOduGfyGlkD3P+g0hBeOaQIxy8veJl38QxRL9W
fKW5tmVK7t37tiyviYIHM2Av5+6H0Kr68wyRzOdwoLcxUaghKaWQ93HStSVarVb8tqqsFuzI/pl4
MJALP+RRqzF9jOAD8lq1MuseHT/H98I2OXUd9QFkeqq/wBS9jiIBb10MLXadwB03cC11lCjKXwhk
0PBxmpeFRCzn3CaUetylwi1rz9rMhn2MuY1wPFqyR2WuhegmnT3pcInqtZ58Quzw+mTxWKKuOPSq
cqPZeqGfnc5S5Fle7EJFjjNw7RwpiiST8rtoaJ4J89y9J7gSpNCZZHh0ibYZow1MQqqczr0NRkcM
GLvBeI8DoKMTJUZAAMN5AqcXzpgKV8y3ZdDGEjQqovYMhc3o4neOlsd3HFhbER/7ioiQ7NrJH9Rl
nGA5joVaPOM8q2DLkesCnsZBOXUhO2hSZdcA0M54Cxo40MIaurq0KBWHkRU2WfQ16Pyr6KX3sqAF
Xf9yyYW6FBmbf3Liy7AsiaBnQ84VEa2dMNPfSTlpVs8pQgPb8jiEOlDEcbIljgELkD9kWxpU0bSQ
WmC1kynlUhcyfNmHTRwtknhML2x/+RmvSVHCRqtxZ6+UJ3b9DHmBX0cXxLzM9SsEGa17KDEG45NI
KXaX6eeKGmKjlHsQ938UHGZxFUWOe5uJTwlG+OnPbemEp9zV8IGMmJaR2FJl4GcSegngZ/Mtpmhq
FaLRNKupmci1ugs2/Wv8haqXBZCYGN2TuwRTSFPBRjJnSstC/F4pBM7aob+uvW4D6HSN0DzWHmtH
9/B0ycOvh7O+iyU3P0k74WlIbgHH10gfqo+/wWrToTVv8g6yXkgZscCDLwQgja+7v/EgA1ID36eV
4flGMIhHPawfztXbkpxvW0o6Zc5ItQNXmVRtjucVD37BJA5h6fsx3GRXO22oQkskGi3jGAH5c1Y2
aVFu3z1bploKhlU/ebmPkXcJl4sT0FB8+QrB0QtxkfGXiUPgmqSIFbd3MlvBSYGMRbyjM8qIFwoj
iWW5zg4TMCHXjEBk9nJBLVlCI9pqBFFC6nacn7C+OIgc+T2nCOLR/0Jec2ngd94XCdDBdzSCRlZY
DDGB9+rHcylpQPS5gGVAgAr+zTTuH+T5+sgsD95pGGs6hvk3vu+KXE40mFTCgdgoCPU3b3pKWVqa
tyCfz7XA9CyCWE0h8QZ36HpBj/sSY8P9i9MurysdlXLG5j5QTe9y9ODSqSOTSmqdwpkeJdlDoN98
UyAZjlqOejWnp7bASQkcHCauTR0PbpFlzIqEvhyrWapThzwleHuOKrBeIlXLWk/3TvLCNMagTGRy
2QtygQcRdzM0PpHrOWpN0QsbQLdacqt+ruFkvrTP9vRBkE9DkdCQBEyZuJwUqsCHJYrxhk3cBGEH
1h+WR41WX9uCp+AMSLGBRGt1RjnxfvFFtDPhcfye5Ql6vrjcez2AmU1H6ROSQam9NyK2FWA3yKxl
KdUvpGAiDv/mNrI955hl2TN7KOGaf3nzPfNKLvg+0oj4as2IIoHgiOnQniiRT8SVy9HBfqQhlzN0
NNVcnYaqg9HYti4b2cYQW58FMg6M8ZB9W+lgPlDw8nULvvFmGlyv0mTUfwBQp1nBw7a2hMHqyl3t
HZmpFw/+F7FX3s/aymqQ6UUBiW2BVWAJZaZ1mrH7AIWifFs6SyhOd1+eseZas0qTELXapjM0I3ae
9xa4+OnKep7DT0iw9HFS13hheqauEBxNIUHOi9x0xNddG8gUaWSS0sDfgsRvxFv9W2cZzKsYphE3
e0/a39L2zR1CPBQTDfDCpRxzOeezHdQ00abjuWW75LaxPfyKtghG0MIgHHy8N/SqoOuhZB0/EW4P
rRMjON6MX1CP/7b41kMMwUGiUOF6nDQeQ3Hz9jPr4YFaZxLxVDGU5HUbUEAtWf/a8lDrs4w0F5BX
e3cj9DYbrQ7qp1VI0Ltj990DFTafds+8jMi+Q5l+plv4jcszguR0knBJ3ERrQLhpyDpfUkZOuehi
ztgK4XcY+ldEU5GwT6m/Ip/BrPKjlJDR4Tvvqlh6ZUjCE8zAHFvmR5zIqas2lS1V3jBEWCVzozXf
zPkjeSJQtPn6l0bueiPpFCFpy3VrFtpwUmYghlVyLBkmUngUUFmvHU4vXdaFu6JHb+9PCDU4e8ml
YC9wnFSU+wQ0Qb/DMxODsVmj83dYmm0bqaZqD46U9eFXCgyYFqpJHUYiNy8K8lnIjhrkFOu72bYf
Hi1956EAfNhGMejvQ3LrzUr3zf4BBsE35LQbb5KlAwVdu14qoKhcI1qyNH+jtfGOp+H9eiK6dd4F
qUey33WskmmFdDmzlcChTn/H19VAUBKaqb0xl5PA2aRhJrQR8CF1WkiM3H2RI3Kyr7707IWB+0Sf
88BGL9ZQNxGt8b9QXqWNJ14fh4XVrvK2ZjKNcpBhYkGpeN0+evJ+t5/gvoZ6XjREsWo0fOxYuwZH
zrcnEBYMDZgR4/MNQ2A68fapLIOWA36ftAh/lh1SDTJKCn/1uBKr3k4qm2FnQ3MUa2x9/gk2/mIX
AzAnmTrHIf1cH6hsUv8LyT1tJRz5LFCaXSD35JMGcQM3T7JNh2KJScPiU8p7j8GjdH3nLDql/p99
i1TIdKnb4FyO4NAlkHxh9JguaumHhJQyigfx3TppTtkxiCLXUA4H/SYA1MWLOe5DdqierX5WD3qR
YakMEDQY6YQrvB07IiFMx7lnbNDskP0kMLqOC+GcdDcgRX7ITy/mgVm5Lyx7tpYOK+KJ78maVBW7
X7QONAj2kg/tHegbiZIrYRrQu4x5sPCWkyP42xGv1YZWwDAZbC0YagsvuyhMtBaGYXNOiyqfT4a1
xN/eiwOp+A9MFzAzoiuYZfjT3owrUf/R6KzoYeW6ymLcXLtoJZGqvzPx1Iyc/tsDUZ1cjqx0vlaz
uyQ1d2G2vQHxXkpprjn9Y0Y1D5yxfjRdgIGVZH77aIrwvZsIANe+wvPRLTu1MrWCucClhsXaE/TW
CMTpaA/yBfstXsMtn51Y7NZZ+/BgFSRpN4OLT+Eg4+ChuHgiX1sojoSPUFp5bRXs4lLYcExAgamg
mwrt1Z3je8m+GQIb/Tjdo93C8AWJuK7o1Rer/7gB1nThWKm7HcifzJ81Hyt9Ugdow6Acb6DvPzXx
MEt7+H03i5MaB52+Cm8nJZzMVs2H4vr/FG9C4hNGuKupN1VDpDBLiQKeU3E9V2SNCNL0JIXd99gG
L0LWif3fZDxcbmR/W7lBPYBsXYWNsaFE5cb0jrm0Q5FUz0R04KP9iVpybPZkzhcyDdGlNOHRnaR0
9tmzrWbcrXmapWYHP3gV4r2Ml9cQuY2xr+rP92o0SRJTTMyJJHOrLgtR+ek1WcvMZXuzU+0xpoVg
2GyvSVWjEXQR6wRnzIDNs/j4a12bNurSDWxBLWB+gm71S4IOPzIMYI9URO47R5DYVeNVXGxSjJIO
LvTqf1PH2aOnHA0pnUa/OrG0grqaaIhSLTeMr9mMqL2vukY4HTrxJUBSuOpi9aCQrVi4J8BhBPJN
L5yQBahKO2JLOLe87oVG4Am8gbmncjOhCdANMDUbVDK4KMINwCfPxTSP7XFKH1eC/6w76eQHeo3Q
IrBXqj5dBBX4od1FFd8aqTgt5fNdzwStRMErpkgu4lfdpzCtle4eozmCB2ML4qvx20R1J95QiYUb
7UIl/B+JbhwjgM7vTbg7qPUGpvcT0rW/I0W/MfOGb8522bCCw5QAPZcqY6OynqYK/OWsitY0ttUI
z3DDk8udxFOpk3Fc/gWvIXnhWWnKVfd4cIbGCaPdGUvQ3m/tR3YJTeuQYi7MsQTHV5DnJwM1Usx4
MvkQHhaGnyKgxmBcPPOwqoBdfLG0BEOctUry2t5xYKSx8lNfgfOltRDnDeKEq0py+PflCRH9UCQv
OTwDQLZXkiAMXZWwQ54foJgWnV9k7/U4KchGOG5/8DmBH2dmNmF9l0DOk++R6qflnK4Nd7U4PuyA
fNK70qxcNB9IfrDhD0crPLAOjmomWDK23griSeGRIlzKNPS6LfWRjgZZKu76zFUJ1djEsVUI0U8G
IebI5cjaRguM2/psnNPXaKk18IQAmL4kbjPeA0qqk0y4QAQsstcmYDCTwSIANK0qZf7Hg90qhUjJ
mGqLFJdYZrEQmNUlNIn5Z32ydhAGwtDxD37moTcps18ESc7sWBFeKYO4cNpttoawOqXajoqCq72Q
S+I7eMb7/3EuQ5kaHPRIeLBejHwVPD8MLJE/N53fQFFgR1OsCAyMq5aMqDwU0nNLmwNocdR4U+7M
Dxbs0eULkQqinwdfemvtEyQEEQPKuOwpjvmVXOLRznFsGJRAP5ZTEIxCct8n6LRIoYIzHb9HPnIb
I0py/YLa9FrSqnT5AaRmt0M8MIokglUSN7qfWvmKOY1hIGrraeJh/8kt0NMffNYzwXH+peqKBqa/
QNLTtI1O6Fy3LFtMl12ume+A/WB8QvDViesWi6HlGn1S7tmD+MDnR3mNLdqkAXi3VLTOwtejx+1q
bt5qvN2uIrJyEA7FZ9Tow4oPnGH7YM5AkYR38sm4NmnZowdeu+zSCcE3RLRd1Xnn1pdSu1SGeyKT
y7apJmjgC0HrlGjEXFBx/H51iYxc5S6vl45pSO2NGVZus9KH71J7ieYWWkGwhlhz3ibtVQemTZ0C
wqbyy8/O3Hw3GLpXaCbRK4Ue1QrEdBYmbLV5yth+Fv20aGVk3WI4Bg82QefbCb8XVldEw/WBuDEg
YzPUq77GqlxHNTFozuRg3kn/nvwWKi86kw2KnLsTWCf1UCd6oUD3R5Ihl244V1F5guiwgPYBtZyp
tcCv+jaMwq3ccBtTtXz9oaI8PqoelS312JtWRmrDnlHKtghgxn0sNx0uKIyqQAPhJziHOR6Zo3Gm
C8/3Mnny8psXB3jVXxkcsyUJGBDUM9q2mN9mMuXisPSPFimaOZsM8tXOURHx+ZOQpEhM34S3d5LF
eztK0j+EsfvWI4uShhGl3lGGmMZLaVwZARvIUdX2LqtXH7+BTjxcHiZLJsuSOm7p7c7w+Am4dJbc
AGk0rQ4HNfE+QBs+pEpwx5V0IM/wyT2mfilJoXWieZ69YGjGcN8M/valU3j7BW26sf91SDQdUwrn
ikfPfjFvcDxZGLQJVayTnr69kj5kdpZ5BV8uMNnSrFqwW4bZtwDm/9X/KwxdxwXAVIz3cIdUWLyC
GQZ2Dt8cCMmvu6MekRhY0w0jhuejOkWHsR3HHq9xP9EKcPJj5NtX2Z1l+2UZ7l3Zfr5SRPZeTzE9
Z5lAiBBVrAWjil5Mc44JL6hG7W11vmXYPQw9t2/rCY8zaRhfo2bVW5rikwgo88PQZPGGv0Dq3u1v
0mr8ZBwctpaHVmJyrV2ZWSJ7fxSQU2dUKaN9e32TnMJCSLhdUfTAtRLP162jym6ZIkblWg7xRw4n
b56oXR8ctnph7h64n9VgBQ1n/6i5K7bWWxnuXfBa29k595omabwEfC/t7vPQ9tDQMyJQlu4XoPqg
NThJ6DucnUFCNZTcu0lDu5z49aSQ2PhlwAAZ7DsFE7gXVLVjn8sX9kzgtM5hw6IUaFEOl/Wr0tyk
20Na2qiQdh1CbKzheA2RA5V1WxKCrqk4CUOjBcuFsXJRR7Wn3/uVI+5xTTufzsX932GQKtFtyyAU
Dvnb9aEVZYgvTtEoVKIafVkcQqG6kCpaUqXWpNNPoMHU5vwHb0X/zTfoN04Ap09buVt8791BHZV4
IIHjmM7USgQCbvG7MWn4BFA6gGmkwo0StR8X7ULpKK9JsBL128r17Y0wM/lM1v6v7j+QjaVzz/tn
9eZ0v7JD5gD6g+zYsscf6LhCtD+7CnQ0YvsWW3lm5S447af5YXGdg7f4WK7BuduVNBpWwhDvRYGl
YheuZcXO53uvcCyhkmuO3wmkZuze5tnl0iLiLrrwZpnX6F/kiCnuxVSp1uFdQaCbcqHeu7VixVpH
GlHmm/i1GmHECtmaMO/V+yDGqE++hjFLh7BkV8kEq+FkLBFrnWvfXLUFBlZLPfU8C6eI74UBJOuH
fH3nhUlmIvpLM3TJ97aOlLQG98opCFakaO3JMC5d6PQUVsbuRQz/9SVdPERKpBZCE7VcM4PXpZcO
GHtDHiw2hB57xxyn3BQ1rGWpFNPcssbve4sH7hvATSdb9so62sYJoGxDQMA9Mxwxvyxe02kRnKQU
vdIFn/o72n+DifUKXCGa0I3y1r9sDuiDkvigEVchaRwoJam5R4DH3D9BiuaOiuH/NDs0O4VJk6ei
DVRYuqHOeNCNRKcJtPj/3TyvMJ0IGX5Uz9QWMoXjTpSxhE7U+hR9N9YJSaW5C5WSbKalvnJExJ7R
QdbeqUn63o1sci7fKPtq+loqSMJR6LMvUWC2r2lWlodytn3LIlBhgsBkAvURYVsWACCOUkaPRobM
NMiIAzrLI+KyiCmWkyb3XUcfN8TavNUfsrnAcg6eFiiy3+HCGyZ5K/XlKADpz+IU7f9S9VF2ub3g
1UaPJ6PVAQLLOrL8Gwz3dBmpXcn5QgwE1VcljSVnvKqHs5jbHzI9fGmrmohCUeag52ADrEO3g3gE
V7gD5oVPaM4ix3ZQWbiizlgVvMEnv63wll3uzOAh3VugrBTMl66RgPjKrmpW6+R98Ea3026n2tVY
CKddfIYxJo8XaBEX6hxnq40Tjl1Ykzb8D8k+PE5ENK6c/uqyII2IyFA/Kf7a5i2InYmPYrYbMr3J
X++/4WpZYG/+WDtcXx3WJfqJVfs+HTW4r8cEZMcMKm7vxjnV13AMPnKIsa3353MLpwNtXaXyEQfz
HI0De1BDR4vEvM6+V2bOOPYtLZO9RumKwJ4AagDh0BDyYdNKy9P3oAEQPrL04L6DrMYClvVtSoEf
iL9NKTxsRjM/urEh3EO4VmBu/ARfynULOAdDo570q0r/N8reUmUAUnexK10gJ132qQjPeGZzrfAo
3xst/QwsbJOKLzIso/mtvSa26bad3dzxB5mZNGwXEgIcqBn3Lr1RkYHYSKMtDTDTFeq+IXMLVo/k
k3awlOEp9W9nwTkCSY8SViBJ8kTTuNomeSXSjJBCvtv57Otj2sLfLQORq9FtlSN6ampJNBhBnpn9
40D+BK1VD24hoczRBZkoDfqTyON1OYIwYhAj4inTO/2jpqghvv+/KONCAuNk9L1era8LppX/3Kp5
VqgazHSs/l1VrGXldMTW9iIcmrQm3yvy15UGR/Pf7PoE0ZYfbrB+LPb8BdnVsaSbC+2hYIFK7Jnv
Dwl+7lfOxmY7NHOmFTn0QiaV0C01xrVVGU16hK7QGKgWqLPfHRlrbYgQ88Vt4KSGLDRizqXgNTpN
APVmP7En6EW928eoOzq2czXjMV/zK13s/RCyTYlasqt+P2Z36jn/Uit/psI77COjCODYg0CtKPRj
bVEU98Q4PTeDh3Mw64dqhHbI65tSLHvyf2yE3qQV8uBhF+Y7xHMlzh2QyIJXJFIACkd8qOCJ4tYh
9ZKOCz2VtBQ7g2UwaLYm8vdCwihwoX7ACMHzOHtwdu56Hszo8EU9TExfyqZoWYrlW/F10XDxHsbU
4GNkRRZ/Q7ncm47d1oCfQwEZRB33BjdHt9w1U3CtjreC/i3iuTmWMr1diMhYtFQI8kAKDa4FMd3f
RB31SQxwGtb5zqtJixJzOVIRy4n7UZUTb7c53sjyvozxkERsDTvjdAIGG2egFjEQ+QITlp5n6MxJ
t09UpamMn9lO0pXAJTm8IzK4iTK6g4WkoDU4KVOlbTnPU4Rfv04QsRBcsCb4pCKQbRW9mvzq0xWP
QF50dORrKth3pCAUHvAKcHQ3CO8PHJaUd76E3bnQvZ05FIJv+T+Za8rWRJHi0L0q/cyEFWxsehbO
nP3Bci79AP09F+JgzpOSmVBnnxUH0J3cgZmvtuH1lbuwwhhKhaKiq973et6drmlKDBf7wfH5F7NG
3QzoJO6+KmRnP+hb0/e+rNxLvDzCBy75P9Cma9KIaTRCk5nNV1hSneAmOzZSRCqh9+jtG+kBc73U
C1i6meRuXQpjHBfxImCC4eoxfJy9eC+0+SzfnwDa8BrJxZ4/aljiw5aY1cfgK71LIPFjsi632mWz
pgBj05iv6JZqHOEKrJmC1bM4KO/hTbpO2ZP7T4FNGPvr27mfudeB2KpMMX6vIllmeNw9pBHWVAC5
MS3TiV7EdQGrLeWD7oNzT6RjtRTMXTuDMSL4btQJuWH2zYhuuthIDKQbd4JAEDPrg8C8o10vvWA4
mxDY7uj0MCsN0S6nxTNKA26e/e9/SOuzNutb/Ah6nyRSYS6IbWFFAu6kPghmj8z99TlZJX4zAAie
gF1LP1l7+VboRNzB1Y4oJkCUGqgbIpVl8tDDLrBh19ylqjR0Ox8o1OehYNWU9s4f0EN71fk7RQt3
hsAiAj7duLZBkW3y2KDRh+b9XAX4BOTQ8Xc/G/g5ZZXAhnLcw4qZV6dcjnAX8BOrbZIcXO/HSLvx
lvx0J+UaB0TxtrzQpMX5DvktbdggGt6x4XG2hKWygPW4v/ZcLIsTL8EWhqGIEfc8sQ9wXaHKdRUA
QUymUy+cCfnr6DmW9jqa0NNuQaeYes4zgXsPNhiZvILVqpyESpFyoqaeC1gH0dRVZ+WoMKdMEW/c
LEiOS0h0VPdXfMbdKelNeSIRvBqUaevm5pouky4x8qpvWquRqG7CYvLLC8/JHmGFJcJEsHrNvzuK
4Av6+Cd0nk8znNFKLkLjHFkG74/UEi3AZ+azo3J//Kyw2HwCYBj1zHccH1+ipi0mriCvwy/Dboax
l5gn1iI+dlGOE+i7Yk5Qr93QkbxnQHuryqavyR+QzQ5kNSejakjiy2PFyiAqjCx49CYMmV7tgiJx
CoRbRRsFyneZNdwQEd7RnwOkV63ulPjggSuO1xayy/YwfmIIE5E3gQ4GuNE+m0SXCL20IUEs8l2q
yFgK7PI9hVlw/IOss8OCpIBqiuy/M5crvGxUlN+c6Bmq8dBDauafxDouuoYWbmu7IkqJqVCqwAUz
C7lzrPlK5g3w04Eg0gOZVMjFMVhGmnityN26x4/K5F/OheLdp4GGYUv8QkoDZBJ/oggZ/MO6huOU
yegmtRXj/GJ8475A8Bjb4od3LZ/Ygw6G9I1c9QHsvNwBcy+ZXRiH9GuljUW6tQhWIenJ8vFjHVh1
3QwnwKmtepUlCCWPYArWwce6XozeF4o1JxM0fdmdfJaRw/iVn8hXU8qOYmyMcRW393DOJbkmw/lR
tq8qq76kwIhBc7/RC8QUK0uEWlg68hejsRwTS31WX0B0De6iopJN6WvrwP5zLDMN1VWJGIfoZZgA
6kvAb/m9NLzGwJ3tgwiCRp1OMbgFYDk7jl+J7ZfEIBzgHNZg+0AxM5VZEwkFkInCzcC3Pvb9Cn4/
DUDLkVfxE4RMZ5wiLjPqAjUyUAwGYES8Szt6N+TaWfOKAKr6oKMS8ipcrgUBWCUg15+H9Pc+z9VC
CBRN8PMpyJN5Fm6EtUBmQegtXuHXJD6aVmVuJ1iOv9rPatm5XEmzTIrYijkXQZCaqncJbInSemAz
DLRW2jg4C51Z0CzuXTc4gkRz0bFxKG2DLNThsNqcJK7ysZJzUzE5x8HpZUSHjtpLMJ+6Ni6dUF0l
ObqRgyZTX8zJrv1ch9ETvenLS/aO5xYUei+sXMoVFS+4HNhBeq/cLZV4vlT6J89jxX4ws8klny0v
87j5eG6QIBTYlDX+/8Afg0lVnahNQsn4VEK5HwmxvLkPO6nAm9y+rtPc8A9J1M7nvgrAlwGd4kJ9
8kGMseTA5HEB4qo6DXcVfN6Oq8yeIFSnt8DT2xuOSNsdO6Sr3BfJz0nrpa3HUDdyVtNsCXjL7fmd
+R2O8ZTlMVTuW+PCx2D2Tk5r7nYeg/iiVhxV84iizE70O9L2Kb5QNqVG+GWuZ4qr/qiAyxvCb6FQ
AvfLWOA5r4ami+8oR9gRejmasA8kXk9uis6ZrQK+8nMQkvTKaearWIHEcmu0iT9/IVMNAUVHoHBb
iDuReHCszPS/JdjvW9e8eUXIEe++qeLb0V+4hC71qfNla1en33rvblt7YAhtcEIe5gMI9RT7NnYX
onzzo+IXgk/RLDFZ0ilfeco57weIz+mhkoROqRr6h4bwgCG0Bc5aOZN7qDCf3IFVh4Fs2nk8Gl8s
QR8Yr/ExFGpjeXd2S+UXHywLXzdjf9C6HtEQO8spcIIDMRgoTqX5tJ95j4hJH9O6OQTYEV0HyKLn
ODpkQfxYpYWiWUJ/ubPD/RfiBSFEyyJOocVaAmWo8fBCyMkdLZ+0g0tRfpuVz1G4lMGlJkYdwdIm
V3yIkpvAllWs6oc5/rmXlJt5KUNkLox574+vOmrYmEmA5BvghTtxelJb7fMrrBRvHgeQXqJifluo
7Hw1IcUy4F4gO7vOJ2wET+SBsme8ZkamO4s5CoyeS/rpx++YV511R7pt3397iqYKKnu3TMqRLul5
3N2SZ3XKSvM9+rWTwQG4r3FU5pB+CoGQmrb9hhF/hQ4NUzZin0NZvMdXWo38fiMUeb1VQ87ydeaB
j7nQ0FD0RNMNpL3sOYExyJSK37CPIzZhhS5d4/dZq5MX+0Cs1DKI4BnWNKbBsjbPTS6FCphhPzU3
u11yMW18nH86qmzX+MMUibj5ACjU/OptoyynHqPxoLGeiHqgszSYH1DUSSfe7QPlGQp8XFprM5vq
5Ohbsjf5ulzCwLD6VSOEQ8/mNVUkzWd1hHwGSDU4/dTQ2BbQUPXP/Fl6Rb0L7twNpgKl4FDVIWYr
wc8z9HfXr4PFRa8TXx0tVHLSLITjUL/h3grkdrtR41i2TNypTIJHGSW4SXtLEn26JjVXoS8unmyV
up6VX+V1wAF7SU4buQcMbOlkhc16OiSGYfGrqtKdmugZyMkVztidXSlbD5AV9C2zW2pHTXYqSXOL
yQIs8oRWcRrRKCGxQf7LUkY5p7Z/gZkbtIXki0BANFevdxM7hUwVQ/eubEZ9X3C8zXlFvfKWOb/k
HF73IwDAcN23up5yBsuVOnvIUcRWuaXfVwNC0hFCTIik+dlMdwjEeqtTmQyXVUN575R9+0pvTFs3
bQrFPp58B6qGvhGWwRtStEHIlB43HWGLpnQbCTFbO3CaN5W4YHlEMEz/MbpqNBD2UTQVYhskFXjd
2bBl0a0ZHSAze+sVlbuPHYkl9xqUSexSL4o/6Dl6g8JW0g/8dq+tsfgeeJmbsb+gt5wiVexfspdE
ststuOWNHqRNfvFxt2DxJiifUZTisvvKQxCmt6JVWzvKwowBm11mtbFl8VJupwnfDpJvI8KNz1+p
jxj8Knz+yiWstMD60xrh+2bHuZ3SyEf5XWYz9hiDsYolPCWb3urVndC956i1B/+WQF3+wFD8FBGQ
GUxvsUhjeBxWXYItdCfFUB8k7SkMMmGFQkE7elKmdjpcMhsqXB4PkKcXqmFVUodqAjeOj1BRrLOP
aH37b21CD5/RL8FPa1RqtZ+iayxrjsylaMHw//9U3ws5qHXZmPaE9/lU/oOcSgVDb0yO5feeFj/d
pPRqh6HigzaEWr4qu99EcUfXsrbDxVlMR0NnmItoVaDnWK/Ipwfa2Yv6n5Wc88ywn1QOWHlEg5K7
IZWouQx2TiNx5IZuWhzOBMM1KLLMGcoSA7JkRe09x99LVPEI/txcNu9McpAK5jBvNQr624RzDT+I
3tgyMQQgwq5/NeAwBXsWr0WqoQdwaHjnVlb882c1wDbcRlkP4MQnUmyC+2uxQk+Gv3zm4uf+hsPA
KTBfvenTdGHtdfAueiSKzriUPsGaCjJ1sMv1ooRqMSpShcdZLzE97w4Utmaouow8ir7HNSN97E0c
GknDHFX2t7BethRgdjYWFv3GI2W9ATF44KxUxMa4yvnG0dGPheqf7RXsT2cBGk7iag9KqANkp9it
sGPkVqKjrj97OguAFJ454/blzC/ppZee0EEMjVwgd62DH9wXqvcwufHFSgv8I9makZJY2ZAIPMOp
2nol0e4i85iy8B9xVy5JjKg7mWyf/JqI8GeUzd65y+/vehTdxXHjA6RAipwkpmseo5cVdXxYeTsZ
nS2HoTOO9fv9wsteoYS5zj2jCgLfSbtO2zd4zRYVbSWoDI+mMfTpdUuCqRI3+FhDcvtF6Lk/dZC/
ikfyKQVhqJE4XSqGOBZfDzPr2luGwH0MdUMJ4RPHTKv6NLRnGqWY5mfj75//sOSkeMUz8zXNwYMc
CvGxtPTuC3y6/fmuEZGACXpeStGSsFuCecu3Oew+OM3SL5cCZTl/eOiYM4x9AkV6LekesYK0uZ3C
HWt4ZUI+kZMxOKXuj92GB06Wh+vf9OfT78MIfr7TzfmRweqs1/A24ZVtkkcLRmztlRCYRnAWUbEs
MsZCCaUW7EUr9MSvXQBgubUfq41ttkDVg1sPKQsnBrXd0HR6vuQw1CSCW1gXObFADkQPANOSqRje
R9uQUoCymhh7nV3fsTugDYVVV3PqVEZig+XT4TO35zQJN7isGGzvdQKu8QlQGoBfh/B9Pkf0uH4M
xl+COt9N5nmb/Dw/AFWczwfOhSbuAD/tf0daEkDyKsrAGFkhbjcaELk90ZqVjb3s0LYiXNpTVYah
vztKu+Xwdnjp4Fg+L/MLG2oQVOGM1rPhMMcuzJiYb4IdRnMjAIgV6a8dtnqzzinQTJBBSMNCtBzE
dxvtqgXBAQVVK8000jb5C/mzNhVxSalSNYxwvCHIVUVMqJrZhZqs0r3xaa0bMJ9TlyEbZEuMyIHK
9vFzaZ0g0GGF4rgnmuMh2hfARXMn+eF6L8GDZYIr8/BBka2h19RcwT6e8Avf9HVr6LTL5VaCCEv+
x4Ch3tRyO/gZakrDI6o2UCTJss0bVjuhO8dCTaFXizO8YsMSrXztWXWf3cvQIZKiCx5xUJIRgpf4
BrJ3mSrO1R0PJFGCscp9Yf5QMjbsjWC0QN1gIRyDfYu/xbSNSU2zJ/O7ejIjCsI6NaK9okvqzLev
oMiZOjGH+yom3IQJ9Lay6Mi81Oha2ki8nYizuL45VjOuWnlTqmLEgMwKDKWaTUgXXAbbOPTrNmN9
1qNBR4DXzQ3dmCEe0wgCFgUmAP05e3Rvzu1CCVYJibgoj3rzURtLAQVCXUhUYaqtls/WtR9thb45
Zr9XHNbvfBuhamsX5yT4o5Jd9IBm82rj/v06j2FVS4PZVc5sXPNzIRu01Z6Lmy+cr5mfSDhfCRam
8FZ5o8zUJHq52bgLiNWkWUJO2uGAgCuUlHt+FnTD2ZTY/5+k0PuKphwVJsmUwO6pkDy7wQ75TWgI
/nfxUHf89p79xI3pjMRQwhhyGAMcK9hwBMngQ5TzSzKJEyFSCF6vfaIxnEamVGu0QOdXxu1HcsZv
nOjW7z5vq9XhjVWx+NWvRqcj5VKjfuK2wdQbfSSpxAEC65S/jKVe0j6+bkuSJZcpHBfTbvNQ/fxX
ghcXkEwYVKNLcLDuX5ZB9EPcZ0YDRyVbao0DgnPN6uyxRMACllUyo5jS07ibOUtUBzw8sdalJE4b
9f6Gh3TjlWPJEDupPAGeYSGtNjswngj27T0kHel3IXJU6oLZTkwSG/UoI3vb1wANske5AFE4xtN7
QkbIYnuBDCmWoLTF8/Tt4ik0uajf2MJ+wUeb1QyMam/mtChx1+t0bIahBTTdtdP57hJz2jLExl2s
iov64ZAEfWxp/FuAF8vDzp9pcYh67Xr9WtbOdu1kflOwxPpM9iAiHPhhgMAKfxGkJS1StrcnkckF
ViBEjAcWd75L2j2LD1V9a6UDcOJVaj7Zc3z1yUH9rQBITAKd0UYYdcWQfRgzDv9EPukYuWOdki1d
UU1akRZUp3C1izZABCl5QNn2Uv9pQVT796hVPbCOHVY1MFoWbEcsG2n/V4RQpRs3/kuD2evtgsmR
i6SgQFP8HdGRmzt9q+p5jBpgtw3E0ShIRP7vyFeF+44eRJm3eWsLkcm8SGkhnRmnHGJkLneAGpUz
jcW8KyjwGEoEKEx6nWFJAZMvU/DGIrO+fb+c/2Iz4kD0FG8yQYW5qO0aUMDR/xceLeLx8mG8RbUZ
EAI7FLP1k3AVuY4cZYfzaPvElMz8WXgIXDGSRN9PnEzjEeClE7lAbXF2PcVClp9FyYHl7MswInsD
RGd9RzNSv7fKT4zbkYSfQyZ45JTpFE63RslJhfQvXpyZtccMW0JbyN2duFUqe6HzinUJAmAG5RiH
0A+3I0m3d0vPVaQKYS3Mj85fo18+9J5BT+8oFodKIO+H8TrXVH0BKE+6Qxlk0MY5ObJBRPF6ggKz
bf/eho/1aEHWznj2eKOTnH8dQxZxtreYuxVxaVyJOcGkVyn1bzDpOiw3WC9oj1tFnBSpq97UNt6h
j8oVEmPH3jni6uXedd/FHSxeT1auI4L8Ao/ykq2uA87806/9NmNWewDnjiV/4/k6X7D9XpmjySgs
ffYfhEjVpj70ttDG7MDWPm5NVgmDpHCFIlmj8FrSKsYFlSTqhQQfNAGhEAPaNsS6qO6YIaNSk4zg
RsIauL/hlR1ioaKFZLYZlHZw62nK+5Bw41/bkAVE0PJg6hWMoar0KdSTFr21XCPdoBgUM57/Mgab
OeC2vlrYxfPWMmbpSO66A1cOvWfXwF6b5rxamS+LeK2C6rl13tfrpBq0EnNiulh+j+W0xC1iEaZ0
7SS2xB3HzTsjXlTRB3QqTTuEtL25SYdBZlinIh0w+3ugKWVwMOE+RXVYnysbRTkQ91HUNyNg+Sco
5nUgI2NLMOjD7h66JpH/S2CLgb64crUNqr6xlVFSm4n++wEuSFaMJ9bf+a4hJ5ud8f/rZb30eLVp
DmsV8RV1Wi9MgENrjABT3czBbPsDN6fJECCjpZjb+ym7RDIDIN8BsaS54KRXdQUUtXuWqvfgUvqN
q3kzRKXZslcxv7ilN+zhfkW5ouTg5lLy4/sHYZ2O/cJGamib+NzJ70tFTURMdubwvOQJrXE8IfKS
cRKpFz3nJGYbnlCWoGlwz0s8ll+XTPb5d44Ak2yhWQWiI1xdW7gXjPLwg5nOo3CJYBHu8DEc76q1
pMQgJpy54JAsKglNn6aFB7tOAmxxAbYpg6W6HE0H7FFXjPpQPCB/H54WrkG2SPiPHw1LdERT+d1t
Vp5cLtckC6Q9LSnFopad2BKwJ4O5BO4l3mTrzk+ko6KKGjNBnEc1scG9UiHn0j0YZL6/fqG1AAHT
LJuC2DW96pGVgQ4sOE+RpLucNoBiIrj6RVHiy1+vKpM0r3zZ8enKHtRVT34Gey9OE3xBHZicAntu
e1EoTjgyU4MQV3tpv9MR5ivdCcYUNt67iUxUgW84qEaAeokyywiG9mzz2Wwm/8jZe8aGaFI/G/fu
kBakdx6Rl9JUu0UfZRinuLd//IQMv6vJesGlbo7u+Z5oy/5kmi5gHEE9zaAW7y9xIWOSUh+wYoVd
IA/fGTgf0Ol49IcUVXf6ICKaYUK7xYPnQU2zr8VYTtRRLoWnXsx4Y8jxTcguKTCHhOV9glZk24U2
Tx2580X9rqVOPi40yEnl/ZKZ2UsjRmBjCxY1BLgPJUnihUpV+RAmEO8hAg+UOShNl2VN9iAfevu9
c3DmVc/cvxEHTVJ5mkay9vEFviA4h+NjWVmmi6oARPe4snieBinzlruKgM9ogD1VMz/nLf7ca+Ks
lcKBvwvK0OCgeerQwunrTncovWhKOmt2iEKN0L+miCdqec96Ro/Lwi2eABZGox/qmiBfFUgPXfpV
iDIl7xxeAhXDSjlfkuXrYcseqfAyLgKJoYAhMN/5IYqz0eXA3EH9elEAQ9KjNdSgU7ekYkYqpEb8
+6gH1lJpH5i19N/pcHRqo1hGrhShjm0vRT3jdpwNpLYmTsiIiFi7njYChx21JWRf9q8aJHk9lP/S
MmQRlj88vsTC5Fc7uK9/cmbwwz3rU9zCj4cYuoa52opcaRRdPQLpDlNqosgzm7+shoIb4dBV9Fj8
3/KW3BUHl+8QqfE+Nv3srhKNGXONXr7E/JCmChfEaVuL43s/EcS68KS9o7JVsJmnNK/nzCPb63qx
avCaq3tljhgOsEmM7fOfsRy93uPdFaXLF0B5DQK1yWHcDdG7oSrrliwmxAlp9lLIDhpw15EMcxxS
EzR+oT03ARr9C93fo1Spa/M5t/JP7aaOpCvorb1Lo7fz5JDuGStLhAnpVH20kW/9yyg9j6JhwwS/
CP+xlzJo2wi+TvospYhQy20W3t6utZsYqnzwtiVizSZxe5AqtoUCMS1m1b1CiFiH+qKJ9HjJQI5/
rAHhdeX12OGrU1752a33i1KVlXP0Euhe7RgsD4Ozp9RmlZSgOZKj7wvgo9pYCg3MmU2YBMYPtGYd
dF10rsP3RDqdJr+9FIP6vrm1xmxaX3bcsRNN3bz8XPY/uz/aB4DdnmZNXLJ7rcv5x8AOHAUqCY1b
11JIyGai+2wX6PasMS1OK4xuhgIlV4Yv6u4EHagvfxTrMrIvCulER9s/hA+S2Ap2WV0INphRbVip
06XXFWN83s3XEmP5DKyrgWLYWkGAYVECCGTm9nuQ4soJ2VdhtXR+omqtVyA5N31uLqAcXl3frxLi
qyRuLJYKcw1HUfWW7LQ8Blo3oppxZdRRXeBPkVQFYXXYg4J2+BCOwpeo/z3lp8UQlIHG7YlDmsyr
v1NVInX+GF3Y3OKmyNEBZ25ZIoThL3K92JUntPFdL10LxCob05h1ogieepgvLoOC/ASOdSlfxnXS
9+Z3xO7pAfnSnvOiu60692BjkTkGCTsk4PvQYNzQCNSD/HSlNnqhbf0nhrHHjNbcxLZdHYgYuTcM
zG3h98IY6PU1AEGUnhJ3SsXPKlHZjSzEDNfeZI2Mfs3Hg3YJcgIvxiHnvkO/TK/ZPOdo1TDaXyUC
9IDrCnKCrBQUMTu6iOEyEldBzM8OPxB+m4kMPCFRDnDdraEr+ZWkOIjES1QfJxkNp0wq3v7Ywwnw
FMFbdrv8PDizFbvlzFQBmdFZb7r73osCNTlcqKAW92CXRHmaOVeQ+NpetJoh83jdcxJUiT82iRcg
XQGwGIqG9c8E81F45yyxkdBm4CyOAc5lAqCcpnSsJ5PyiHyjYmTZ+fQHSSsp/YhEjcEfjSSdkeQT
z2+WuISLGqt0x1wsEZOiBFWxzrYvN131IGzX2E2Ji0M9lv0lQ4NQTEEuudfb5OE+59WFwSjnN4gq
iNE5GV77MA3+718xCe9L6zSbT8ku/efF4ZBN9edQjEmQGTvcQdtzfCsZHG/qqFxKFxRA/JSi2a6x
ECDZrsu6Hu+B6ZrFb0a19A+DjogRfrSOg+mf1TIMxD6/hwzW0fAnQup69Ca11owGmPXL9IPKqPZ5
3UYYoc5hOsKHJXUIq0KkBPii9h3Jm95603O1yqScQOSiTxCoE6kaoR186K5AoSuydXakg0bdcNVs
PsY57AsoJOvR8JNJVT8Gn3od1M/IwBuBcy+CDjyWbLZ9QZjSldL8iO6/3esoxzdE3vQmFPiDX2Zx
ialY1MCaqUwPd70p6XGgF3ldFZm3B2ldyD6sAXQwwb3/GaJl2vsHFFwyXaFLbHrXva5Brn6NgP0D
ngcTaeG8AnN0abC6SQ40SjMaLVUpoYK8RhaOaFa5a6HQyxCIdEymPudcZinPLznmqcdisAaDIVir
u+ko3BNCWSiL20r8a4Lyyngl1myylx9zvWHP89n7d/5aNLL3H20jTwTFaHmZfVGTQpAth2KftrYe
L61yESMTAyzS+9a3+ILpTuW3zUgOmm+kng2rbWyFLCkzx4TaJ29PHLDddV5NXHdnnV9zelx8fJtL
RMtI19e/m3IkFsPYiH4rwr22NXRXac3amueG97DmMN3qxviEq7L2DIaF3wxMhYEg3tp56j+pgRVk
NnbktDSlldd4Cptfyvv3HboNYPQ0v0LzkUVhYZ3OtNkISoqBGoYehTRN0mj7RoWiY6n80EM/JZ3d
qxRTNZiCGLWzpoys6g+3mOs9qG7+peujVR1B5If/vqSOs0gXZuU110DBAkMqULrAnjyku6ixadth
H9a0cf8V+MISpvEv/KcN9P7/cCXjuEf/KcmQWXZFjvS3HPRzKyvkFgHBdhyZvbf0mkE53Zeq1LQs
Au944mzHnRZf0kdQG20arndlrR2Ze211BQd9m+xlRn/HusmgPj1EO9x9dyWVCxQNQWcPfJZhVn80
ZfAaj8AtZOJzMIqjo24HhsD6nG+pxLdBv16ApU/VcReLqo/u9SA5RY7x8Np+0LZwDoS1QHOQWuO2
FQ0GUhMmrYCpv6CUB9lInIsOW/c4AvzEkma9zcAPfIXANdq5ZA15IY8cRXUnlm/s8k+41jQAFFh7
EfM5B05rIYGWmRpHs6kL/5z6miMgOwNPJvqDiLs8e2Enb6iO4jf/0UKHBi/gmvMgRPuzKSnXMei2
Tx1b7/4qMkbxbNHePUTwWPNETTWd1UzmvUFJb4bb2MGpDmpOeAcPtIOz9tWeh8lW+h6BADq2RO2a
0OIN6YPC1MUs+9E5yNkBJYAnclth6Y7wFSsXyq+P0bSFpptlj2f7ujcoypQWtrIgwclIDb7x2RWC
TJrRDfGA9Ydc0oUGvNbipv3qpE4dZuUvZ6tpRQwVpNQQkajGRBvD7BN0SiggssnXAVsJpZ9lW9kD
R+Ox17aZLo0wScGBpHC0C/DBYP7xqh8AIzbmkA8wLGQ508euTCCk2DZjfgmHGnX7m8QPgkJt18FA
PBEHFnjQrLNRNe2rwgOl5Q71ZLoN/RBprSbQCj6DDR4TQOmtFkV4DAb9wLGD24gtMRZFvP/AtCk9
SbQGPraNqAgkupkbJPQ335nAOCkaeRP/Vm+EPyVgPuRWcrUPb2/zM1Jj+UJWJMp6sia7sRsYzpM7
4Ztnr4KbxGjL6j+ye9FXBBctPE4SWIaBfwIukoh2/ao1rewP3FVkIc8lmHSpNgWG2puZqoXr0mR5
iD6FNPhMpTs+SevZhvAKe8vKb5GHr7sQnd42A/FUWIuRqqoEfRijtYuUhotypHS3xP4oEaHAYdJt
yDYGoXtFDQPAtrkj+mN+sHcco2xgsM5lpH1kGO27kYt9xXLpYHPBDsRRpkvAdOx8NSDGm8ktFN50
BK2/So7OQibkmZGK4A6Av5MBGShqvcUygMfAAq446wkFoVVPQeX48YhZSoQfcMJBs/y1RIXuNi75
00ZXGRJo+kpmd/b99VvlRrY56y2ZwKMvALG5KHp9I5eNr+Q1qB7NlLP/4r/O/yRizY1HNUQDQnb0
vX4nMdYvW3LJoCKvtMrQuzb21EAoeG+gFAAdAB0UefHyc8/vKvDy+gJ+wslF6a7S/vofS/DGxkZi
u31nPkpViEfb6pEygvIgE9nvdvXkLRzsHErfZkT5wNuut7qMuKpYOPr5i9slmJjhpv3aweYi5Ygz
rv+W4aDWWLPoIcR/0ngN7K0fWVfwSydDkKx2HdQY3LzzDdWCah53fbWZBPeUAYIOuORzxZImNeBf
h6+0gqsCIcNByCSncZquoX8/IwxzNkt861KLO6rArEWX6ABNRzeSbYMG+uHJL+w4wDhzS/Kk6KuA
qOP+u64f6sI0c+HyUvtKyez0TEPY4kOGDi3eQJvAUV2C1guuPtBIK7bhyu+XL/XAlwKz4vxNh07S
/nQCmQ/4beXRaLNCExDLdb+zkkup4YCfS+qA+Ux9TnsfsVarUCYyaq6Yp7IeVUdvqjwsCNPag+zV
q4sKDiOyG3o5Lj6ORqYV03kqodXknGHd1OD+cdAPcLhb3FCHvkHoQOYCb2p5OAmuJvFjvueZ/Jlz
XrAHU+dum+plvPxx7PhOZXZVKO8PNWJeqsYCNLC+FVj6IvANzv2HbIuUOFHnr5NR89chDFA1jTIe
ffSGe5zptVuLrksCweXcl67DD1qhjEM8WQJvRefvkMzAlyVWAuq4H59LusHg/bpIddczsnj4QEIy
IrrQzNVjt+BNlzUPRS7PwmWedzTgvDQGuZN0OaFUAIPzIg9RwSZBXdYyj3kaAkCXdAGhD5aao0cV
l6fesIVyHXOh7jiP9Lrh5AYI0Its0ECo3uLcu0+/ecXkjWTlrZ6bw9lHBQTtCbs1lkX5xpTA3mJs
pra9HBOw8DSJ/v/NpKWkfpgq1VP5VvYGZvyVJ/rYlp8ZrEkBB/u4wd4CVNRSlcYMxDTHOFayICa1
nSEQY/vRIcUM9PuC+e4eXTwaUe07eWwLbzowHPSdIvis4v+XYAOpSktoTu2KLGj481IWzUeMcl6U
YCJL39+GAul3U63RJInte8OwyEdjAxn7LZTVURKGObsU1yypXwPL2JDf8GBbCUejWzbhPsAhoXKO
riDwyKuC6ueN+7QQ1RY9UOJMsyuFkn6j7JLSlRrTOETRG6mIeo7y5xWonNJRZW8RCE/Z4SQB/ceI
/SP3trh8qU/YWk+JyQ87yNoUBWzEJ1+7kRqmBDMR5klsg+LP9Qt6gx+4qbE1EqVjYCLKcgOlwtt7
DiU3FPu6xO9i89Qq9odnakrxotq7V0GOz/qujhwY91M9rWVOloJ6drKGR3R6ASH0vgq92PtLEmiV
LKjveeaC1LMqhZvX4b18HIviVN2IWyL0xvJNrC+VoIW2ogxKVzVaIAPZ/k7i440M/WFckwwoVT1s
fV8zNqzkT+xinhsvEl7ci0njRhcmYRAFeI80lzzC+wAXzeQHjzWJ+tuM+10u8jpCi/RhtnG51Txx
qPbyaTAvgcG0uJVTjGg3iwjcMcep9RkAHp9mU7oGZqJz7KCgYNa4jCS1M3rxjJ+TujFHXprH1bIJ
oekfpURLFv8G6AZbwIkk394zy6GK/Kv69LkLqWrqQ75ws9MiVxH/75FTgUQZLGKGryEoleye9gaw
w2aqlPb5HJLC2n/12Ay9s16n5aYM8z/8Q0nEoRbSq/p1PmxmCGkPCYiNVqhjU+z8FQllTV+kfuW+
zWWoHVzlLsJSyZbK12VpzCTNZ/Nlt1G4GmkDbG+DrMJt3p/REBPn/cR2MR/BD6UdkdtS1/MITv6l
JkeU5l53nDV9Hv79tWFkpJiXDl/IS3K14iqqZeVkAaptdIoKGdgAWpjWgAEJhiMroxOAXnDo2jGs
jwt4EexUjJe97ZFVWsCvzKIMQIYGL9Qcj1JyWPn+oy8JOr6O+gpB8Kvjzg7uiRDqB8EgmmGg1WAg
w8jSrgMIBs5p5dg0G/pOU73+6o2pwfbdzPZojbIaNAgcr7i9mvxveLU8dyUgnvW6Y/rcABxSaQu1
/lQCwWSEL03G1SFuRjm4TccAGmSPRzdW+D22lUAs+5aYg/+CmbcQ+fiMiTwMOBNdlGNEubHBBR+y
Hpuzbl578m3N3bVX84OESYgd7NyOcMsL0KmLxWSSjIFNhuAuh9Va7xi7nprvS4syoMs463PI32W9
sQiByunrYTNNpctiWRapmsH6x9SYGceBLuvAvg1wqcrujj5mythKBNo5MBslWe/7U/8JW8ICOEGo
EWj2udbRiAIQ+QDeh4+LKo4ozqsegaxOQ270DN+Q+WIRApHgS+kVKTcxJnJipT6gVfs6PbeiTSwM
GO+GDqLOKk6nI1bbpRB7UrLjWpY+MyKf7bGCRrwuTX+Df63j+LAO3+Ouq806/jt3iyritLXsDyBZ
6FHSfbfKXe+gT005se5k8qV2lM0U8VrJTqlNTGQUlx1IlARXwGlxvKlQPqRKj2wDljCyoZnYxt/Q
Kt6H+7NklB+UpL/FtxBhxBgc0VytpWkqd1EllFIwEcWLihFY/Rx1gLPHTTbT3LqvleUXDQHRvUr8
1jWbPdUX0HGoPWmDGHKlc+smmDikdedOl7OxkV5EuS7w7iWhHyZus4eJz5F5AennlFJ/kQiIEcWs
ELlWD/NpXHBqctLT5V3WGopXD3PDrDTc3RLGqILnmaxLGV/EjmRgCc5nJZQsJvyQsCk45d5iwVo/
r1DJkzaun1WkjdJa6IT6BgcKIGlllhYRwtLPdtW+JdkqWZcE1WY/fmboqeaoUzubcDjjPnVfpXjz
HRfDhp/cXX0Tzx7MRBpWMONEj6Y7LdkeupkB6wYI+b0CynDL+FmkUjPk1SMfcGFfCl3L8SL+JImh
G5/od0t/zL5EOovoJMeKb2ZvAsFXB3uJhQv1CbeiRI1ch0SwJCPHpXS3zOVTz1//655x6c/37cU5
EmWZbEdYpeGc8yx/aKAsHT42VHSYinyR3xls6nPdZMfH/0m6JH134kfdeiQOljz0bo+E3pgD5b3b
o3SBd9E79bxBPaAWbNNCSoE/BlO1Pcf/CNxM1iuPkORuYQf6FDGUwoo1aVxJT93np499hr640MN5
7EbemcpR970Dlkroqvik42kFQ3KfvSL9lE2Dibh0AOC8zoNd9a90Fd+w6usb+0L6Mt89h/zQecAB
HniMbx3AOq4D5kApe4TsuMXAkfVkJEo27krnt13ZmEXfuWb/JNI05jNFTKxpmcIHitlOw8KqinrP
jXmIWgRiyqsMXKJKFJLuCJfwcR4FKoD+wBI7td1E2mTyrcT3ua0KzIOHDPTSJbbq26AAyjbehfWP
eOi6Dia1jeqgmhXxDAw1G3CHzOVj6+S//01hmXFRBbFonmPzHKemHVO+I/VQBMjsgC/famyO8ihS
M5aQVf/Fp4Xv3L8kvEoNbpFcwuePYwgjGyePduXUmR4EEpR4LqGM7VOaKgYeSqGDy/ikHzPtDLtK
jrWPoK+lM+yK4y4pJMo8A2G++FQ4OYCnuZ0UZIDSH5tauSnypz8uEH/1GMI9KtEWfvyULjDN2nVX
8bXqT4oqF0nKSHKEZWxI50h2gi/Ks3+MpSytDw0K6IgJg1YHeOgFj3dcLPfzqHg/m7/kjZSkJk1e
VvJVKpm94gpII3RMYoZSgJK3nd4C2cBFYdIiKYXLB3jnTBQCIT8jcWdkLE1E31x+Efd5azrcU7m7
aqHbq29Nv+keJmQOwVddLiMmU9NLSJvD3KRfWt6CdTLrqyc4HgK6tUiM5ZiLLYYhXdBrSbqEf2gP
CEqZRcw11xqw+fdEkXcMPoHeTJLRI7HFFN1By1QhbrpMEFNq1c1TBVeZ3tGFfhN2BPEcQcx+70IG
WOP0qgjotnqTQABH+0cxzDnxBXMZjQNfxGsbfBazl+SRxecki4PFWqlvVvf3t/f4d8gZSKr5MzZs
5IU/zT0ybjiN22qMZI8yhbdB2Yj2UzTcZ7x0qtrJlBIcaDIvmVEYBmzhRxSYfCnp7MzWZKfv4S9H
3g0DzewJO8zcrLEO3zdP3UCO8REKHrfbPqFypmx59E6q3WuzRosrmPWcGp1fSAnV0V0vjTdXV5bz
x5/ZTRU0B/sXuzpbbsTtueH2OsqZ1fUN3VFqf1ual5QT8uI5u9+fEzhY5oXw5G59TiwBpPDYE4Jx
YnMcbnJmssEFij8V8jGxh9BYPPq60pnx52MMtkpDFV3P5a0CxW79+qflAWUf+RIWjo1qE3bnYboo
0KYrHzZsW9YgrBOgTylEjDyASZjmVzBm8r+/zjfug4xdlDe+z6U89Gf+fQmJyg8nanYf+r4m85+1
RD/8XOexrXtH3BZ/GjiXFEKZwCtY2LSEwe0Cm+6ziXTMxwMsJK4d3DatzAEqfaf1ZCudp0IWAicR
Z5vhjgYe1Et2M+LUWqR6cvzjoa4GnPlmqMS0ueOESudnY6/XrnsvYYuN6338JBCKOOpOMYhZD6qY
qNgP7VwBCI40Cd9+Y7ZCNRU4yCpLKi4lDALPA7ynaRYmxjVuDImyR3EHcv8rLRGNYOhBEhiTDiqD
Q1eZSvIg2FtVsclWFwULeJCTrWEqeN3YSOnsPDSH00THGKCo58+5oUPJQr0zpo7gTp1548Be6V49
M9AyC0IMsLcnOKalQUElAph3GSf7A1KbZp3OKvyZ+mD6IkbFsCArgE9wT8I399VNQiWh+b4uwDaD
HcOHUhQ/+LFU3cVG+ar8BJce0ILQgsaDeAEnzpldkulkwnrndfDwhtryFevIhLnKh6BXDnWGQkJf
5Qcsb+Opd+YAtWiD40uRm1TWM1hrCs6HJAN4TcS5K+QZEZycOlHpnyJWycWU8kph/6ARMDV5do0P
V8ZjxOe8CK2GrpspulVROtiG6QVSeHVZESTvTMQLzExETS9DIH8FQoBiN+vAH3k9AnMptm4FAdxl
hhFFCrH8F6Dw0tt2C2nuQXj5+Pu0n5xSx2SE/5kobOp3h7Vx12/XJzHEt1MybZ2un1gzdNlUD5V5
mhfi4hUyfQVUgMijxz3W7xuoVzjljQx2+joC05JN3Jtd+RuCBUKI/tdxfE71etintWHwX9ldoQTD
dnKDxQKu1fkaCQjQslt/KkldUAWtR382RUPdq7IFsBC2a+vxf6gn/azpIcbFn05ZdPOrRwjIsHo6
2VO3nWKRiBAcR1TxQI7WKaBIX9Rkn5cbVBs/RwPy0qLe2yOnAFtIzku5ttbcIywCTnv8qL6DrOwc
4kZzW0WamSZPhGiZ/rqYVIbzEqR9cq0HobCfR3oM0tlxjZFsnrQ4IwaXSI+fiwVaTDQVg87+2bhe
0SHG97uAsxSexK9VixTVbsFakZjapApKkwsZOL3nF9ZtfpU0hxB6EDdv7u+ssMly8lCG7ignyc2G
qA/DJYhxLvJNYxTOzp0ryT9gZFAZxp64WhhE2D1T+MdWjuUb6B/1epvsL90Yb52QjQNTDu4sydm1
csMjF/qz82XTpi3G9ijQlcn/ibYNVYRGhojxGJGQQs4c7W4a6sa09mc3hzXo+fnL13npOoAEJ7J5
cN1BIGYRcNr44H+7AmsCbBqh7CWKH5fSgQG85BDT7QpS4z0gyTNyz3qvw9rg2LFm4sd5MNEB/fBL
r2cRnnlacExPccdjYqLqJOYL8vVD99pOnKQgiaMlIXPofoVmOHuqWySn5AZl7xfYEFdya1Vg0ndA
Z9FxjGzQsIK4lp8j8ljU5t6wpslf6RqVLxy7j9IITwOsMyWpPn9HVEsNIR7in0hLBhXBOPQz7u+o
s3KEv39Egn2O4C38+CZE/q2m5hyNlr2gWtyjw+8hU+BJurnlCj04DZndqdMzcKKpFyg38RwauGvB
xf7ztOdYhlGxuTY2/fZ/pK5iQs5xgsu/nT3L7XzJsMp/E+8Vpg5OrnOu9omCkezUEjHpWA9fx6F+
m+K9l2hChlNpgv6RU/D9/jp3rsWZn8jOKVhoyn3hivJoQdXug2xGhF+7h2lFq5IU6VXTFQpisdlf
PWzfBpOqK387igiv7salTtdg9Y5Bn1AUi6rFmMQN6UtljfdQhAfaDxRN2EqmY2uW4B7p6FdD+PhK
hhfMVvaIE3o6/Y+PSohIFRO/NlSu+ii3IjNa86WXnrHbkUCliMs53V5O4S2XhpFFEHydiEuWK7zV
EOcBlLPo1u6kpOGF0iJtop3cCq7K+gQjTJa5SsRMtmh0teWKLBSGvBwsl/kdM0WBtQm7scc+mp82
IvikDp329zBjoq9BK48PrK0Dc2vjFQZReI4f/b1NEik/yIURUoqvbxcfhg5EJ3YQ/r8V8e9P935s
UQffonyr2GqneEc7zNPEuWUaBjLY2iYeL13/6OpXFFbFgvCly69MZorGh1/wg6SlkmCr48kKI4U9
+nrZKO+QcKVE4czDkq0sk6bn7jVGrkZu+SnBU/MAT/khbXwHvipuRWMF7FVQnoTpZi91N6oHkgql
GEpTuELVr+ewGYVY3CjYM55q5J1fRNb63IzZcI01R2JGaVBFnod9i86hyGfohDpmVFieqZNIOW+Y
Ubwiss954i5gcjCTIcAAnqsJuKDiZFgWkQv32bgfChXDpOC/MSl/Was3ImTRCyds/W5q/Ae9pr1O
cGGx0r3JmPNqv/2/Vj3DTDv/f8ljgeOxuJBFdhvnXtLG0RWBa3ZzJG2PlCD9Ng8qpodJ44J7J61/
SNHERDHPiliGBD6HAFiHZCbjptAz1tzKQkbky2yLVOzm7uMqTfZeVI1Hw3Ldfl7FvfxzLp4CpPhJ
W6gz+RS0SatjN9BsI2v1LNcGUjiC73DHo8wC9D9jv3JKHLH6r4wQ63vQY7zfXK8SsK7LUHjAO6Y8
SPFcEjBTucWz6AaA4dTavl7MkHM+HbdsBpIZuWh+oZRSWGI2yJKRLp+AyVcZL09sUKgTMgnYekX8
QGL15R/AM/Zl746/0DJYuuqzeeHLoO94eJjxmxGLNmVkSfPeQanQLPosP50ed0+h5IZwl/96jXKO
5x3gCnDFfFmkQ5HVAAQtVYDKONWN2/Qy3AwHLo2uZ5/zG4++acn/zI/DQshS5zE0SpxwIchvGeVp
hH7C8CpniBgYjQN0oGUI9iv3jeicw4n4WN7QGiVwyEePUBLkiEmGMhpEBk9J3pvxzYXWzQ7bnhos
4o0rBo+Nu30i0g3LYi/AbAEIqZe9/lhuJBCUgTjGygVyR+8+G//sDm48diU3B2gZkckuu/IeXvUQ
3XA2lran/QPFxSb02L8qcQPNuZiUzc8zGEOb+1Rpvoxy2Zh0LL53IsHd4KCfXrgJMXF2OfQ9t3v+
dhyCaf8vqC4cLOStVM0Qni6Lzet6ukg1K+c3yNicloIPVWa5GtXVDD/tf+FwKid+F87vYQ3iTRkj
OA+sOMIf++FQ5oaf6P6sp8Y5HRelc1XZCJ8i84ZkC9p5HbTrNWhDZZCcF+qU1ZQif9NCATuNiiEf
ahnsDyhR29RD/8CmVYU0A5FH3QGVFGW+2rUnq7cSHJZUTH6osyIic+VOcpWI0zAFlmJpAoJB6sqw
szSYQ4aJJ+TVhBfW//ivTTqTQf4UebVTy7awaYVOKOn2ZcJey9/E3HdIjh2XBEJsVCYS71Ip1TES
3oxA+8Q7Lk67TK5fnuVofvpivZrnd6YkL2dZcFuzmlQmXEGrvF6ueCFMglxdNIFrwnh8Atbx01Nu
aYxldvqNdkyOJ7s55bsvs9agqR8bgQgW0CXqtquS1vvmwDc1bXYVvdu5Tmdu5hSQ/v/rIDFW23NQ
0WBqhg2IeN+zKSV0NaezTi2HCEq50bG+kTJ4HEy82iktKEgN6KQQFSDFgGWTgofVtxFUxTO55Z9E
80Nik0Qas9fZsYGJ4g3N/qAfx4aBRUa3nOwponQLddPD5Nl8hf55E2uGkg+ti3t0HbnUinJ23HEk
K6cpLnEqviKUTF7lpDFslc61RZZh4i0PmcZSZNUpZaeBsuwz4QlRZvDGF9O1Ar7TXNViOTu1E9r7
v2zqVXYrWHsg6oemUsbS1NscdogWSNiBdcvJ+VTKXW9kn9/IJ8j/rnjQQDlWCEIqR8RvMZp9J2vz
ADoUSpc0BDVAgwu8Zw3YpRdfmPeoBbMSwFeBUZkVctzovFz+nDQREijhUR1ar3q57P/C+bV4JiCz
iTAfA8zzeB9HF69f2/oxocnp/cxOEEzE2d5rmDtL+JJVgIrwFw/dpBTN3S2UpH/XVTQV8rfybcs1
YLJqI9jgj4RW9L43lAwvemkL0Sgn1R12mj/jSqeTC8C/Fa4s7W2RGAw01XNToMAZc+CF9e/+LX3I
fyKFik++VsfeIy0DwaXv0yU9/j+HtrxgdLRr668nvU13putTexqFOgnJHC9H/AfchuMNO3JpNg+J
U+tDGmJuvR552obvJk+q1ba9XopbbIhG+z4hCj61vNflY3WDdwOfE2ppCFF4S7gK0Db3wZg1lmtn
LXKhFkNkd7rnQ3pNq5CQqS4cJJZA4zT+cUfm5zcr/v18EXw7CnpI+X1/rE8FIBbzDlScn7HyRfsM
ctLG7c/IHO+uSxbEAB+CZljGvj1VEu4ZZNV9oaxicJfqA+zOb4a+1ft34cPIF18o0eYSmlzOjgad
jSUYzKU6YthoynhclzSg9CIHWGwkeaAddq/3So11qL1zm/m5hi5fEE7o0F1fQdmWuUxm9waWXJzp
NVkG//7iMp7LbzYJYOQP0DNB8JOdcCEcWuRRYajnreIOuvUcV9Ea9FCi4c3998cFZU0+ow18/rGm
cGGRgpapgDTWALHXKCbQRzhc3CEcv8zqv9Ut6se8VDZ2G2Zc8wPnPM12rO71AqwhUlPS9p64vJQt
H6LuCDoRT6G1OoiT1UeNhkXGGtpgsL01m0/n3WWxyXFzwOyVw/TfGkVlsjdN2nj77wp7mOj+2FDX
dqZPD0HQBPOazYh6rb0E6CRrNYpwRTn3kJtVNVaBgFJy2wqG8zqVDMvIQ1zEmAUPQiU5Z7lBHxdD
CKcu0rl+ArBHqsOGoVs1OCaeOBYuff0QY2rHU4uJ1aed+MjGfuCd62yDhxSiWCnemb1Rv87Kasf0
EUdcFEN8KE5jUpqdLUSTz8DK7fny6jBU7ruEmx9gjfsTQmajorfpg+Uz9gatslGqBGlOjH2rH99U
ynS6NlA7XKXtU1cwxRzRY0S27gGJ9pEMNxSAPEwWsMQXHtzWKo7VGa57Vi7LNh8JD4Pcue8No1Ug
lCyioIn3P5f5KvfwF304zjr4bWUfvqql7GkympCgzD7km6r3UcFP/mhMY+SXH8hwCJEr9LQ81utZ
enYqN8r0LWhNCLF7CMhfSyTiqyXUPQwle4Y53SO/6nU+fwrHx16ZR534R9aac1vBpDoULh2hNt5l
xwuL9Kd/qrX+ua5kR+p3jlf5t/OWRvSJYLf5F2tY87jOoXmfNkPSoDnqmTu4AZkAQv7d2RpfiVLO
wqnxnlkFYQmk/YwXxW2z3vi4/G6vIEX20+OSRAsepbIj7eH7/17tvF9+bC8XUcGDzc7kB+bRszwf
FNtHLF1qtk60C6tBRBg4hCltgAnAhljAjoCufPEHDKmmGAz0aZTRRmaQtSK+RCgB1YQX4t96EgJ7
0Hc37oz9IkZ8mDGol1eRxFo+3iniyKogWKr3SvZyWMZrB7/1TPstI8VGlZP7bA+mkRkuJHZEb1yX
aaIweqCoXbyxytj43G9MJe9cqvvdohy2QIOX1vUFFGBgL34No7aItKAxq0Tl7XUAi8J0ffH1ZCgu
nR1Hz1IezuyjJU1ePJertSajRUhvjZG8wBipdnx6KSTabNwzRvykIl/oR/OJO8/KKC/h2Z/wc9yn
dBjnv3K4reDsNgRfkON6/fiKZYftgK6btzkhs+gN76zgtNqYJrXb/zC11ar472RCgoGK89j5TsvP
lO3YtEFb7oScPyF3P5PPo+JdwuVRNI6Qb0hHnJUKriOu/q4qTybyJQUW8fX+sZVFs1I+6Xw0xPFy
e0lbhKaE05wDAykXYFQIdJR7iFVjzBC1HCupmCtUCGMXCoDb52uBsz5r5OBeYNf29ORc2SHGUsNQ
SOdLSK8aPtsbaZSZCUXit3R4gSOuNDrKZxfHyQEtd46uVeL1+JTLiV0+VElY6NV94gJPyEhohN1i
1v6b3eO7sR0sWEMxNk0ZUOv/TeD4FPMMnnl4p+Nsb/laSoCVvtqJYH9vgZaeuPM92Qo3q+T3uJan
QAkuRqn9A0LN04n66JZjpJCs8oKMCLD/D9NNvsC9TRfO7hrxbofs0k5mjzIB/ZlR9N0fUoVH25dL
uhxJlhMl4th8+qm4Xjj5bE+z9R/aN5l1pYrAuCdJELM9tqjgK3iHPnOGZ7f0TrnJxcQssZzES74I
JSdR6sgrQrmC99PznjtoIHecDBRDQmGG36bQDXNfz3Ft4gjGkZTtcYuQbdnuV9JyfQ+0JPT190jQ
aYT5qmByZkA5J11btqK3pFNMTMZ96QsRpOPOiVYvCl1FaVAuQ9WRgD9ai1tbdXwy7xfCp9k3MFJV
2UJvLfzr4lM87YE3GebBBYJKaygx3RoJ/eR2OVFMK+HLrRzZlruVWbBcLa96n2hZ6/25Y9AEc1oj
tAeA8yvGdgDF1BdIBZS+udeYZG4RrYE39VvX55v1UYrCkpyo8O3hSryT9kKP8yMSPnODAgFdEIH1
DiUYToWUjlIb/xCg7C7/yyksYZhjrZG57YnAu/6NYzNKEnJMDTS0dYCW/Svfd5lXnwX8p4+FPURK
UnaLk+3hSnjnKoxsyYb+5xhO5uidhqG3XFx6wSodDfSaYI4lsW9Ja6ED6A1v19AKjuaLPeXAq49d
yVwGiTCxCwFF7D7k2DkM0eyg653MnUCGbabQ00ZisT+/9gdKlDcK18Ge4bEKZSwl4I8GZnVEZHCU
4OA0eg7OeKU2hLdog1DbRiBqexwNgo2hxrHzZ3Us1LzfqiXT0SikrfEyhntbHRR/wKgyMZ5op8Z7
dUifba+qA09smXlFxlPKmG+65tD65YIyFHp1SzAIVMhab3wrLqYHVeXxCBBdyiCLYDsWWS69u/j+
mBm/xhcJjiiJMy0oGX3Owtc0FCpjsEW07l6+elfITzxX3iWZNdnqUZQm8NNeyMwV4GElRxV51HeH
NMGrV/KJKaVtD00wpeYAgYEEpJ+C945M5sK9I/2c1TaT1bUsEVoDwpvwk3T5eo4ICNQJAwfqIT8j
mUrS6uSeAyA42YWI4RIj6ZDLlDfB6mgWM76JXzt4sTq8TZkWDI26SChvMlB4ZF9alTKubSeRAF3z
KelNNfzOjt6/RNe+g1He0XapUdaa9TfQt20adwujUjvD9I8o9K6fTIRPvrZ3Q3zwz/0IkS5M8owO
i6ToBxt5DHzGJDe2wn3QMgZYpa3tEwoFC8RTnBgTKdDhVd+GUskj3f5w/0ekp93uZNoFkfCLc7Hi
zqEmlzTb2Ta44zVxZTQz7A/960LIznkwX4aQW6vnxURSzyi0tIjec9dnfK64wRBro9V3HzU5X83k
HPZW39dDjtgDNKdjmWsgj4cgoux/T6SKPX8oB4BmLYrYsNGBnk/0xehBFQQwPLgbOKHCtUoynY9U
Sl/dLe3EI0paZD/SXZ9OQ0+8a0MjnLmXeALmwDkMrWn6njohmbS6DAwK7WOH1RtBuOOKK8Pn+YrL
Y5XHa0A09gdVcpa5vP/YA16OYqJPGNRxr0hX+wx8w5dBKU1Jp9jvXiTpSXur3qUak6fCzezW+1sk
Y7hUtPrTjQbsiEZGhRQiVF9IUmlPF78yzb94jjJK4ha79YTRmYGpDCs/2QCnMRMMnpnnlXWzVoXP
rs9mbNV8UBmeEwFNesGSFXiNkN3XUbDU3cGkAVlYvd/Wj3H/0kndtLsk71fQlGGW9uT6Hc9YqEf9
l9Q/eZZV4GgFL1+/FHRWr/01D++h7+WxTHeooA5zZXXvHFvdvSUZL/OHkNZeN65Pyt7LD4cdJ3pl
fh6D/VNssSm+ES3Yqucwi0LDmPZQbbYptoQav5VAjScYBbNkuGwye006WCLvHib3ZwEtakOL1Vmg
w7HismgVJOWA1IaAvCKtTwyQ0WNaSEqka0X4jt0TqaEYNDgjxnwTvAYSccBl2Mscahn9WBubpCd5
cothx/ftmrTMreTbfnwmTlwqPCfSoWIvL4IowFVrgvMRK05OV0IpM7zDBj8IRoB7DqqxAmGkwuTI
+JOFKpKm7XUpde1cs75uTiFHdghJrT7JNPe1O6cpGx1oJJGgvFvbNECGdq8jOTY0LWOeyPal9BSE
jPha8sV/89io2z5bTOhxNMg4ATqt6KJ4GKzuWmZr2EhPjwEDzn2BstDggUI5Ebz/32CpcFxxnnaA
JYaz+BMCyxOkdJ0oyLgSVSF+wyTY9Dei060849jbnrHtpHZPSFUNGTakwEop+XrBpM5Qc7NI+0WG
Gh526i1pTSQ9Ysw/FtxKWB05dv4GhZ5N1x5A8mc/lKAir1KEPRrj7uYjRErKqaO+MiwHjfmQWUkH
HO0Bp6PM9RVYXtx6mL7e7Xdrqgx7AQNNOFDxbzYFeeiTKvVqoI5gs+Ri6QzT+hQdnwPGmWG3rAIH
8xk5aRq9wxHRn44zOiunXB9tftLAYUM8F2oiJxnnqUlsdY9B/EvrhRlpUBrOJGUwa3+fXkSeYhlm
v6itcl21Um0eLKG1FxjffbgnrVWtYLFjXZLYXnQT2U4d5K+C3VhSe06YQmGcrXqdroc1jlxen6JW
GUqX9k5kEQDVHB8bmWTVM3MY8k7frr45XVr4gHlShUhd5Q/mE42MTv3KBhjKzNpclzAMiEG0LwCM
If5sJHvUOIiDuEKXZHlee9mWxMB4JoxlHfEwCg7bI4Mq9lswqVBd5ha/DYHpzS49vVhKzxy5NJqQ
BgBmHHqUTiO8B/m1S2n1wNUVYJk9BAZHkmZSeUEkPdfrtesVz8ZKl/Npj54ei9kbHIzulABrGymM
B5gFu7568GgCRfGjn8KltIqvntWXgakS0sfFFo4d6SbC9fwCVz7mdsgi88x4RZgG33j9ylLSO7an
5BDRABA4wu/EXlYkpT/66hfRhyWQzKBCJB5mxL6e+LeqOBErPUCUgfX+KjBKv5QcClVK5/bj7FY1
D4a0BXxXEX9WFTmAXiYaOEYFrHvTp3i7JHHbzzhRr31Vq80VY5blDnU0/5EOne56ZaGl/cWtbRbE
4MlOw7ZztzynnLCVbWoB6k+VnW42XdUBt8uquvPJnqUo13OKep10hpl76HCbaTRHfwGoUlhXmuP7
wYcOd6uMBugQrsPErveuPsOlM6sJepwTyvFzwj4yA2G68qbckNjn0v58Xx6IotJo3rz5VUzzZakM
hx8O5BrpKfEbiwgX7cFcZCWSBYICyppXFa+ZCho9yNw56Evt7z4KYsPkig3YQdhajxH8ZPyJ1Udb
sx8xc5JE5S3lmt3dUOzp/GyAeuPHH4goqfThqBDbx/iYfZcx/XeWwgZXXE3Bk1UlujaeflJfg5zb
ta3erxo9FMFa87OnXTjSZTM9ZwCw/p//UL5Idmxwq2yOP8nQgOPZRUZyN2NOg9Lq45VX/7tUBrTC
zv4gXbKXh7RTguFc5T52YKf+XtvARrvnQ9AKmrgymdP6uTu0xzo/aOEjXclH2BPp39APqeWzffP7
VszU9wBVX8Yp3BBznKuR7QiQmlzdzGbkPku0NUEnC6cO6rQ3K7p/1sCFxnFCVKUQROlgQuKS0RuX
4prSHAwU9EEih7mnu+nbStjphMQdmROOsNL6rDlQD0ZmLAb/M+uF0RiniqyrS89yVzFUMW1MvSyk
SkCWDcH2KUeYsC4cPICIYb3mVSwr2cgKSP3hXrbonTN7m4kUOWPX29afqIKjWqzZE1wbFczdJhtb
5xOm7Tvr9fPPnnaQiRRTyL/llAKwppUA3f7TaN1T9JoOj+5x0C+50GpcLo2Dgqlb3ciSj30JyZN7
bRoGFelPsP2RFE/WX9sjpS3zdo3rcj2Gvdx3qaMQatMsGIL0wEo4Etix7Xf4dwFxp6jmrfiuGQa8
tYO5msyjZbnhcokez5NaUXugb5x9r39Pl+jxYXDqTErjpEwG2r8lhEACbcetXTJvUsycQ104H5eR
yxrn5tQghkesxuwsF1V3okPSzTf7FWKMU2kKDryccvcTX6M3YJMo4g3DIaOjBsyJuwx0MRTjfr5g
ggVCW5wtF2orEewQk77nMmH5qrTf7nMOVSRq2OXeEMu8sH8rn4ccYSeo2yD8XB5opJl7mZOLZ2oZ
NoqDHFINI2RB81W4WO2ym8BWRLbvkxpRZ7dVdMebrCWkwq1bizSjF56ZuXSBOaf9202ScDztUnUY
1SwW2JrrZoJvMjIV6iD0lmljHUdtH7n1Gr5IMviVzbqcbLYel/klRMt2XUIln1autHPa5+OK9AhY
D6CrW4AXKUdBd33HmwKlD688sjMDqDK5isZAiHE7B8ltoWPpTX887Jx/5LBgO2jUZVLXSmfpPQpr
+SdhJp8aOoVWQsGsdZlJT+Eirfs7YKmcKcf2Fsn2tFENRUL7wOrWHtKhOGDA2ctBdgcxuRiANhJi
TqtWjVTnzzP1VRfu0E/hIlJ3eBX6kqrka+vDPJEiTXo8FmRm+KxFHM3GPk2lUq3shpkOECIfVlXb
/sL1h3x+G07ZUNyeVSri1k1YmzBUJp1W8uph6Y2iFuZOAnkWei92QwFcfOVRHLSV9J3+gSKsSNKk
ieYggFnp9/V7HYhbOGK6uMlIk37c0c1QZQbJFqMsfL6P5l53Hp7Ae56G9lAjVZ1/HFnLq9IwDauY
6U4EPLWf6jNk+osj+bRENF0+9PcchnxfOMlYa7vcfi+6HdtsAh3m3Xs+BNvYJ4pj7hnmxyKtWl21
CqyyGpEZzb7GxrHTxuaB6dm5xvaNnywqjR9Juq0WvR1EYMGPUPPdkZ8GvS4S78RzJBDMqVo6V66R
u8qV8duprsA/O305oEpwv/f2tCWA+qf+ZGB0mSJu1YQ6oWtRXaXBGLo9vGk31Ali4vMaTEbBH7NL
yijYOwgTMvyhj0eQ5p6ruznJUMC0EpUbDVtVFBAaSFkftkC6MJNud0Qyks0glQ06+pMxqmlOe0U2
z+hSZUd2an5DMgDzGMVcNBiA5qE4Rp17Kx8vyy5MQbCGckqgsX45LstfzIuOE6WJDUN1icINNVyg
fObt1BhpdHtZn7fLXOIY6BtHLURs5mgqDg0kYArljjmOVFlJbLnrnPMgNJSWmfJBWk1LmXzDYUZg
QsgGoxiGaexcFooBpeaXR0hViEkwRrHcgCLdnOEtVE31FVyAroGvdmiY4JMlMa263+v13NfRb8U0
pvndCSBAHG2uv0Nn0+rO2M6sNYX/J58K3Ky0y8LZ7e/+G3kns/wjUrq+zL9k4Z++e4AaBzSyHV8U
UR71Li/h/5h5goC5j+/xN89ichF031obVtFTTjaZUjERBp6HdbkrCTeqDWIFoojxR6zR14PtcVv/
0tdOqxCDi7O53mgAnRjLZF6EoLfnFyREiGs8xiVih+o6hcFLLDyirqu4unkRYwOapZwqjeTCfxY0
owByuAFw9/Y2l8yow6ez1zaMHiV0P0Ful03HYGcZ54+r+CHbdcwjU01+l0z0o7GC1JBK8yJufmWZ
jm1fQi9IupSfkBqpIolMYG3UHqXsUVVXJijHDEOj0uzeZzZZHfZQhWhS69JhAPHtxyp5R0EKvK/9
7W0acLS5CNjs2bBDMhEikFsvl8HTk+qv+jU+Fd87MSk2IAjrHah80yQ9dOOUsDtiw8689a5r0Sll
Fyh+Uyx2CjDsqXVCz8R1XeTNX9z82Wx5xpRBRGCy8NTPydY97v9KIhBJ8bIiZfXOIUBdLF2wNdFi
60Nelx18Qu59Gvv3kBsOkZdwe2MlC6f9uuJU6g8Qw5DZ1ai8G96qDtCsiAaxAHpnbBn0AFUmd85V
K4OirUBp0hcs20xqDn5rTt7pp2DUQgH44xusnVj4Oixwrr1oAHl1EuVYNKiaaqkAKxyuZ0Kka5Be
2LlgRjytt9nXoV52oxXEUDX6CSAc7qwXebX4Jo+yBZKuZDXQnOpSnF5D9Q+guqISesqi9IZ4qD1I
gsJukk1Q1ekz588HojY+yBovN+uXWZh+8mFfenQNDn1beYZQ8vNo42U3bCKgNwBjqerLedAIw95O
VkopdaKuMiORX7/Z8YF6JL8BwMasHe0S05cpwfivk+DoY8G1q0jtEefOUw9AWHCsRIr+C1XCCIBk
HnMOETKsoBZFN1D69rKNfUiRlGfcXgByiTr8xZBLmcQ0lFN4bkbaYYhsoLqWx5d+QwKOZHC2BC20
xbI49yyO4alqam5zVc24eMf2fGVteMoeGwx86/7m8w7BqtdSR+CRH/D54QLP/Gm4BaTCgfXa4MSD
uZzoA23mweSbhKz8LHTHPmW42SMs5+3MANZeD99MjFFo92wOv0yGiUhABZfkqwEyyqePWgs/ftdF
VEIehzyIja6z/HrdGD7/8WMyshNRkXXrKvRjw35qBxg4TRMnKCAPVHuVGPoq1fG6IZGtfuddzz2m
4Bf2CyGzlTbF63XhV6JrDV8yNx7/nFtPUHy3brxsen6lqvg+laikHUCTdJO/ZqDbybzJtbBEizJw
H0zFAfFP/o0O7pYC7gyjFXkZDohnmdF0FzW+RdarTxNR/arFJfANOVJGSEGVI3JLvMypPCDbK3np
k5Y5ZbHjrXOUTqPlx9skKYNERI+n8pjfBpwwRO28PB+Z6nDq/NB8Mk+VfoMONvz281NtwUp6Tq3P
ITsfdEODiBGNXClWzeja9x2DtqEyuTtbTk3izPEj+ctfV8fDVGx2mB7B2tYqOSuDP6tQE91niAnp
SwEO1rhnqxmmDKnXq0H2V7n8w0DzHqO8t8UGI9N0OnODNd+D/gM17kYjE/3vOF+0tFeuEXVh+2vr
4pZf+BgTVal3SIVmOF10Ha3578GwAD6u8AavEHHlDjABxhRzXvlzyVay/h/+s7wXL0pjFUeHjFGB
PnlsvTxHUk5j17vz2NGV1Xx5cjlaPkUzyc5MSZaBvJ1MLzAEtsaMW+d63l/s7jwc3HCqCjqZ/9GW
6JbvHw9q+HRedtZwjHbuYeQKxJtkoEDLhbZJ4iXnRxlLCpPnke5PO7Bkk6tpiY6tRdGq4gXIE4eV
bV3GksVWnZTAPHVhsN9WSDxRf2lfUIOqll9NB7SRmQeqXLRi+i5R1OTNYd5tZ4WfGOQ8FIBEqNcO
i9sjbf2N1ocUdhdMUcOoS06DlQA/LnuF6LRc2FjE6T0BGMTrwt6o4FgIvwbdQaxPqauVQYhRrU6T
E4H6htAku0UX19g+ha6XG2Al0ZvSkYOd6ndXj0U33fY8RZgukIoP2GvyNgIee9jJL/IIb2Kg/7Sd
NKRBPzi6L5V0iazR476KGSk661Bjtl46TKpHWGXxczpS7vl9Rq2r5e7sT8TYqptEsQjLM4EGdFnn
Xm0H8tmkWPoMFPXKEjmPRcNBsHKnq7rH8fLZJsT4Jl6oxLiHwh6ymufhxtFBsQwmKWI+TfSNdCo7
0h4xcqP7UFLkAVAgou+jo4Feu1k34nhXs1hfpZxGnpcZUHCdwKCE159b4jPm/DXnw/LSjPWJG65b
nUJnb0e+u8Mg9ZT121ctt8gJPc4IkfxHq9iJkMSw8UJOQW1K6lpaKRAVHx1x7H5fKbRpEZcJdoyx
zuEfrfN6ePLSkf5HxpyMp1xi7BH0AGg2NUDl0PvUvVH5iOgV94UxGSYZQkqpbLVomwk83xuuSeBV
0tEweOrAK247S9ekkpdoUovGtTVbkZvDCR35BAPMoh98rpqTUCp+lpfD4HmTqsNFL/QJ/dzqi2n0
Dq2APpBfayUDckvnFRAMr+YWMW0r14iVWwToPdrqyf+YMhNVEnenYte6Q0/8MB+gnoLXWvGKHjzr
ERKtrCd3YySXz6w1xcU6NVQD2arU9xG8m88gL10sZoBMzsyQ/lgzIT+arzKb9Z3C9maFFtzcy7Rh
jQA55tknehAD9JH2ztUBRrMJelSAXyyPqvAF/uEk9H82/34f2GRp/RLb1igMnIl5/w2MS50BeZRk
TwJMNtnyi9nMtW2/p5mQgYKrM9O1Rj10lbG/c+Bh8hiYoJENyWE2Kep/n6GWG35f+vxVK+7Ion6q
a7KMU8WJpVrQx7O9ZH3kH6faMg3d4mHfxtk40vWjhCXRruzOYEbXeMoiAzLC2esaBpeorgYVgdn4
d7tQoLOm396Vi7qNUeZDG8VBk4gn5Hg/1LXWzgkinFwCC9dy2dqVF68o2rU0e9xihtydIqyV1BAA
o8J3NW59u6QvY+LKsA44gPmpBkkiDPNoTiwQ19f5xuiKgf9vfQeEMP8qQJv/jG7/myjQyNPH9u67
RYnQ4QJkHnVLlEWVyH8k7Svek+p1/MAhJI3ij4xIXQMzNgFMsn//X9j3moZnPV1udztJxibLign+
f5JE7kK5p/wv7Qq1UqpmBzGv9Vtz3fnH8YMXqiUiOAoUm50C1WIpO4RSgjOw1NayfQW8F1dBq6+H
9tbmam0jrfpPd/++oLQ4ajhdK0y1TlackZzwxQb6drk5m+ER1oqZU2pIH5Ct8Lt6U+sgeAfFD4HB
RLgjcyYH3j7dPTLfzMqJ/ADoqaeKy2YbjnFQkaunLrXiCKGXfDOevtoRc69+63ySWPkm8ALTIgbf
vwgJPDOniei/n7mfc4EK4vXLSFk1kK5JrzGwNV+ADu+KaiEz4I4oHhC3lW8FrqM+5L+04plnOj1B
s7gd2F8Kf6ddusmE2LBncysaUD3HA6aXVJtX5mUOZl98BWl3Wb3rpovNfL1X7zVrkvH2GIM38jtp
1o/2387SKaBauh/ePdYdZTRUv9zu31Dcd/bWPJCfJxHOU63NnGPA/A/h0sWGm0ltYbJrx0fWt0Sy
7igvUKu8WXBitk3+aOUgfXbnPep35vsQF+FdO9OgxsWuUAz4K8oSBRifSiB/p/j3ydKCRnJFtdrr
G5I8ih1OkQmGA8AajmCBTPH3b+gfggl/XOXj+li96vLQXzkG/nr5M0+Q2W8958HQ+0HAowyOy2TL
zqpFYTttGcbQAM6FP0UmfId20Hg9Pw+ndYdZW+7/yLIvdOvF0zn/ETlvECktiFHJwqiXPnLFbgqX
I51mehlKQetcmlbI5SL7mp0cVgEICtm3uBLvUNHStXtWEJ9dYKKaMZKq9p4bhFNIXpuZ22IzrJhb
GYX1fkdz/c5on5A0+7aYtJypg5Xp1DdN4lvcOz5gWPEQpY3k3DDbMJJvFVJRaykrhsLUQe5vk7Ia
HHb4Ee2LAzY9/+YkskIt08IoWu4VzrxUp3jGqoO0I+B2CXVzR4JiT6c4vSiakp7kQ6PQOlLwpn7q
mhnNVqabuy61u8dvAQqbNJIg3MadIZ0yG9heptXWY6TDczj+w++569i11chel8k+x0ES/Chx4iMZ
FMfD/WhRO67VruEBzlVt/U14B1P6U1yJBOVwJyeLZ0+sUT07vrRZTCZeGjv8KfthjS9O/pM0PPPD
x30tnAE7jvsH00l+BrQO5YS4A2eouxlsis8Uo0Q9a9FeqOvrcAO8Gx+JGR9S9hoAQBxaKoQR94Qj
EpFgLFGNYMU/o1duVFp9xrKGpCHUfbcjy9eH+jxJoHgOsrbQIw0iOEUPtN/RraHO2F8ZQff9twWK
+hCscTocyOEf9QlJcf+BJFi2zcIINNAszRDSi5olKsO46QIbmtTPb+0tPRD4C2Nf3JYv46GxcTSN
AvrQ/kIsKmDacTeUHULdfKDD/E9updCRxPdp+0GsTud3rlJ3KUdspt2e/3b0AnS62/4fITC0zywX
lT2MU9Vu+Ijkg6hwirl3MhDzSVssBkTj1qEcfaXClgHqb/MQ79KCXrMXEfu7usfdjaK25H9HDh1X
TqwHwSBjAvSX/Wz6CuiT/qa5spsZdINpAawd02I96BepNRB4CRpZHYNfBhTZEMOj1e8+5h0kdVzI
By1aDyvMQCZ66UOgJ7az1R5oEYcVJRIq1R5u12yABVEPQCtYiNHvmcuG5Urg2hJGKQW5u3dealsk
qLQHBH+1gSH32JVSUu8ZwwbxCiz5vRWpcUS82QZB1M0hPviltf+AegOuDMd2zYzRYOlqXDgrRjLN
yo3xdTf3b3CShPU8ASAI5F1EO/FolKZwzkWNyl8qLrrgNCHm8PqVtzdhnYnajqDLXiN89khiVw63
PTsPxBQc6XqOfdr6IItiD6jPGC1BQ+GEkzm/2eMdtJEOVuttiVLzyl6ZOl7zeFYgvLelOVjFNRQb
fFuekora/sl+K+wVPzL+goG8urrOSs8N0sNYlbUu9alU4G5Nk4F8DEkLFyy6xsGsCz2myHm+48oS
Q1OKetWkszXtdtYm12b6D6bk6evqnk+u1ElXiDxBK717GILGkHdZ8rafZlsTFRLkogKXpOUWe2Ri
qRhMpLXwd7T5DsjKLk+WrF2dX3ojF0fQpP9b5z7p6tY3KJMdEqXfphZIWjN3IOk0H5+jwYl8P3a4
s4P2HeBe5hN4Cpir9Yx/T7qi2SP+HDul4/ChPuW9uFAzw4gPeYkXWFXOqorBvwfEAfBlcg/01IFj
ldvNhtLHpuuO8UZXcLmHkQk7lxnS4V/p/riuNlhrehqAlMlXfKXgEtoW73kufHMc5K6+9VXkj1nV
CPLFC02bxF6zL6bUJmw0PYfTBmA12HH3DOStdHrxG3hHG2gVJQHsVZ2pc7eSXqyH9enrfM43Mk6h
tEsDvnGWs1pisO6DyPTcV0A21s8qazrxkKv63sYZCuuN0LjfmEIzZ8iWXH9pXFnyFw1bBgqaPSik
DKNJcUWX5yKTuJgZKUsTIoiERHgPZ7udgTboIlrSJhxGUi8Nl/CDAVgIW4637ZgkQiG02VDldTNT
j1NhUNcjMz0VhfQoSQetRuTyr+clAofE/VqNZrhctGdwU7fxAyCBC3VRrtyeFDZ+39Fj1eyY0/i2
j2tB6UUt4VoBdDogFdk0rIMB60icj4tU+svfLflRU3+ML06GBiIVyyINJlNMbUNe2ceeySwdZJSU
T3MOwI1gQLYWc43aeERTRnPQQEIPsTrQ8RNk0Ie9/kU3m3hFE75u2ZwwExbNmd20A2WlYw1NYNu7
CaNW+4ad6v8FZk55ocrC+HcezcOO2JOlvqnb7eluo0U36HtvhjStwD0jCdolxdws/aLlde0NOkr+
nKWWIjXiR/UJ3p+SRMxKubclZfCONCjngpJDeHKXRC0n1iCbmjav6C6QcLg4qW4X9P1nNLTe+W5/
fbVAGeAhp4/uxwHPb8DN4M03VdWaEgx+YYF+X2SRGcO80xydZJgoKcqJgMfhYZwKcmz+LmVVMXaT
gFC/ExXGJwEfbKqGtJb9rOjUm/yary/mmn7PkTqQ/ETtKeauphDZFfHiRDl9L1wczSkh2L+Z1fxX
xB6HmETBPxZBYHWwv84Bjsuf5xeZqlhVagtHjh7l1B8dWcMX+9IsN7ygFuO6CqNh57FYJ1RhLyIg
85mnAjxddO9sPBPoqTyn1NeBmtrisrPbDyqDBr41Q8MZhbU3Wxa2WGvzvo+PoEw/kuQVNkBC7Pi1
2uuZJ5MijC1Se9fcj61O7eNpSldgOmT1ViO5F6YJEucPervsvo0ywL69zpo0ctjFbDvT/e9Let8c
sBwsjKZV8lBoPDjbS3kzoCTk5zsaRmiHnfywXdVIB6tnhJIzYTQ4d3l+yedibfp87ucicf8DOv70
W/zCNRZAMhGApGnQDSOvdZQLxszxz+hr2riA/Lr13aSKvDFHNDHdCFVcvP7zTHdNR50gXgopTzXv
jGcLPJNZgG8EEnIArOb7ZopXdgwl7MXLnTu/1uRHvQyiCve+m7zY3s0gVV3tDifsO1e9v6QopZ2j
BH8g3cXAKS7z1Yt2OAZ9qcQNTIHYgAbjMytoPVtxxDJK5KRhnFiOgjNrwKrk3vcpM+oB5zJPTfKX
0TN2SmVOwNuXkGEft4n3A66QjWbxY9dXapecgE/HB3CYil4bBi+k7jaqRR3ehP/kJ4Al9ryehBXX
/QknOH7HzwbkwzHpskiR0VHz3zYIyk13QCIUcXFd1ooQJ+5fqC83s6pF27Cn6lLsO38nad+0ob7T
Q+fOOb6klUoLY2v6ZfIITu8zqtccRA1qhKK3OjZ0TGgjyQZVPq8kDLgJxDs99JWL6pjby/LwjxGi
Ebv8jrO+5dmfNGb3B1O7Yfrg7etX7UcZqmO2oKrA7ZVgDOefJBoCuTd790/5tloy3iWfIO1RMSlJ
gdYB2SrQMmQfKTrlabKdOAlJoCSF3nClp9Ky4cc8YIQfmBWSjWE3Ba3thDabD6IKhc7wJY285SOe
qOxvYIULIxvD9TdG6ZD3W6RF3GU1WqYWxCq7YscwyYsDUWje+1CIvwcmIDGSgfKxe/R4kl0PVWdB
jMt9V2l+DpsC2EqenUF3GrZqviG3ev/Acsr4nCO0+3BjJzpH+GxNEpIgfqcIixviAM+PG1P5OpNE
ctfXs/eT3Hps5yLtjVnHafgqZqnH3AKkSFJdvTE+Z5gAHO/y/U4AJ1/Wx9MaS+qfUKFaKLfspalB
iaTyVZ0qPXmmxXQwmWsg1voenkitdWJ46Nn5Pi3W35nY+0DULUmkL+hdShm99Km/K312aGSgmcU2
wCWa2bKEJBRMY1pWoclQBShuFw2VRZ5S3i7RZpQXJge29i9nlvTVRL9UMOQHttq5ThjLVZIpGvx1
1G9HaijJ5pxLmzKc3nLgjdWV3phXtfVNObVGqtBeJFJ1Sww/RVuEUXyFwjM4PVGvYPUrzQ7G4dHB
Rj8srIy3AFSFvfMNxtk6Pw1RPSkMEOy4NN0tL1/mnLPkyungqJDE1xIiI6XyDzU4/sGyQE5GQAmA
LzUyHrKSkfSPwtMJAjGej2Sbq6RzS/JFgksofI8/e06Jxli6YWi8ntp+3yEhSr2L6vaq8Ii/s0OW
Yf4dri0GaY92mzZm/uK+7SiQO/SU7nR6ZSVGWeH5mCYOdG0shwXTOAQqQz3PamApaMds2mDUmraw
W7xNgstog3gD1x9LrUYAgjYpuUmNCI6Ffj9g6HQzx500/zAJjYoA3Msq5QNe7ph6LIPgBxrMx9WT
KaNSsG/j4VkWvDULFW05G7y2gktCH3HM/lCkIswHVah/KD8zLDBRpxtM7j09Zp6WsoxAQD5kP3MJ
aZbG3vH3cWpgQXLbAKCoWfJMIvr8kC3KCcLlFDC48BIcfQRACTQgSsRN2GOLWA8HS52RJGe931Y8
vjuw0KKxOLvvEH/cjP5tp0gjSi6plGeelpSlrnXEIggOkZI8i5CE1io9BRosCRU2kREpqPI9fuBt
sCbnK3fwbwaqstl18YgNRxbZZygV6UCe8sooXeSCwanBd7gCc95TSjbPidEzCIMfuR0XnnUBzV7h
6Qen863UM0nWT3ODURiORKeKd7NdxQR2Vdm9hJYJEz+uCL5khD3qSBcp0C9Or4yf8wO3tTmn6d9n
HYyVEZc6PX3K/z/Udsy1EFeOqrR2o8q+P8hLE1+VzLgnGXWqfL+PlxYbNtI4+5gggs2UeaYkdKw5
xCCHzuqv18Qz/tfoZF/GO3yvHm8X3XED5OQ6/QztAFYoNx+MZgvJsKFyzfkB92cSEqjdIbqCO0cN
cCbbn5xeNgNuDIQe2hBu+ZA9XtPKK2vhLSoA8XLIaOS1pqXInQGt9a0slRsawJaKigY0BssqHneL
jUpUra410jcrVfIsj8fjsGiWfAxEWbAZlCI4CxZ9swPz8IO4C4DvetJCYN6qbgnnkYy8WxLtIcZK
v5myy+v22d8i244jnkZQfTg1hTr1rYGWtSx263ONS21Xq0yimnS7DCeuWcf3cR5KXBKns8RyoU5z
1jyFkuSRoPMhOTrVbraN3K7+JHnpkvtzMCiI//OeDjdCMQ4NRj8oECOb09Q+tYuQ1rMYlJj8SrXb
0RhuIY28TQvdF3MjrhWdG73juxuQKJ9ITsaBCso7T5i/f6uV7N21vEa0wwIv4sJ4IIz7QoGssG4A
ZuHI2/hqUixD9UO3ajRsZyB2FauxzAy5QwiOdCv4CQBKRiIVDiwjVAD3knEIOmCIKNsPgd9vGUYQ
tRQraSqUgja3zCXorgN5qzaDUzmpq1CxSax9wCXwYlXkjrL4MU/CwpeC/wAXvJiYq/mOLcMbYr2o
NM2TbHZSeTKpvilh7sL4HsXHmjL9PnBs1XdHskBtBs2cqMOjvY1ZXFoxAYM5iTjmNKFuHcf+8dgZ
FrqpyVF+6gs69MI8XYRairy8FtFx0VvZqNbqTKxu/z/b/xnLyjCXe4w/wQ9SoMc3OnbAfpR2X5x5
bNMCjMfD8pp6ZOmzM0MInAYc8EzTx5gt1E3D+W+t6RAM1lgHBVO6F0HVYj+PvfKOKbhDnG3U6JN5
GIQ0EpNMdWXMH+8ql8EjZFcIor9yQTkitL+6O+ncgOHQQQiusZIET63z1MqPBhuQHNGoYfPdwdDs
jDQCknfEqe9PdVZXqNYFXq3E72MUS+SGgWwozmjhxcrUQV/zj2rx/nFQO7vyz8DNGQrMn64DUk//
WB3PoIBBjrWois6x9QjckaNiD1KWSLKZn2lWFyBeN7AgXnimY7neUxamh4GFPXjIStWRfMsmmBqg
uevfLxg1AmVYHx8NuEMGZ8Uek72+igioaKLzD+9FKjt64uLCiVkfoI2R/RIGttE65N9s2EkyTSuT
G3m7FEaEt8ybqJU0IkOOfkVs8kVbq3VKET5YHDKjFQ0hYrIRKxK+qXA8OWof5CbBe4mjglEOVTjt
uiB5MpmJX+9qkucKQj7lo9MYr/NbCcMpQDw6iWwg5osyOoD111QR2u8QD/Kw5bJDQCd/RhYrccu9
630B3Yk2uOu8bPU9UmV7luCOaslabQuFt+5X9H7dntJtJOy7PhzOtTRlfvJ6EACUr2kS6k62TsGf
JbXFCJ4zfFg2sQQkAVtSf2A/1o1VQdO4UCqx2qWwrbt6Wh9QiB3wLAMeMf4voRIVOD29knDCvYtO
0avFthZ/sWhgQaCLXOQYGgGMnOSlfAl3RhNmyryXrpgC4RG1Bc9pN5UA8KICUQ2tfRHbqP3Co1aK
mlVAdz2v1KJP8xRCD/i2eAHkjTJT5QwCMxJPS2yk/Jh+/KvhHB87u/Scvh5yCNY6HjKrm6nTyVTK
pq3WjTARwsbzIrvp72A+J9ozlpmluOoT1zw4Ks+umaopVesGEQFw4F0TiPpFdlAekAPfwZgG72AX
nTCEkp61n9HCq74CYppL7SJFHj1c9DKm5+EDvMpcyAfUOtrzMum3DcGRdDSiHyQlMI607kITXlVx
aZKIbz6yuvRs+MH6T6Oa0dzoO+hCqcU0EBxkhSvFR01c1bCeC8Xqp1STN1RLB5/MFNb0UqiXbC/v
fXuYC/Dk3Kdj5hlh+UF1EZs4XU27Xjz+/24cu0q9t4PYmTyPCzcgzVX1QcqAk30gh5FokCTFn3Gv
mapzsfDjEcgyC8VCxfDdrp/0SVCwFgSJxav50K4e0Wlo/GDA7MpK5NJifuNqKYMuhk9LPm6gbC5K
Jz0xXnowmPD9nCC9Rroo7RUJJtNY2CPVcymAjg9Sb5AFCgUXaKZYS6cHAhI5lWZf+PKmocYwt0Wk
bbrARz2RoE+Ff1nqLOlTi0LahGUw3Kz3IrcldD5GN2sDedDRPQNeKNmNmt9McICuFn6++I6y/By1
h/JdxTwD4Z4katz7oPMSqJP81h4YqVHji9xb2z3ikELCUcFFLTXuTWmWx01lpEAONPtsecnbmYLM
RUisL4lvDc40Vy0r3T1oKLJq93svSxEJ1xEIXtIxn6wlmYrAvf1vylhHE7KMRzzW8clFjh8SzR6D
JzPfM3gvdQzdN7VnxW5PkT8Ra0TUCpJVIufdWfs4uEMVRUojEQCSDBTwXJruYsD2jX1ypYeES59H
Ih8/8WlVc58gBpJ2s2vM78DtJzWf9otEoaOTq5+xboixDk1KgW0bT9uSKazPnz7ou16j0L5Zsztu
h3Rbw9P4f3HYlvzeD5vBf2kR8br+bwU88bI+DdhF2tn4fMTAr9TYbEQoHEEdxBqjEzAYGuhRMNTn
uB8B9s8OefnYz0czqz+mQRqEbfIya5RsOIebpxI8HYDqu8OElbvQAtlQZPEhx6WcRItWI9GcF8Yg
oQjg4bCTE/QhVlZmODhrggNY5ZwjGy5ubKAyCsV/ghSfFKfQ3vTavBE1P/qR00HpjlSY9PYvZ0bY
H0uBHqEdkuC4nxscxVOQ0s8V7Y0UMhrjvs7kiBj8HLjdELl7V3XzvC0dDoOdkEVV+9KTsNIwbYft
+o76fDHHII42EZ2v3z+3Ci/fB/seC2wzWzsQs/UXwW26KMALPPpu0MRO8odNMe2ycDTmAN29cQ6I
xkId7gj80O2PcqeCzslnpQIo/SxZfT2xwdK2nVfFxvThJ8EIPl++jv7KMbeXHglml2MR2E4GJ1rR
lWU32JCAUfR3nnluqCoVmL863dCqUe1Y2E8ePsj+BbRIxFICAu2N0ELrtvdFP+YJAvTMZ52QVoCn
E+wlLHFqNefQWiCRpUFVDFEx7lrEoexBY5keqAybz2k31C4bwDPgYhg8INNAheZsAecqooVvrDmQ
+C+922wA7kNI5V09lQqtzOLBb+HPi6oD31m81s/B0uoirXqNmX/StcmjJIdYj5LC8O7vFq8bmtTE
ohkKKGrycGBHVN8nMkKuJkxZx/9ZpDJlVG8pFUTpIV9GTnmlwbghccZSec3xf4crTySaLrirqjyh
zQlYzCUXfMpNfO/9cpt4O2WWjKbYCsRKtjsvCI+9xgMGFJb/lAdrjICRhMdP2UA2mFacT+Ybc5Db
gFEDGCO5GIW+NVLxjHuDebG97BVpHJBkV+QtT2y+EtP9/KH/eUxDLOshti+I1Oe6sIH6Ur9Igqxg
qhU9Do9zIZwZM9xR7IdYzqhzZx6IwPuBxXNjPRKS89NXtL7OAbKx2dkPZ545HMVgeACRrk5PZx3m
LjOcshG9/IdQ8QwTwQqM+jD5hX0HJfLAwvkc3EMVEe+Xgu3upbiv5YdKkMh/1LBQXGS8UAbb53OL
7parWS/u2NxNVZkaLKYZ2K+Z1cSzV/cH6bH/qNhivVorXATxjHptB9/YKtRtqT7BVStjE6SzyGmr
gNTgWISUi2DB3geXSwLxPqJ8lowWFOaQN8zfHg8DB8toQkkdcWi5kjyHOEzPl7KPmfmqTOUF8V65
BtVdld2qhSWQiDwReFaa8CLe47zkz/1kX6Y8RTZXjbAUpliyZa2CZ0haj5gSkturPCXCnaygylNY
mvXaHql/RfAZgBZMkQK8EEMq36OReW1zUf0lND9LsZwONt9L7VFjZ+4Qw9i5mXGK/KilgoGioJa8
60TjqUR5YRrM5Qr6IIM1piTE91Wmf6qRTTf5vBeAz/lFYPqP80IYMDaS/b66mSrAr42miy9aM3AE
3mPYRWOP5rWR7eYkeqp+dX5h9uVek5jcjE1AYH0kzzqF6cbttX2tjMOFIzlQWyWVq+63kEfoVcgY
ZmuPG7cJwb8f3qNZp6EAScL2LmcTZw2sdHXKXYdKkxoKahMCIv5CTtB1PRqarzGFZDzHbKGob9Lv
Z3Ug/Ag1ejwXb6+NnUwPPRzo+mpO8gTXhTsOp3h9ZilyIHYb7MIF42ZMNx9Kh/LLMMHKRLaSlOrV
K/AApvO4H8JQnKCjq2TBChU+MX80JoCP75qYPPHSGYGtGGcEXGh9G8Ohvcfcfm6bPrprXZ3TOyOl
JW4aaZCmg0UP/wx9LnjHlC7WE9oLrfz/dhLIEF15S5sBJSnQ5Vs0DfWVFnCMgMesWYHeO0F/Udc8
tGgPy66SboVD3q3RrWJlvpJ768ToTEwdfKGNnGfVKlZYsrxfWlFwoimbro9GttcGVsXv0d3EM4MO
HC5WGzAhkzGEHdfmVHvIgHzOQMBU72ikyasbqQu01rORh8fiNQKGsfXitJXSH0+SOgxjREO41wvj
hnhmPPnOW1cX5durvwJzeRbk2uGESQvE68PtRhDKxse5QmZgaCELdb+jNbFCcxKf5QkNc4FkENts
cBmu0XEyALwTF+GVqgSZ0Cr5QfxLms8W4QpyINV62xSppxXdoiNltPk7qFNWTGOrBD8VoC9KHEFf
JB0xNNIFidlsnHXTXhqkGybah6EewaSFHOTMiEWoWclT1x7LrtlbIBqczdy2Rdpxj1/Gmw9oix6k
veJYpGQIQ+2FD/hPo5WWNRgWj2ZjkTzhQYnJuyGF2QMKfvq3gT2qEeLvC2jSygOumDeh647It1Lu
wDeiq9jueGBtAkjPljKFiWFQZWSW5sJOhglbJ1ix4jnGkRrG55hMEaYQyULn5oRrrdX2Ec5K+ZbT
MwS94hHTGhaHmQKSqp8BBBJ3L/k91WryuVlHK6HTX/7H6pxs43o7U8Qo2KmhyBeoH+acalGTWDQF
5P/Uf0gNsZ7WgD5jpY2bG45p1JAa32nv+Ysdjrjc1sFH89+FB5JThCcujk164oHpWorjMS1k8gDp
JaqJihLF1N/Zq90WcIMam+CC2RanCJU9vwVqw46NVXblmxJuBUgoi5LzxjtAusWfeCy++YcIEqag
0lAbqxmhqYLKkLvJU6Gp4fbEYYV0htp5Dc78SpOL/JeFhLS2t/TU/a4mnDOhkw2116CmYgZJpkrb
Sqp3pQ/dxMR6A+Gq5gW1n6ZyITJziKhSxI6lC2vgnJuLjC1hsdFzuP4SUkHSaUGzvEU9p4YnKHhh
clsFyK4/EJ9orn4UBHpgGLcQYFgnvMhkADUuWp7k8Ie8NWKYVkGMV9eDp9zjn5RITMEurz2YYmVP
A2dEQBui6iH1ojNzLO1i4AQixWGl9SLHqZHl8hXXtKpDEmtsJep5cOLo0ymKw1xwv8ms5UcwsqFn
gxpWde7j3Q0tt7JINz4DLnCcsBgs359fzQAQTeJoI3G/rpKkXgpjCZFp6sPXspek4LzhJeCt0M+M
posoGjJFcKKHM23cw76IP3rj7Yu26hoEHoZ5vFUSyeNM+8e1z532512zodFvqmiiDFblbbGv649M
81AVQWJbaWaZum8laccBgwO4ikdUWap4UArFZg8VvKDoF7Uo2tAmn/ElL5eDEZX2LxO1rJlH/hTM
A1VrK+VPE5D8lamwbGzijHCMuJHumf0vs6tqJ+JThDKyBgmzA4o4uxzt2USOGcIzMbVXFT1kcqth
VtH+LvLu7hETJTJj804kmGyeZpkh4XIrWp/vrhz0DHux5rBu82M+4eQmKex7azrh7eM0Kbk78H81
Y75oWv7VIFBZU7t7zrbBM/WNIbnS4jFsERGlYe+IzmRactyBZvyVp+t7o12PKjw5lty+c8Wbvhav
Tf0Vw4d2qHzoG13z0xsn7ayZrUlgKGJO+0neuxg62J7FTBDNJMZBoW2wLwND5X2hFu4Vpe8lrFQR
kWOlkcaHArBghkw/r7Abcy3yH4kplcA2ixWnEQQ8EYKxjN488au2CTTH7Ogxxp4OxqHuCnaAqbmp
Bbb3KDpJRgGuJnGuJQSIVe/ndGoiMwhYbQHnlDyTi70V7L9Rv4BabZPG+AnIMUwBcQSFubBQhiCp
fVWJTV6Hnyhd87KsffXs/OiAq1CInzbq45UGHSdZjkHR/0KdXQqclox37yBqJj9dM865B/UCjRgk
q3RtJ4+Mcw0MD2TsD07c9uU6dMCjXd7qmwzHchheSYBWvh19Fd2HXd643GrVBawcorrjXXi3pGWy
FKQEu7krGlD4oOl6zVbaOYZRY0QGQfg4rQQBK2SVphDLAGtue8SpabFyt+Vyp60g7GOEjblFVU29
F2p+giEphbWemRepoK97eO/CmP4j8rhusPt3lSepWFhBoOhUpXnhiP9a574f18OMQjwftst3a46O
JZIm4KHvRYBbHRp9sdNVtiwYVcWVtnHRvpQGADe1sDqi3a9S9sRK6IgJ5Gn5BghhMpdJyxtkkKZy
Qb6yH3a2C7J9TsZlnmZFvXybHYwaAVb/XktfmV0g+opV0KLE+JVExhSyeNKhcA7vkg/X/7dZVWfn
pG52gzUVNSgKIflQKpv43c5H3JRnq2BIrs8RbSVgVLAmb1ksE6btj45v3aKeJsanmlH3C6UHtu/l
Anp64CwdyXuZvpSzGnrlgv687uzsrHSa88r+nsxo6l5Z5YJRwWYv/P80Jo9BfHgYrY09QraqbOn9
NeVJJQEnubCdmRziFDi6SJ3TeFIgM/yTsmKuFs4Qvc/xlyXqOQz+AFwbRlVR/V7MiKyCx5vKGbfq
MXZbJqnlx1CqT/aIx3ikjwgMEU4I6NrFdQlL7qBQhg8leyOf09Rr/ewXVmsU6wROQsbjHNzv81NI
oeN4EJy0wZKCEGnonHDOh32M1bnHsIBXhL9JfO9zgL/eX4um7CRbCUiU2p64DvnrNVas8Rq9N+hl
qVjvQ8VjQyWWyyuXNLMHCX0+Ox6xDBBF8tPJs6MPt7v3fKTtYKuOYWdHFUchl51icOarxBJBilrx
Ct+5kBnuVG+sG1jWY5XadLe6+YANsOqxACwOf6B6I03Wm+KVFwDcqfHiLa4EKRYzvq5Qc/tL4r0j
l/a11UMOPyOsDpW6yP7E/sTq0UkZZWgBqd7RjUKFuYgslbVqTDwaB85P8rwRUPbl50qEk2MUyG1S
U5hdThslE0DuMuljHC+H1qXqLStT6RTxl4bPJwS8vRFamuFrwtcwGIpPu+oHtLb9bVHf3gc9wMQ5
3nnHo0i3bJoHv1qm0AbAd18TWSQUZG0F/Vi32L9fsYXbh5LRo/8oa4wGny/fFo0cA/2EP4rBfXxu
FEIkS8fm75IG4QSFxLKQ50oGikNmUOgKvJlK2gPENCK5n458+E/g8HtlAZPRX9CwIenD0CaXx++I
FKDsLQThexQmr7FWN672i0RfzIq8gckjFDehxYIjhDfOXiMAM5JxTUPGIWHvudyGkCdwjMRwHDkk
xvhrU+J60lb9VKXc1iX4BJFwEM0LmnfVYRXyBCeQWUadAFB2XveCfqYFv1IgCR8gy7HbGU58b2zu
J0dK/myxqi0PZetHedwHNHjqCoCCELTQ3gCVNE27R+3Y4uMAs6YXKf7tjHTMEUftJYqbyCtLrFEN
IaaZLAaTSgYnpdlAay28RXcI0iYwE+BFbJ9a0/tVcCJVYmaXvrCUU9cZzOf9s30bYleVQhH50Oyq
H92qmjxpgFiZCs1W33ra4rFDn5g36+fpdvanrmv2rCd2ROOG4PHsI9HqlGqmuuFLnt1U2vu4Kh6z
4qRUR2Iv+dYPXnxMkna3xnmlCvFB7UBNKCqVB8GGud/Dsmu/0lbbWKTxOmjSLEvTQe4UjkNRmDH4
nbrg2lvPpvlI0YTCfxtm4HHasTUWgI1Jzk2jPHIHIFkP99mrgAnpIaNQv2zKBQCDqM4g4/gqCDFG
z5L8UFjcT/NDjz684vQkQxDyRt+mWpmx38bkpbVitrDIOrA6/lIiQbmF5XE4J12gsYUeFVYamF4S
DHal+UkfusbYCajbQB/oUeb1L0STqsJfi81rRL1Y4zw41w51DQlJXbek+ODv6jHsKSlyGaCSpvHc
J9RtVMrwL5Zy+GGimzotmBsnQfasgFdFb2qsz08Z1czFG5YjFDUePxQ0l4SddvPVqNu2cdjnw3h+
PNDmn4cddzQ7vdUs/W0f/+7GT2FIwG0NYmcivxxF+F+WEvAS6hGPXMtdcAVMNibofhoFXiAGkRKA
ndOTmbL14RP4KiRgSdTgas/hNDQUGjC3MeDdOTOccTDJrTTIP2AffAnE8p5OxgWt80uK7CENN3KW
35mTDi+umO4PVW+qgVw82sn3W68vO55J4Nw/S++V7cd00+Ova6tqBsullwe51+SU3f8arEPyWYqS
XZNBFbFyetyinkf9JsCzAXreag3hQJJNTv0u8J5g42f/kjMwUWtiB9pn4UnZ72GyDTCbES+31bPu
vS3gOODTqieRdey2fdjSvv59NfnuuodyON6hCNtE4Pa8NRpmfDMUIfdU8eB/3p+1794heNDSMolx
yyrc+mlY49ccs7nVNQRr8R2lY9lL4u2Ffmkcr0HhnXeHIlwKbMEXXygdYjMF9m0hNjOqlwzNVPIv
wj398D6NpLBKqnuWU3rhMIn5LYTTO0Rj0r17mH2sT3IY92spbeMaUHiYIKdyslAUdHOQ71JKbWsj
iZOswKy6o957J7yZZ57nFsW86VQWTcxUCe94s+3VhusphPy1Yqu1cNhMdjArfGW3wCoN8JiFRxhl
80ASm0y3MoT2VjPYOoW2vDPkF5+Jiwb+K6+smLPwoETP3708FC26Egu9nrqngUCC0hRYhYIaPUD9
zNQ990jbvOxflaT9kpnZHEEvdPd6/OiHcDHNRVQOUHjXBb2rStBxPjANx2Gqon+Via3x24Ijf3EI
qvebgyCrXqVlV8ueg3jG2m69VbB/96R2TjyFzhSgLHjCfD13JOBM5azknRwpXZ+bB9ZmZw8zKFJc
oe/D0+qdG2gXwwEDbKDcDgNTjsl2mLgN1uPrhhvObmb6iRSgJXW/wSsii9Ohppg2/HQAcL+9fIti
qZjM8E/Gbp+YylnZeRY5iJBr+GQ39HZ1mIZf9LjFd5ABQaDSk3r3+3G+w7EqqlJysCaVrkhq6puk
Ut/9QCwfyS6TA9ksVoYxOjqm6CBCgoPTMFGOVr3B2DN9/D4kw4DXk29FrYNc3KJeWuDMeWtjPz7y
z92lR2tEYwRYmM/xned1T9mh7DXDBJmWRfgyJXq/EoJAYYBg52nnG9QvL13B1XDzMAFODyEdBLv8
Y4v0gX+PO8m2v0IMm5FCzqk1KwXl19Q8RFCqVi+I6pebVuUKUrirCFUNf5BnxhigdjzyAlosm3iQ
mLBbl36/wMnCOEgidEu+kQY266CXoru2lPnAoJR4yCeHKm/+j9RyZA6uiLACvCVeWDoi64yYoQi5
OSP+zrj/Gn/XrCZByd/fDmokL9wytdy06PsB3A+LaBb8xAppqwalQ/uxRmkg+yFVS6WOPRIA5Gce
I7Mw7of/2xROVEJAHwNhOjBmYkQH2B5UjstDvCop5mvf7R5t7+mWbddbnktwNWsM3l609nhkNqPW
Pf28twIw9H42GHolB5X6rBugyXLEhhLhHQamEfftPoxgUSyZxWvjokr95yxxkm+5esOwKQnIesj6
7ll9Dq8muGabFRbW00QJ/7IKAQsiRC4O6an56IAmifRabKRKM9tX54RxtsEa37Q/rK3gOM/iE+fZ
AGlUyHYFUsSC4jRLXru1MFKOE44RS+fJneWHUbrVQgVmMjNHnRMjmMFxk2VJ3Vg2qrRg+44C9lSk
c0GPd4qH+Fyke8Io9Y9RNRwkaY2PEKX3A3iUDtIea6YULHn2rb5lUPZVHoH6ychs1ZyNpnl+sSH8
d6+PkfIF1TmrEXN5v4G5S4dFos7Z9A2OinSB8W9QcZfEbOmOwePq7HNTIKXZ8/Tp8Yt9aULP/wtD
4cW+CKHTsJQ+to2/R2iGavGS0XQh1Wu+B/4dtvDxvH5oHWI21qf4YnANilB0MZkrtIv0C8DRAsVj
4FdDaIGHpARtkB4rS80ssC4sX5cgOHsbtXiJ8tsIJQpRMvIPQ/pyp5jAtuHWV7MlVFL/aEagqDaT
VYzhaMhF0cdhpi7wYpMxhzYiuNId6ZWPqXGvZTwTLSNHroBM3SFLjFEjv3jqqwpYl9VOT3R/BoLo
TTRtSmWsQCHHHNurwCIatzXPCOG8DWDKr7WKfzqBYDlJUZ0ZMYVFOexj2Sm6hOCAmY7exdWwIysT
464tH/oTS+o2i8XxJzCYlVCLPQCQO6tpJb13cEItyEUQ40PwaM6VBCJMmKw4rAfatsqgZVsaU7Hr
s9FNo/rOBoOG1TJ/FkZypiKreflFNKSInPUzFHN986MJ+Ky+zOLQcEoFt9wRGqedVUlTWtceoD+W
f1htcnw1wU8ieNjb8b3o8aAmYdEIMlXuVe3a5zjZZssR4ILWG4udHcl2J4LZHVv5lTasKTJc/Nta
+5PiNB7kI/25fLsrj/HyrbydiABlsVp11lVVTsBcKP2nojjblpMxRBqQbfvaPkqrJ8SlmcZBaxwe
/b6PA2TEyLfGWS1MWiED00lYCFwOIWcCKu5Fi8bIgUMQlfG9Pp100LVmB38xCsZ1y5gzSQXrkM4G
24AChLka4LRb7u1YdVvJLcu99ISC98b7WBTKcAHKTTK2wNrpQHOulQUJ6dzaOjMWDgZWLnA9jgAa
NOJCF1mztS7+LcYyJwzbLMkEXAlAyzsg+RgT9svR/XRp40geqbwt5d0XvfbuHD1PxQ6tSIZZjKpZ
TXhqeC76tMUGIyQ7YEiCxK1WBdBFV9dDz+Q7P/CrIAJ09xXnX5jcNQqMnpLE2QujljgkNEh8vfZ/
w7/1IbXCMCtP0NMb2WzwYO6dYE+QAqGFvMzjURtpl1a0TST2ds8xwuCYdhnk9CPw9eXAEzUeXy13
BjtQW2f1EylF857fX3ozqd5XC0F4dEjwCIMdqtp44/l9WdqIR/gC2cyH8osUbokHnOU/bMD0KUC5
RT/i7RCYEANQgnhGl3jG44e75SI9V7W3W0xet4zclc2eD1h9b8F8ZhM4sMLCcwbXJu95JlI+DvD9
Kunh5iU25ADUBwc8W3Cn3vWya7Irl7uUpVUsi0XlLA7u+5mxG2MoALB7l6mPRz4u15/OlCZFYvus
AGcau3JEX55K8DlilSxy3k3ZmTpa6BcAZJaR+gtGXJQk2ZVgBwj+9zWH64lOr3DYP2e/yvfyXmWg
1Y1uwrQKlWQLEEPlkBVon0sWRUAy9+lQyWha9K81jJnuT8ynAQfMxkezxuA4NNTcUCLq09eow0zZ
dMSSdSs1x4KCaWsPbXD9jiFnKSsCZDmE/GGkZrNjrqtTmBKDD6iZTigJheP8HV/mC/q2dfuPL6XQ
rnKap2qyoDo4JIBVwAUR9/Jf5ZB2fz7nu5PJxuzEVcEq+DBCazAjY3B3IeUvEdDphJmRB9lLt6lO
VdApjkQ4+TK4hkUod1KwTpSBezGEC+HK4BwQYtbR7lTf/S8bVbDSplIxHP8A+80r3NAt16dIqNiu
hj5YncxALpV2TjsZ0ILFNHDwOcsydnuhSN7d9TcRljqEoktj7OnNlXUgiEzateV615NSL3u7Qhq4
qeW2zGrV7SymdtfDF6gKn8/zBHNhEVxvZm/oZjOfN8IeuwScvbQWuVQmA3kor6C5ONYJGJ+7QAoG
gS6f6O/92QlSg1jJy+8e/AkBwrMK1T0nAXO4wfy1NZ5Mn+fNlZDiTqlPppNYQ5+wisJhIzThPSmG
53HrEjkGk/t0/Z7T9IguyvvhvAVFM449NptT3WkRYSzgIdDjD9JMHFa760A5brAfJQu4HErIwHZ8
uB99jqwPXgUfGCH82IdRsdiEu56dYfft3yohvnX8hLCKksov5CrJ1VMbWG4lBH4exRLG47a9nN5o
3Aa5UffJ1AIEideklZFYrZbZftgeG/rCmnJ0qthusOtjwCtA59Lb4Hh+vpQRiOX0XTOA4dxFzQfO
cYTu1TSmajEEeStUhctwH8P2zfFP1J6YSa6oxbE8mzdqkdKxHFs6BUJZ7LwTzKvWvOjFSHQi+pLV
uQMsGS92wfw9mKE48hAEtwZykM+qEe3xkJlU9X+Or3OIa0nrKJjkPJxKJdvTaYZ2JFA8HMfPC5Tj
IAcFbHHqvk2BIhjoRMcbSLjg0ovqdagxCD/5f61/KE91Yb0uc7ZmQ7jocfjtdNXg1JRAHlf0/cps
45UFnaFJbxqtOGQzJZ5xD2Nf5bQbHQK31Zj0GYWu7r1hkZfPV4Dt9UnbCxE8KebNAbV3h4wTod/E
w+rfCMpGd+ywAvcZAPkK/rvJH7Dy13zKVGFXAPlFlGHIRSN70mHlfEc92AQbCvK0EMKbNNOKfqdz
7or2Pb5vOBej8T/TQPB16pOConGNZbo2ECB99Gi73Nf95unm7jRkXjdN3GH2TAUAoPwg5pjcqrnM
qbHu+Yx78rWLQHGd2DwYcvZmZ4vvuOGPQZ9cOc57+Wp8r8ehNNxzKmF/14hN/3h6I66sa/zbkEbo
PTAvMwdwt15MWjmhv+JwaOq4QavouJvJc+Nw7yufpF7XzkYKPW0M4EBIszWkNH4ENnEO3z3Ol2+z
rL6hkGcYfqFiZo9kfOCBiWQ0mZOz0ipshgMt4Rfq1zrW9a7GaaAHnLy6fZKpZqRtyeuij7ElV5N6
JWu7eW68GcJ1HClp6p/bAQRb83KEsj9SQbjxokLsDPENfxL2WjhJ6WTroG/w/c0YDP0FgZiXRH00
u80eQJXvzpp0CtIzO2kHybf98xdYBNwizKYvOHhvGrNfKrTDtMekhj01y2EPtuWbR7ehtGFWNvAp
0/kAr/l2JUTo8LEnYejnmY4UX1qV+z948LQmzlBxa8PTXkJpteGMwAi7gEcsEgHoQld1M7apIDRS
/+YmS36EpycYaAUfbSdqoZjDJrKDKiicqiZvUzKG6e6Y+5EJUaEKF5rYlCHzP6olrO9n7HjMUA36
lI7W5WjUhkXCdSGdZ2By/JIaYcwjyoO2kRxGqyCceNM2shSYeOVgTSO7mYRmR0YkS6VxNUDjBVIC
y9yPI0LMNDe8irhl+o/09kOokjw4hW7Dx28zHYinr2q+XXtFYZTkSSnel353H0pN9qf1KqW86XAZ
JDVP5jZS6fezBinjbDQEUCZfZ4L2hn6t2jvOcm+coYoO0VFT1MeA7VXtrNFjq8bbBZVSk6WYdabW
AR0seg0eKy0SChmQ9bwomZrsuOQCGb3iKPxlGJMUuFLBDWYrsOCveGXDo9RAJtAoCD62OnaRVsm8
Upp2NSk75giC4nNNxruSpeJCAXIxGDX8AMOmmwrQTxFLILzJrjwLXrj2KpAqRm3cvfKifivfSnH8
bQTNwLhbibj9f/aAmA0Io91vG08eiCBDgctVfNZqQ7fsWGAvMSneflF9dF6rr2z7iF7SYFHbbFKG
KMzjsQ7FfhgeOWv0O4H1OdXF3gxDP/J+8r7Z7OhHgqxj4xnRbq6CXUmExDQsurbl+VuUliMWvlBn
skRy3cvPmcqhmbXsfWEMECZGwlxQiQJC7SBc4+7fcdiZNtdSkO1rXIhf/1iKTYMkzrUcW30ac029
SmdFLyluX+1y+i0LsHpRyZbHbDZPmYntqubM553zJcnPcuv8c5uPDj/lT9peWWorPf+YSNra/vqJ
iAX3NS7f6eTaWJaI2Q+Hp4ett4rtQF2Xvg1EDmg4yB5404Lt7VvpjH1ZxtVvLqzTnz3rKsqkflrg
5V+l3s1IeEX15rRrAFKknJfMtexl7GW6RoUIQCevCDgIgMtmqkWM6YcdbRTKWaYlSelzHP90AE4C
320ZYw/6KH0BG8fvaAmvl8EDoATkdfbjWZmnUblzFzpfBcO/ukidB3S63k7X/CfBl8GQOF1iFg4v
Cv+nLW0RPzGGQyvmkquvFs+lx+mC1rq6GmxnxffhKBnIvocIL9aGmY9728yKrPxolXRaIY70VcVf
d9vqC5mlZExZkVb1z43HvoKyEAGZYR4ZULYeKddK30GsyyDWPh5o9jCSCWlOQ0jrQIVXL+WuhewZ
npyVKyMi6Y188dC20JV0J0MVpwLoAnou7nNvPMxH05TE5kQcZmUufwJg34hfYREImK8v9ZBDGETC
S9NMZc3QlEaCLPv8oCrM0zBDN4Kur8VO/XLMNpUkQEABKGOCQG/xKz14Ca49A0ucILsCpCsYXLpV
X129shVWw9qgtUGYBtxzzq01V8bgvFTXVXSr3ypwUJAPor3FlKOj/UW7N5BF0H0kpypxhsClJK2u
OhO6KRl0Ve58LIhSHuyZ7uy16eOMZY061LMwTa8PAbekU1GDmhHMYm37qP/56BVI00YwWaxvWl3z
hmNgiKI/UmwFN0+b2aVyjzg96Sx1Q/RbDf02qQ0zVILyLrFIshO32UbgjvELB2+k3ViLnZ23gGWS
CxLc0wrB7bRl6UWGuMqKt6V4ZWSlAcjTFhH56BGhlVddqhVxJsFpOGn3V6XHELqJZ3cdktyYoopt
Al9/9ZZ/i0VUF4uELXb3hc96y711qMUKJlWoKLCdmvLgMJOCKCUv9NxY8wyHpoEjxfyVG9Hg9as8
yYMEXKbfAF3Qdcr5HVAvp0RNawdLrUXCnFfrqj9QUpQb4pkWitdXwfluPjQsHvgZ5RKtCUiAR5oB
yHdnRuq0OjWwSmQzvcLW5qt0PhJmUOoAPNMtEt7ka9iDzV1Ry5kHNzXZUPJ0/ODB8UcK/XuNgEdx
dvGsglSBcuI1dQmqJa1MQcE2nvAC7nE0LcZ34mLe5P747mX7JfZ0iVLJlUpBg9lVGBDCLJekgYlq
TgKCpLPwqh40dFwYPpD3OL8mJgeTKHXvensprQHmWAyByGA9TSsejtaj48bT8jhtD1DrfJdfz+BS
gEdddefCcTlnwp+/XoLkBja99v3HefKWGZ8zeFHTxEFmguaoVTX1MOxCPs23gT96bxE3l+CxPMLU
dGKHBrpKU0PqycLBLioljc4yQQE92KVJ4hsKSoAauMXxfPNY3fmeVK0F8OPKZxIQMbDCyQwmdJ3t
nPV/IY9R0idZLoEqIF9TxA7pK/9TEsEBIkzRXO4saswdBM2trO2w4Ch1sB1xPrsfCaqwZNngZOfq
rXdxw2tk/mHyynxBd/LHysAlZnLWkoI+BpfMchVCqA43EmuZQnkriYnh5GyRr5Af22ONYLoNJV20
i2zA9dMEqPCgCMR75TwRrcClaXCJdaNejgK7rfpO+o7R8VTuDNZzqr2g/JuvLTNjNDNEumUupvGG
ku957N0hCV/aLRNL27TXgHcOwDPHchiXfosAg9EsB/kEqAU5Jsodvb5JZ4IJlidAOODp//D4uFM6
4lJ4N3hEutMXMRV7UXTuTcX1e7FS3n7hBhpRhk2Na6SMArca6XdFso7zHodOKwiNHW2oUU1Crqxj
o3gT9gurwysC9N3yADsgPgWryQXqfKHnqov4+/yLedxOTfRpOruq+fBpQAyggj4oZ1MTo1tbZ41J
3QPwH2SzNzYG3gWstlAm2j+FZanDwjAvGqly8tbK288lFZkjY3qlM3ZzC1IY5Oor10ZHiRKRWMUH
wBGMAiaFMNq9H3tpCGrORprMmuNpxaTfdYSZyvnsytW1/i+be1XmVneui63VwP3JZxqCJsBcTRBC
yOgVfm0fJRjSpmSBkq+LtTsUuuQFa8rjPpYze5m5Ay58fdDDlfXUK6JN14LZ8D+AuOcDsp3Aq7CD
KkTqPxnbr/LCHduV99cvqDjkPG9fsMwRarhQsr7ntR1AEfiqkgvOLL1zhc9rLUWMBuKdyBwKKWGP
TjlZZx5ZE3N+XmbSnUjRVnhiqUFidbhQy5HvO/40IosdZ5zJ/1ta+Q6SlgXkc1AWI/Cb3G0/1m5c
Ni/LVTArbENv+u42VXI+jt/mbsIJZ/Uf+LtyU4MeNrFARi2EgoxEIAelw13j+le3h924ng1MTLjw
7q308fRS4MHb+X8slT8+x8jG4eYbWkOzvaUMuzL0anQmbBfoMckiCVoLLCvgL9aAfDQBWRSsomDc
+MGnUrqgJgINytG4CzmSr2/jQDUbS0oepkT4sljHDgbrn4Yino8MLaH8AUq0ai25682DMqHiVvGp
CK9KeKf55nMsKp9qNWDN4A+jGdrBVO4VFkjLBNlp+jwmMpuE0QfstBuKKMZ/KD+TClCpqrGmtEZU
rLM0AJSie4dT6O7Zd/yn3j4LdmC+2jpnX3M4ikfT78nNp8pQ6DzM5Iqf4kGTilWyEoWHmHnUd05l
BC83A3PgHPVXBYL2tGO+6oIyOcrL3VugU/eZYOs758YaEZ0vOHC1GhV6ckhlvRo1MNDnnmqH8FmC
+ZIE+grcH9SX26LRU2aaWWtEKuy4oYwYPit2gSO2f6LvBX4SvdOTEcZYO9jIsws/TJYYYiW7uzOk
Ln/R4a266jZ34/DQjuX5odSngomwcg93+U/Oluq6XehcDY7IPUTH21iDx81VkJR+Jy2R6X/G4UZP
v3BaX6dgF15YvxU+gNCKUVioYrAI8h9fE88FIaJIEhyhjSQCf5bDjvBlK9Y0Oa8ixy+idlVqvuGE
Qq1uwq9/uQF5rnSXQ3XXfelf6lPLq8xRPP4bN+0cN03bOrSpqOFbnl6jlac75QSf9xqc4R+d9Jo3
aRITIWvQFN5HtvDt+hej3A64EXickQPyryZVz8uc/o3dXFQ0wnIzxdVSTnnMUvkUBHl/YQAB+dR4
whHqcvyt7g1vrT9g5dFkUVZCdJ8Oeh6udxbKJL6AA7SuwAuWJu80ckF0QGqKlVmpCTQYM3YUJv/g
CFBV/JPgXenzxXerlDvHNsFnuFJjLrXTJLrUkNjQJ0XMgtLG1vMDJJwfgN5E/xJY4Qhdr8WGCOf7
T7cyJR9xxGbcTmYIA3eFktytuxmWs9XRTT8j1ewa4j2hd/pjQvxTVkhTf+6rxB/9OhZNvVKK3jkD
rwqW6qnSqeSqu9i6oKUXRyHqt9lR5OzgxQDVOOOHiEVQNa6DUztF2WT2O09Wjg3mM2xfDBYuT5U9
Wbn6+BaNe1n/vvcB8NlULpptsKXZHLPeLg9AYrpsHsX2osngnVomFVnTrguLlyRm2EWWLPIRA96J
1yEW3r0uibF+XYq7konNYNAXqnyG2je0+NHz58pJf49RKHxsqZtEgCzAlhsq1DxAQUe6uh8PwhQ0
gBnElcZlWvmQTVMCkD2XgnGczisagVwDy8VYB5YecSB4jtMlrsyfBzZ2E9YvXpLkSivtrcN+PjmV
A+Wz1/lIEUEOQf14E30sAfYo2qgkD5PevcxrSOP+hpegFZDsdW4sb+A3WV9fyWt3xjQYAx7brHBG
1rwYjSWb6AOHgUe1nUFGfIvkCLfIy20ELH+45MZcVhXAVb80jxzOheNzfa3N8ZhWwXF68etS0Wrj
FG/hrAWc1VmXYvma3kdyI/9t8PZO05TCdKtFO6R+RbwHaWKO6fO61oEzBPhUl+OMuGgeSswiJaGS
F8bBFN1ZXTX6zJyYb9gbBq/IX9Ib5VVd2o4zFa7Jq9Ejv1RJ9hUyiUwlkzVJB0/yORzOG4utFTeA
+I2yM3VIpOwFRI+OEa1IuFGh9o6h49Vy5WlLgUJO8QwO19CpUEC60mDpAdT7CLfP5uQgKcXwqZCE
9bsZ+HhS4Gss2Xo7+2hKCyPwVytH/hyVuiy348vMY08dIeirJrYalFyoV41JV8ogNViqTg/9iBeA
HlK7gQSrFUwbz+q9PKGos5NbaPk03+CW9HQyMruGcyhaoSLofaPaOtD4GD4i/KNAQYNUx1AA710o
OxUHHYCUwYrDjhoJR3EFnvmh5mychkAI8zWYyfRWnS4KmNPqlxvHouQlVE16uw839FUaCeMi1V3d
y89Sq3lx+Ii4dYLOEzvphXt9F0UOShdBFBBebOHAXSCKocw2JmEBLpsen3OFQtLG3sE88WHAMszk
b755sj9xi0mC1ySEh3xJxx8LDHXsOEsN3TSSWPKZk/PeTNe6x+n6gYd5Q/CzgI0J0IcFCg40WKPX
DQnUztcnU1mVwszv3XBJIQ1GNJwQViaCQYa2E6qLQRjdFT7mnVPXa1f0Xk3QS7PAAXm7ooArhqMI
kevjovm94IdtfXc6liPasGlx5+aWbJ8cWernGJbPao3Pe91rhGknTWa7d7X0rNdJMTzzj8pCUh97
N3NEPqfmH4RZYLRCl1G2MXvpChTuQnHaoSeCAPtDlDS7rMT6W8arA+phG19IXsQ4jgHXx4pcFS14
ARjUHTlCgeM19dfTD1WEzNkcFpOC34DJBiYvE25jVwVuVGXEe4e3+L7Z1yAZWEZ5zYytnXK13gha
CftTqjR/JFp/EBYk+NUV6o4Lq+uTLYn4hI7kgp8iIYpYK5mLKUowjNgPO8jQc+7r6L8/hm4D6Z48
97nm1AHGFFV3uJ9iDl77rekNwIRddlXMEM/OWPCS/os/2pU7MfeQ0hH4kBgqFiGNBfIMNy5sbPjx
SgrV3ju30eDoXMhe/Qtp4F4kc5iszocATjI3KDjs9KoEpSJEGSu8Bgse3egEmKtZm9wOPZCEfII4
dib5+U0rOSj/f3mQj3Qk6s1M/zE4Y7q5ZAbYlllB7GkjpkCBszoKI/YPmQFCbby7BjhgeCaYss6i
8NI+JG6Ii9YjrN8XzTheDSrfHQUlHfMDy2xEtSM1/Jk8jEWwHIh9PwTIrlk6EWNTVJ8L9Tz8BKaV
/0QIA75ZGvTEA/AK2eQFxFr7KR8uNPlf89H46Kt59skMqducFwbF++ZuHzCKbNgw55GOpSx9uTGG
MqZYbk/oyKDJmonGcPMrP40YlIp3BU5BYNi2aFT2X+UXv7Mw0NYPlAKsLDInsyDBjYCpTiALHquY
ruwu6Kv9vZKKlJPg9bwkIbur59PA4IU1kUWUCy36924R2MASlkgGpWzqOcjzZ35nuA4F1H5ayM99
Ny9D703C2alEF/erS1tOfcroQkIzZYVcmfW1yGlFo0kBKbg/ro8oYwArOCKchs71T5nujya3m6aF
B7M5PMaYv2HDplWERSfjuFLYjV468CgLbED3wp4tKBFZGvfwmqGgPJas2zKRZfjfWeePZ6vw7qv4
c8WPefTr7AheqGwppZzobofB+R+23ajPaxzL2lug0zStvPrshUFqAOMPc841UFqsf8vK+QPi7/W/
CqxhKhxqJb8a90UHLYOTdSfuIMM4exU7qPnXdjGCQzd1anECGk7Mcf+0Od5DaLR8qwamsf6u46oA
DKdBew6IbvRKQqbCyxAUi/dka04GJyINk40eLxs4vo8r5vD3Ol9FQheJlA5tdfublrDe7kAySCod
KFL2Y8b9BoxoukpkJ6JCjwVun+RdOw3UKWfmFdNIxuJOcpO22mSGXT/VFpP8LhEZJafP+iYAWAI+
cEWOV6JEA5H0pK+L128v5GkGq9qe6njg3p9dapCyPtHN61O8eKgAX1oYxNG2uEhqkRRNj80q1vEb
sApwvuHW37hPj9wkWnMZAmkGM70Dg/hMf7EdLYrohlZH9vy/FQSLs7JthNCX/I4kIdOa70RpQXqH
U2HZ4UhmneUDoCoiqBI5IRtvxCNhNnrBFbH5qxpmCJOHgtMkcPvTLeHdGDhU2g1zw0HjSD9OUX8Y
QNEKfoYR8xn6v7CoeFRkMCyGW1bTqE6BkL4bqtYhBlLI9YL6OpaZntxfrX99JkXSkq2R8qEwLdO2
8Npohlq+BVb1cEfuZCAd+F1CtRm6uxGUpH6VecrOrb9Bp3AJVs8yESbyiqwx6KeTL/3QnDkwSWGz
V6ukVPmZNj6y64l5zJc56rx1hk6SLUjJnefQE1b/48snnvCaStd70ZVmvlyjIiV0sTSBTAlmKX04
TGQd1iuupDzS79gQLXZTutgjKOvsNQtVR03lZ7YhKjHo2CwF4MqN5qauvXqTBYuQrtluM3hjhjn8
TA0eQqLHuf6T8YZt0oz6cyQSpNTJaaa1CnmJ3pzaeWaDsjuD9Ys3riB+QbTlRHK/IOn/8XrmVsGj
tz3TwYn+K0Pwo0nZSDo2lJ0EoIMMTSsLJLa/g5eXb6cTLlnhV6gFFRX4Arw3ljhW2gZ1K+bck2f8
VcOKEqwJtYaJuHGAcZQHCJ8fUAckKnrodeHe/AiR+4838A7WBbgZLQQt30rLIQ0GEkqjMIzLUy/z
62gSEwwjHNiZNbs4cHtyR5XSCOFVltvib0DkW/yhFAOcSceEV7dxwPLZahc7E1YPZVUrlzjeZpGB
2/crK+G8c0idcc2b3aB/dBWdPk6ripeMTcUnHwDkigs3Cprd+apg6mKJ2yLIMoVFLW6rPjWIFf8r
CsqkAl3wZlzsy7AN+xWv2rR9B/7IXk47EPL8umQb/H2YznR3WQCaR7FT2bjhaKU4XZV3SZe+JSF+
9D+pBLINEQw4u+veECu4e5LRKdBAz/Tm1mEBls904bhAxEJI3v74VEcGAtFG2DgErjsJSLcc4Asi
pf3+tbT5yaGn9TV6/Q1Jwe638r7dwUii7XFGmf1vpMvmAj7MZTse+y/MKUYzPCxsaiiivdkMfocR
AZJA1IlaCdXiU3N/6b8VNLsELlKmMtzikWd+In18ttSQQBhT74MekFMOmpnGX2zl5i50JLllDj4P
HAPtXixINnmGOrlwke6K+feNKUyACAcBcXie/x+DK1xh6Q2MBAtPiS0i9LSn3CNGLwyLVx27O7F0
llZN2RHkV2nmcxFmsVvsIBYuUnVwj4dgln2wU+av3+l1N0Ft4ylVlZPM9sy2huOH6CUJic2oxHpF
yPechTjsVo/xfP3/Z3U7xYZyf2b7gdjNutcAuUbTUXNt8/6LcpISYYxp8P065kn7AhZUWneA6OR4
5OIj68/N2MEC95EQ16sKRp1+R6c0j/CEH0dcAF6KmmZcnKFk5FYvX+lJaL9FwFine4W6BA8D6zr/
SqxFdtS5gZmqQNBAgmAIccaw4Cy9SHSGjQYKobCwi+Mxh+uZk3A0mRIhAqYA9g0zJwhHzcy48mTC
YPRQNiDFhmjyMoEJjGZBWHrncQ+0EFIna213QUIhRgbDngOhs9JnZkcFsba+2cRwdu+wwvV9I7pd
Eu8gzqlUm3oJMVTeyySnWvSaEk8KlZdlgCxGrmfTIxEFyALom6jQxTS9PuM7WDQZ4yFDUUo/Ojr0
0zrawfm2w0sL5lc5+g9BcsYyIuiMtimLsycqxWsLFfspmUhqGF3a7GPtEh0lpL+6p50nr7HrSVeg
+hoGkcCIq5rLde4ngkGUfCosY/neEQ8DXd9eu10BVUvxy0hv52S54hk0CEfe9E3m8Rj8zMBzTSku
xzTYZYksPHaJPsvdQ1n49q3zTWERgEQGpnJxyQwZbdSxIN2uMYRuGmek0ECkMTeJlA15qmG9FoNk
5mOPRi8IHiIbTgpJJs2vMp2Y564TAI4WPX3llw4aWIrzXuG9NjLY6zQx4eTg+iRKSqrL1C20VEYe
OtQb0sB6KACmJVk4TJ+cpOj3cmDZuWukUilcvOJSZNngg9+vnyNFdJ0+4vYA5d3UbN4Q3LFbX30R
hfDFhnxsh+QKy7fUaqmRImtJSjWWO576WaXfsa2SdPRMVBuV73HAS+UmVbxYj+Euh3deEU6e+M0K
5UJTDzx0oHsYr/ymcOewvx7Sz37qcRMO7RoYsQoBsQavCD8hJXTlO+N88RWaD5LUCS40zZWE61tx
iF0qef8LIzXPRm+iRizI3ZGBpsjVlVN68YDhApqWvAqcij8PuAuWKy65geIIzKNlDBwScnMAB0cB
XMSyBTR9Fn9XYtgokuStYxKU/RoRwu8zvH3yazlTzpetTS32xrxUUjnIFewmnFEvo3PpWARUJJE3
57AT6eJwXgjNRkU3Ayy+twF3N7XfjW+tKhdY3MQkJujEeayAhgMXqPRHQK4EGl66KrgVr17UOVbA
30pG3pPvEc/M7iIKzirpBTieYNdfHJ6E0yYbTpLvpf3kEoS59hRqn0Wo8wlsxzVEPpyDLr9NKLN+
E54ygiyXEUSOcUptdkiIN/c9IHJLl17eSIybEpMJ3gIibcn9bnKBAzbn6gxFVo7EwoKTOAXI7NRo
hFSdIflR4FWrZ/eS7q6CVIPrr/R+2/pN2UjVP2vdyIeATV0GwGM0Tc9jlEdIkUtZOAi+US/0lZUF
JsfDokC6EnVclyNdEUa+iYaac9ikcHmoEEsA5AbrewVreJu2/a9aUXLBZLYdxf+GQ+3kwuv/l+A1
jgR5u23hne+jmqJN3MUFtTdd5F2oTEEhUqfq/SMgvuwRIMACydrX/sBJ/zFDWuU+NIoUO5gSvOw5
A17Pq1dMPAYKAwD82cot5Apu9UwqqGY3Xh/mtlsTaLmy0PEUOgRtSn2F55JqaCzOgKG1gndXr87y
fADpxh8A4PPcz1DIsS/wVcZvKP0//gLS/humUnNSg9CtgQpzh36B2+oSaGOPOSU7uyKP39odZTGF
40mQLrw0621whljCfEsqm8ozq2RX3VhNHQh8xKiYa30JxdheFJohM5g6x2WenQm6qroIDG/vkb1/
o6vbhpWjLhZMDnfYpJJ2nJ4za8s9U5CgzpCYqGWzTVOxFqP8t9bhUeqdK6rG6/sQE0ek7daDoVqe
QwGj2iuDQGqBHcZ2qucgIWEiMi0z6v0mxm3ITCQmlNcRUq7sBo8S7hs04JXQHBnNjXCjt7ZHXRiN
5iVflyUXxANARXJMMyUB9J21NA0oNJkKy+x09lTtrTbTDszzCzYJobHBGQl/uAptXHpmv/8cSvNH
fYYOY3/XHJkiIkfTdN0Li4WDMVX/lfUP66hywlj4ZGrOgPTUH7CgN8gpyUvDbx93DexUw1OuL7Jz
abKv/f2BXv4rHW+yt+vOKGcS9FnsCvyusdi3r3U5PP/Q+tMu6HKhrAZ/uUDRxDqXhuM+ke0GddOt
WIqnyrfwjR55VG4gtzoHwUhwzdhbrNzjs2aH2y2/28DPHQoersot2QNZRbMuPFqeUkbflSuMIVXe
K2LVP6IGoWnqNQzJxa3Q6q7nQ5N92sh9Sr4D2ao6RVEhtQFjJw6/A4tOVyRvJooEPxN4M36BUcX1
HmWG0mKwo2quPZmYrkLJvHN1nP4FYDsmz7NcaM71AOy9MZvJFVf7BfcGz2F/wRYMVKsJ2+NiAumx
VXWRM7xg8zss/WWeUiDNnyjdV8LyPE7ukF0V16V36Rvt8OqD1s4fIDx53uqYasY8/8zyeqH9jpA0
PDb2MG+Xc8/qURp1/z2Fnk7xrMS3WtjDSm2mdChd6WdX8NbDQ/V2uFt9DbxDW4KubZkha9n6XnUv
tYOvWeXGnB3+kY/wn4Mq/1gXkHq1nPC+er6r7RDsyAV0IzR1h4JGEkSgR+/VKlOFA8QeE7YQLHkk
+pV9Nv63My+Pc4omaBfmtO7xDfrx1ziwplhJ8RUTOBuBwKKKrGfCo+OUYAIyPquyvX6YapEYhzpP
7uhq29010hbozPvnF65ym+OEf+uCz8bJCcV8JkDIT9JThO4YQlIchN/S5+miD8+ljBpPX01SXDQt
iXe6iLAdzKvMyqPOKb7BZb/wZgaBXG6BJo9RfgIC/p/U5/bZGByBdOEIxF23gdASjwKzyHwXlHfF
PhTawNnhVj0/yV3feJc21m/ENmP9EQPyFQHDPp7AN7kEaRUx1mhQIFqsRDg2UOOqqrgjDGJXelSA
IzIp9ZSg5PKWOZUxfDs+gnqia9gfcrrscDzNEC/e/K63mgvjMVP5f7rhcwpSFdmKfUncXCCiDAxX
BEZsp858k8UbVulORjSP2/EU0/LWIsFpfSQSaWssI8Xai+bkBAV1SCQpnHwHE62uJDL6cNZaW/EA
jj4pju+cAnOnCldjNM06h8fmaC/QfDc7jWNUePU6+aTZMFahS+bWnq0+vsiT3KepYdCN/LX3QSNv
PbQc+Kys24L3Ka4k/4+FyH6MKRXVOI+NmYsAqSgUmWoMjUhq87yJxWAZsqC8Q/K/ezdLsRhqW0Db
u7fe23ilp3pm7690tUbGU33208fF6Mim87bpVxs0vnxCxBOiR9y2hg83nH4tBC8J5DsQ5l2hV7HF
ZHKxBwuLrJoeeP6UHD0h2OshjjwHpyN1X3/cRFzKpCzqbjqEDMfAH5vUbk42RRrkiYDZeqd0sbBj
D7ljCegJrviV8WHLM9atb3lk8Y7EVwOkDRVidoxoC/w1rj5k2u62hWC1a8Hh+A70qWoZhCOmuYto
aisadtQakb1Jp/9N/dPrRb6DKofbnM19E4QQOuiy2Oa+OMkZinV04vyjD1NzPjXNsrRSSdY4lvr0
uvkWfqXQjXrtBt7UT9ircT0ctSZuwyiycVQmzyman5Zv01wpcbGWzNXAXKmPLpQYtw0zlGOt70ls
k0IlCdhgxX9CPrGCYXHAiD0O9p1P14OVkxcz34MLVW9XGPLUABWmK8j8S2Fps2yGtQm6xNJLpO4/
bP0sbO5gYtHp4wjxvPI75/9TyW7XKghiIe8m2TSZofO3qFpbPmOk0FhkAV/x4YMNLiKl1ihwDHkK
FkM/wlrUWemt0qhZ5URPAfFiwIf7qGOekHaZSVmqCsvf0Y1AcDSxG/I/jzRc03sI8k343pK2Vz+y
NEkixv0i23rElJaCeh0NE8LqmfUePKA+5lmLav0xH/FqZBDEzkNOjLhKvyyUC1R57RQkHUo8OJtm
OTl/Emvf95Hdz5GivxZiA/EvjuRqeZETzOh8vFt+fKC+pD/kbpGm7H60Tw05AaPHju7nOZUZZkmD
rFpWRbHJj614Y59S/pDpfCLPTXvDkCPbynv6k1PXbTMVOTGPno/LH7Z8YZAe8X8oCO5hWQZesIf5
8L4tWr1iH51gDbrgnKgKzfQfzMTliWDT8/8Vka14eD4e6RRdQ48HISCu7YNBS/rbtanqweSYT/FC
rHe5JWDRSbigvo5DXz2iyI36uZoj94bVDjlFxk8nxbhu4t0sSJvaW1fzvQlUQYCis1oDzs878gYH
Mog5obYo/1KzcSQHNJnV6pUAx53OwxZmOAJj8PVAmOn0X6NkrgCTzXRdj7khPNLIsa52p79m2FjE
MsDiEBDnMxj0mKJ5/nN2qVSl50ksAYoTr8qiUUh/pVb43Au/UgtSkJyN1XtS6YMei5b5/seY5HV9
ibL+7pxnZOsFPlscnHEzXhpml4gerqxQUvA4vqDDH5KXuZphBEm00numuC+GcPgziXsvHCU3sdXn
2xN5Pi+BnKgNdoeoH2cc14agJ+5T8LTwxTEjdMcwm1W1G4vvpbWduCqcrcBXUvj07Y5RE1AO3CJQ
3Q0q47rSEvfzIVagvpiS+6prip0ri1c8Y3tnC/Kmp7SspGH0L5KAPy8NRu++frgVNWVdVZOvH0/j
O0/A1xUFlu9y2tgR9iMnbbInSGk4heSF3MXTG1LJ32wP0XxH3zOjkM3pCJ34/xQ0S8KjsPOm3vgL
c/sSMy7uWazGqNKfCOu8pMLCPsyAwPwCLyjMr8ew0cYw7RGPulxdlOyFw5VgCt8thiSTjfbHLSGc
WyuqBNSToEEd65xKpWUjWr+52k5N/S34ofMPwNCx3EwWlX7Vp5xNOoq5LCnG++3+jQJKPCzs/ooh
f7nLy5rseXvQUqZVMAs5gWuVr24t+3TiGJPrH6deOi7r5+x3wW6L4EhrXGUzLwCQzd1HxrlPT9F8
QJQYcnuMRfjZZQOw4JOxvk6puHSeEtkbctB5lf1WVbBNvvw1AEjO86fSUIYZtwOkQdAHAW/t4cc1
zphBYtwTnrvOohaBJgj0Yd8WDfJYeDOaggAOFuEmo8arDm3bw8gR79YlOxjJcD6ulor9kAFvub6H
91ROvWLxBrfhpot3CRXAjOCY4iYg/NYZr02DH9s8tUToVj78hgBDUEvBZrzhA3rdkj/d/3/er3a6
oCDffjIPAKI9tRifBnBZrqV8UZhBaFpyF5+c8reeq54/aWwh7j0LcPwnFZyvF4MMaDMdnC4+H7OD
q3VmHZxCnOWKbh0Kt6KK2F/d8zUSVNJZE+sjTnpGnpFzQ/7LtnhSWWf4ZgWp1Gf7qoQegOQLYrbR
StO+mMFjzDzqID4MhDHfBuLqZZHMfbjoH0dBfzPpe63speKWr8AcnYU4v8nJ90xgbRJYqohYPYIk
M7NHqldevd3hYYB5UKGtDsRv8q5nMHNOJBeJcXC0FZi7ne89WG6gMLlLyyk0yR4EOUWE26Ubi5gK
4tWjt42MXnSp36S7t65DEzmaPKxpQLdP9FqxQ3xU+deCmCkuazXIIfnr+NOP31u2cF0JGHXiCn+e
obh0ZPdHGz3uSHX02Ujd7v9yZxRAMnCID3yoadeun5+Bljb4rIb2T3IHhdQS36JLeOOnUFN8isf5
tcbOjBY5XTSl2u8hnD9t5/AZPG6C+RRfw8/4s4YcpgFntj2Ev49tdN/884lqUngMypa6pB8qxvnI
QaM+PATVSqXdmtzFukUCiCQvMOd4eiHz2Gs+E0p3Cln5pic3sMAjwQYJma0qj82O67Vh52DeAuZD
D97DTlIpVXF3ZXUACzIRCz3CvwxP/TrdKI9p33nsMKeBioVotUrmbxj/6gNvG1ovPWCxOvpwL2gp
ip4kZG4oxMk/s7IANRzU5S8331A2WIGeNb7AMiKa8bc4hxUHnMz9w1aJoagbONxMGcfxKFmaYb6Z
Mqd6iahMKWZlX/GJASHCplKVeNGDFB4+vbAteyCydwR+03gZoZsYQRHzEzdagp90S5bIqU7tRA2w
tAMet23NTMdhKNOp3keq2f8xHAIlnTFEoEncFoRzampZCaON1v998u5Tsi/Ss4scmN/WwtncHUej
1upALrgfOaYIVacJ0OgKmaWrqkbDpAYqaCljItfVCK2slCDG5tBaM5ySicKJ/Bv8yMzMZLzn19Q0
iWXu/4rHmQoIvoFiKpeBJTv11+x1fHC/MvQl7e6QkH98qpbMnk9ruVLSaPxUYJfhg0AFZef27Hem
+BdgrVkxeRFd889yPZ7GnPAiKYQinrqU+Ifo8NrFya3bg+0U/WxDUCLweinnulJzy5IOOnBVKxZa
DpRihGFZQifkQy/12YwazyV/bH9d0qzspm2WkmU9H+If024jk2OT2p2b+fB4+Fftu/ocxOicU5Dh
ZdDutvUN2HFYX6fN4ZUbGImsRvlu2Lp8nKt2xzRu1vHkb+gQcb0TcbGYLXiDaLzwUhtlCPh964Vs
m5pFuPDD+lXWiOxSXADqR19T5SxNS26VSU9pBukk+LDwMvBKynioO27+klVGjkIBUCrGsB5iHKPk
P4wn3uPba2wbGebpAtFV0VPq2GCde2K3sF55MKvS4/7X9lNy0OpTuLI6k9bSZn4/mSnK8HkSXT/I
ytzN32DNhA9zYNqzeyOL5vV7t7FjnGlV/0/Ns+prfA7nM9JXWsU6MP6u0pho6xQOEnAdoAtfhduB
QgAGk5YYXHxpfG7JdaB/HCdkwH842BfPPO5nMaJP1OaK2Ad5okFMXju701J9X7DWJGXgfoQYVzll
aI1rWk/gcIg5pshsJ5sbjb4SZMykh7Uwh3S7mrx41MxSWIMVldGTeQUkeVS1ALKrKlgRB7w9PtME
Qn8VXV67QAvnxwp0hHcnzlL8cx+AyT0SEtAHFs4Rqa19Lz6Mr2C/cSvKDVWlbgMXsbIVBW0tFxGD
mGEWCe/Tobj+KnL/KEdvs+CqjQuOnsYWR3IK6t4AALriPeMH4iwHRz1og4fiuu9Dptg3H8NyTxXX
92w7wgxSuQmJpN9OJMTajKp1NXDifCSx+ECjIvR4lUe5QT1QBMW38JwPTbpAPtJNihAJAv2JXYOw
FC3EzITXdqFJSTKyI06UOpfCSs7M0glYjdHvA0Yw6m5CG5OpUQkNAg9MsC32FxQrbjarr0AAWqWa
+6lK8bj1/MyC5amcnZfk7Tt03MwOgGtl6UqOC6L8X84b5KudN7ayNmDjs/h81eVENe2LAMhd+xDC
sXV3gkkgafyRi9+2QLVrN+rkJbJ9cov/Vdp2o2FDIJPRhn56tkd1/8Pj/Ynj7iD0i1mlqBDPC60i
dVV853owvvNYuyRhbsvjfxR+jpNgPXvd3BRgeBRfNs9t/1ewhDhHht20LfAP/HTdCvUwY0AC4DHL
QbF8ZgIw/9T8YeS8Ufluz1b5yREsAVq/GXwclmBIkzy91JTTVQICmg9akMzIVfM37v2jAKahXB3s
BL2Zx85cuvvg1rzLxZPt6KR8QLm/3UhsTCtxes6zoRRqAvn8Vf0hXQsVKUJZrx8jzz7pjDuRO+ao
VIAfyqqznyvpzH3aNRRweUY66UwNsaPBe5/O9o2naZZgXvIWNF6On5QnhwejW0E+gKC9bpYnF1vK
rwNnkNks5GZyysMToyVnSviumuMevXotBsjBMcqNC+I8UZfBb4TG/F2TH7le6Xz4hukAiazkY4Jv
GTRy96V9LgJil8t7aoeUZ4fHIAgh1+rA9se35G/NsRXxEyhfZ65/0kx4shPHCU4BQFgTHWNQc+kD
ZSRdFaBrfM/wCAjds1e/A8aRlBMwgjSPw/wmMr0b9qd3mpJ5rZxmsDPolziYQodEGl+3RrSVTBe5
4y0htyJv8xdE9TxK5cpylUKu8OfuEnRftn/uD4++uphtPfjoOmbSBE64bH6E+mO8x57h11CcT/23
OOePHRMs7BgDRIKeeCTFvsFyD2Mav5yb4tNTaFQinLmF7g6/d2Rz196Sotx//XTpJE4YtZZw0jGG
wNZHYzekg2xuWcRRo6NQdUqQGTbmjtxWTynd1dHKAOujq22+RDNZkWhXtmT9qsJxaafVfPlqzwHl
g/o6lg0rFA6f7DYd+Ig9Iyjl5nuzdShM5gam/5sapwiCOFBbdMifQ5DYLwEIHQ9VJIBnHJWcWC30
7KMPtDve+6/vAE1+pGrbEilmAlcwAW5UalLYcorxw5GzHkzk6xe4RzfQ+yS1GwqNOm98E3UAADbV
C32XehY+F10BJISG4zkbRqfv9fMhCZ0JA7+MkfGMKjIgeDN+wlZAk3IfAcdK2gBrUIUEHEBapJIX
OOaKsGZeF6r3GD44zExEKXas9+qf1c4iCQWeZ/hqmfpMwxFWwEtHqgSJy/sNMGWraItheqQrI29D
xXN9e5CS/5HU4QuMqz2mUA3Wx8D67GYsT/pAauBs5d9+QgjoStksjX8ViF8SALJizfkByDCP+v/S
u9umPfqKzw9u3dBlmA2hFPuh/eqIoO0LFTCSzHAfwffCkTEdUIFIeUOMFYrR/7Cr+qAMiBOkFYe/
tVWBo6OtCCUhiNGWMABFqoXTehtf1nRWD29B628PJZwNwSdp7YHySTn8iQ7St7pj9hg8nMzF9BOr
phI/HqtlyLgqRgP7SDzDAHecLITlH20q43KIHe4HhI5oNi6W6rPLfOdV8Yqq3wZrzCo8/G07IOOp
B8RfdF3rLcnHlFV/vj1qpkQ6pBfJfCPCzrxs5eMzz6Y/Aunjcl1nF6ey0h45VPSfmRNgWIiY99Y+
Qr0N6YE2fudpeV7if2X2qgzJRRHGp5A4R7pOWtxLbwhtHhfSWRWJBXMAqtYXC+1b1BkKXHse7vWh
IxTu9kYzh0U1vZgDImHEZXTGLeW3emgKldr7EhBzvhIvfGRu+VnSPy62lu1n8vpaw+b5EeAnDptk
JrBfiWAsxDhJbQ42u5NlyMPoubipaMsFT0b5yvEUEfmWLlGzJjGxj0K4y6T73FPTvPGVPd03nD9A
XO/MTs4m5ClF197bXMeVD+QLyiRC5H408zjkRY0UpmmsGBqF7SebsGq6qlom+3X2txR1CQEmzWYc
XlOFCN8Oba+bYZn6EYZtCe8HkA6cx6wU5KUOxTl2sOGw9LqzJ7YJpJfV8wag+K6P/AqIYWrib/b7
wa68JOXijdYn0SI41Y76K4QA2rLGTjB7NXJajqj/cM7R4KsZs3Qk4mKhLQhh7zoQLvXLPfDnEl4A
xZaxdaC4OKA1i7QkQADyMhbprLn8ZRqfQ5FG2zDieE2AkTYs0wVufFl43aoCsfgeVSpQ7RoqVfYO
6Qg5wA8Pnytr8FWMAXCRPixA7ffUTWqk+WAP8/wMwYPULejGYyeC7ZszUAHQO9Z1H0iNF5pyjq50
TfrA57ImW1otBpLZWdH4+I+NPmzv6X2J3cbLhhin6H9BXXHiQt1ryl9HUQiKiTWZhE4lHdVQ01eN
k0xEuBYToqZYaHG7kLG/9PQtALef475l7WqlVFdZejnCKrH/UEldgjeJimq3VPdjh0WJPiyDls64
Wx3hn/oO8vb6th/At1goXCtZXb4IdvjGmUKouZDpOkY+MHyqKOuj2NJYz2Cv2Mi9uN6IuxFuG7PN
/z94QK8yROKEsPALchjzOmsVJJH0090R02ipuNO/fV5YdMpoFBhpdV8KtAncZFEXGiIhZ2rWKVia
N0rEaRhKUsrUcUUaztep9ZK0WOThYHvMnD1nj7/87azHXusH2XN7/Cc9b2G0gsTbTufhadk4RczC
c6vdDPXqyvkgJC74tx8zWGDZrEu/kf7lH02F/vS6yMyRddJ8FIeEVDy9/kVQRQdM+LVVNX/FxQ0u
47ZyDAWyXbn5ldnqEmbEVocgJQTWTOSBy3XZZ15AfYj9JFO+m410Rb+XkWgJ1HE1/Hqc1xwhAPux
/bUsoqo025nz3F4q9+mzq3KLcaV+kUZwBr5KndPwoOtOf5oQOIpDFi2AboNi+Hr091xgK8Mvx49B
rkQrGnVLN+/LA4EKoTF5F1Pj6wjwGlSDYd7ZJD61mMCQziUcU8VVa0rlVDFDU/pVHUuiWZDo3X9U
ZFkEdCqyTa7Ub5RTGN6mfLXiCjOxL99JzqO+rtyqmArru3FC+Jz+2u/WCPvwsauNNmrUMDq15KYz
56YISdokKh7a8m1mY3qQpo+L51nG2JzxjAB4ZQ+8HW6YcG/K1IicTQEpvtbKdx4T8VoOwz5sxGar
oZu9qyCuY0rUerLltiSv7YL+EjexrEeschLPd211pt7KPd85dyxqClvUxLZiVd16NL6HK/Ywp25T
ljPP2UkE0J9BRP/205tk3ihn8mxvl2ms3OGXGXuOKBj6agXPUbhsItI+zef63IibxNU9t9f+WWWf
4GbTyeCU5AIS076N3+VK5G7Q+VqD5Rgv5JfVJZdFXHtXWapqlq6oJLTaYI6A8VEvBYBEb1O65cUM
KMZVN1MQF0hRk7HyKSSaG1Zm9VWJ6Yfh4KTaGM1F6XB74ongM1QNCmKqKdd9KNeQJ2EuoF+KV4yx
FiugyjbVoh1FWwAVdp5Xs8LPoU2BrnZazsUvIsdDuMiWRvw63cQdXnA2PddcaMeb9I3PqCbwS3hT
HxMaKs3iE5Dzvdz7VbKuoQ/Ja2x5DANtKC3qhhwsFc3AIoqwdXDHGaUrMaTWzA6zcuFM0Lu+cJnQ
hpBNpa6ARf18gXfDPZZhtOWOngFYxr5nNh0E7HcoclJ2l8hdok7Yaq8NwPflx/pLdL6ms7gcgzIj
ihHkJz/k4yI06UyTRXHybys9SIcFkAFWSiPUmdg6qMnIuSug1ourQXuhnTWE1RjNDKV85uBP3rHp
dzsEtdn1qwB5hTkW971T7P/YtPirRSMbWb49ofjWXc1UTh3dZd+pKvJynZul/NdakS1/jLoeyq8s
pkxVV8jgoroP/W0FjT4shfThMiMUL5PbRHZIGlg+hus+GKysqqHjHwxBXdtDEBJWfFw2vjQW/Nf7
+1nlppXYSppF5C4qXbN8h0MItrvH1tTcrWV8Rrp0jorjuBWDuyf9ucc5F3sw0532Nepi5M3kRJId
ERsvQ6djdsE05TkRa9sQAaw8ATeWu2iQnoJd90OUyEN5gHFzjaFlLxOdXnbGfhi9PrmnBcH+helX
w29L3GnEpKGaQF7BXoWlzXM18WF8P7mLv5Ds3G5l8FEy0blT+5ZWTaoHAU00kTRgXEwKwZNMcou9
1kUJ2NziW9JYHsmfiMxDTHpfK/sQeS7Z1LcML7RjRVcnITSK0zMjgPnZzBEcuKQSs5sgj9ADKjjI
HUUmQ+8CBEroYosTrVHH00bD/mSKOXPL6PLJIsRepMo0XaNsgsOW3Gb/7KN+n1oEFtJx+MKeDUd8
BRKPM0q/mhBvJJ6Yst6+u2/WAyh27eeSPlyUpITTPcyl2oCSP/n5WpsvWzs3WzhtMnVHEWAO/u2Z
AV1x/bEjnfiEZGQLpEYOOU4wvNejUo3TJBKC62Wwsn1tNRKLDxjh0ARTXKLoaxuR4r1NYCANGVDa
g8hHNt4AYrN/LJ3dILTSZeqh7QxtlUGSC758K5Lxv/NAuXhydSeK6TkLdYA/V5DsO7+BsWc5+QWQ
81ULfkxR67BM8kWw5hyermepPUUzjY3fNVzqNP2PAhR6z0evk8cNY+aIXG0VwQsTX03zpZyEWZ+7
vbd7eMLJnO3GiBXJXfeHLLXxz+PdKZLhbHeRIMcq4WRZUUgryjI7AE9NDycFq0ChZrsdwH5uaHWI
QEteEJb9oUdInyVubG+YHH/TOK4rXx5ng4QT8KRqGFbdOBEsksPrA5t+HZ9tMAFfTr663phIPjnJ
hgx34M9rpig9fNGT1PDwSufbus+HBrmRgZH0uwgK7l9BiTD++SUzi5Zz53nA4KY2EAj8CivCiJxr
agNHGpbsV42pgmOG58MKAJX5n52zLuA22mFKd24tLgXnG1YYwENCpl8u4YmldtcPNhKEVx3+eHkH
aL03uWdc48jgRfpfK486DdndIU8e7zYb9+tXQh2AuJOj1Ff4PDUZqdk0YKCz5X9ZeVkwBCHEpSbc
xW/GkniLYrx4jaWs4ckjQLQiUkW8cqWBFgKEHE0H3fzql9oT9mcoCrLZZk32Fz2gJquNx3pSTTFs
jSvu/wRvdheIvGQBtJbOxNL5fPQSqL4AnWaxeyyG1sCBoxwS6O1pFteEPBfgTQ7iT/g7M9JxH9Lg
k7c0tcPL8m/wLH4mhrsPok+4bfs0N/Fz+V7gTULsYVwCZ9GGjl7XPaGYS5BV8/VwtZzV8LEpt4Eh
4KY9yi5C0WwZpNJmMhUhEARnRq6REINrYpcSbjeQT7j04AU7q2KHgXSMzNqfu8fy0QK4KSamhAGY
lPV+0mNRcMdMGVu1PgVy8Z99LHxcEqLLS7AVpiy4meXvkhspLcKDlFbNnBXOMGd8JOXr1zZpiPU0
dKw13/jI2wwM7nLdBW3HfGFnxR/8CvhBirYWGnAngmb5JfK6otb1n7NyKq9d6V57VdI+6MRJmB7k
aoSUErBNh5ct/C8iwImfESMUJcesyIUbXHzucKv6G5L2q1Mx2r6bJlShc+w28XrWTVS2ct2cs7aD
j1xVjY8Ork07z7FI8kxJcl4xr7FLblewvU4LX/VLhRA1DMFsK0w9hgz+H/QZNorNEdjJSJZXqqvW
vEshNMAqrfJoPRDJPtVU2pEHPEoAEoyBLdg8zULGzaXB27faBoARZ0sq+5VHmGFPlPk3oXBr/w8T
6yon91RIlO6nNexbGAhAj9HrYCaDzfs5zmA6SFkizbHELO7wpH0C5iuZdBA7hcSCX6Dnem/47DAB
q8XbLkNNo6LHTNBwLuqb2rWWe7Xlejyyq4BOLu0b07R8zrzutDECXwpkcZKmTBhw7DpP2GZd3uDb
DYSusJNuIPrdgqMi6blI6Xgw3Ek0Hj+Fx4veGA2kx0S2ECiCNyAphSE8hosYF+ATek7hRBqK+EIZ
s6PBFgM6P6ShIREsqU9HEn5r1w8Buw4KY4+AY1xt8vQaNFXudwAxsxh1CaWKOmjpZ+oaLniaacG1
50FIO70AbOFXkCNderDQ3Io8oAnw6HKnMX2kMiJfsHavQI2gPQXTgGiS9j0VNY+KNRKbXcyPpd22
yGeu5v4zDhddI3SKCF9HwtUc/uBz8YV9tSfhfuRancl5boFkWtuhZ0IWRRKgf+sC272ov5//KQBh
HUq/YeKeUKvgQdJ20WR+r0at6lzp5BLgXVO6HiV9pcZPxLDyHDeOJBDdilFmNMIGROw4xV+RT8r/
zOoKYuTctiOKNfhUXzzQbZaEcttW3OcPVg83o4I6sv0noS6C/UfN9gX5pXCiDGEeZjPw3FG6elvt
i/RqJ9InH+oGX8n0582QtqN6WI50qqBPBLStsplfHCXamdZ5KMbIcj0mRFbWvIVRLB09XhHYFnGW
UghEmjlNbuMRzGqqZGzUMOubQQGiAIShjpc7W9y3rTK6rjGZWs7eZ5a+bXp5F+z4LpvjMEFXDrDX
t7DPkwQKCA8z71z6TAZA78MvQmZ4wb5Ae/VIAanGlDtfSsawLYjykyiFAoRn1Sm83FR5pXGIXvjh
1CZFbVnVFHFnYfJGixEtpIm4THpDYhlGdMSLkRNHFPQ7qCf3+YrFFyndniT0vxZRsfc8HcFQ+b99
sMaSNzlv1xV6+VBmJFTaPHYytKQK472KUWoTB8MkwUSz+lB/07qZu5IgdR8KsT9WG4BE/HCq5BOD
6Pd7sbSD6lk6uRB45wl4r3RU5rHJjKCO2J9E6nE5vR8gwxZs4B54qXZEduAI7F0D8v644xDu/Pv0
zOBSG7CXQq9iHlIwUW+yRpoOyQyyGc3jL9JfX/1DRhe70mq/DTlgRd/pXJ9y7/TlwAgCb6WmgW+Y
KbFcHl/3IzgBx4ooZNaSPH1A/6zJneCJOFxWyQ/ZMiA5/2n1sgxN8n2h+etbQUzGwKFNu7vdcNwk
ZcL4Ra1dEWP7QKjAEh83w2fL6XunScGi3aI2MZ34PJsh3AOHcSRPRnD04vLaPC3bA4u5xkEy3UK6
VLXCQpH3hoVIqedWJpTWcWXp/B9qvQ56VYfWmenbbDOyLA6oTejXB7j/0tzAhpg1r0wNv1kJv/Ll
m64AV8EgctbUU+eBdH5GE7Jf+lTKwhnaHG9jk8Zf7yT0xLcQ2KQSMj+bVLWn/uYusSt8clYymgdM
+1B1EVZJYRGcM+PUFRxhLj+eIJdspN/haNKdDY4i8u2U2aw04iuKXix1A+T5rqqZIUHuMqUBF+CW
vpc1va0kdS1raqf1SihCtJhK4hFAN5fFkCjy//sJfK0HrzoXKW8+yYEld9X1U3qHfl2/5AokYI9W
8LBjXSbz/02CTCa7vyz0ifUZHoLbaLz7OdDWAmtraahFa7BB4ouKzFK0TAqW4udAJjI+WSDi8ANK
ZH0kGxQFhn3jQG66rQxQm55+Aj8YgmurWBvGwU7/fNieodZxWmyCswnRX9E9KpV7zSVz6Bd7hCMK
7FLoJbPmhpgGFSvndjHPDc7wkajMhaCaPsmmQNKoxWYTWfdni5aCBWUS9Hd0Pzxh7KSTZ2pWL5fa
wBh5noXQONbjoJA9O5Y7qDiey5HQvb5OXlMTFl5XYrBD5GCc/3Mm0r3ryzZhOzAxS6AeJExCRXgY
EmSTYs2E2sdaVDBwf9q0IO+9b0UN7OWI+0CjIc55j3EiwD8OUFCaG+U1iNKB0pB7sz5rjTZI6Yxj
uiOLVZkDpoRr5Yry2ojX18Y3J0JuBp022GjSNkb7/BqPBcVVviW/m5rRFPytJIcqmyqeFMalyd0k
g0PGP8NKK+ISoHaUaq9USt7Qj44OjrAzhb2LpdXQpH2jllekL5Wsg/E16+zNRot//rAaI3RgfFpu
7C1ddl1ljEOGm8GWkmAYMwLr68PVNhAE82EZsNXUEdbqfyNo0SiAR4HXl0G39DCo9I/22pasERSo
IDgBpNOaGrisGwHsuS+sGJD/OlfcGfiqx/G7HZFiMQ/Y/AbZWE8JKyTgYyijXRqBTT4ZcVcyvoA9
PmW2YRBYQ7mO8E6NYoOIIqWnEL2PAUwxTAlwlsLJJP9DuTG218B1LS0TR4liaYUYtaVTzwiv+kyT
f8iRVSLOkVLKWc6jLU/7M/qXI9PxR1DiQMBKfBrKo8oDjYgvmBjGHKI5jHAdLN6S0rYDfRYlfqd5
0vnBev4ipDMOJsNSdJ/dtVwQ4lGd4uug8JoXLXDewjiqHKhAVr7zLSPDeQHInTdj7GM9ZwCsJg31
BnUrdFblN+GqKqpyX12jvQt2K0b/kNP2nD+WhmSCBAIlGkfgxdfNpw3OH311u0YerBHgaxwRMH3e
HE9jbRoocHLgw4MJy57m+7YACvGAV5M2cOSYdtlnT16MGLmYLsZ71DGMEIfEjSUHTm+jIIe5hvU5
3fwuvpANDaVfXC1NyEfyc/um8AqIj+L86/vlEVKqdc9cZkbMW0xigx6q+fjF8hThScFLG5yNnjet
zm5GR8BEqkFud3pzc0b0+oou8COWsCo9R4vsn8ofT+hVfDVxXlBBqSh/dOaOVzVLzEPvc52PGWZe
NIEhDacdZpQi5ZWhM5mOhahJxmGniqORbFaqCsSGG3lo70jpLtAu131Yi4As8HIF43BEIlhj2xkU
49bzjM8IjaBOYcKyNw7aNeck/H5A/1kUz6CEAHN6qlisTaeowBTmrA4UZuuXRvDtqCXKXecAdwqp
jWffMLYnRQ/HWeYqXNcHphR5Ay+u4swlQiffFLUoSLoaiimOnmP081OQEJL0MpM4sRTjDcQfzFop
9ros4LuvEDoelzDL2s0aciA04hYYbV/ROgpp2vUZUKl+K4CZXPHX8Ul2eEekC0pNCpI8fdTIWmcm
vF0MhJEK+v5N659vqymSru+EMunEiRRknBQAj8p5ruFtLsaok0nduVbM1PO4GivB/2ux6Q2616ET
j1bpmTEpVmocCn1OlQEwR2micFE41Bi2ryVprjFVSrKtBR5I/kTolTkAIJrDPRZcENUZcqU3JVj9
w1hakMo43s3uscDH2oEc0TIEYztjQ6Pu5dv05vxlaFYdeMSLjFJJxpkWV3nBVivmCTVqCRf3w7Jy
+rfQiv7YDy5g9OoTl7ws8RrC4tFGtApEYdSpycc5wU0Ad8vNpTtQCAVITOL1UvurjcUGSm2BbC7+
MYVbw2wnWNi9jA+gMhpvRMqtr3iY9BIHk7umft6D5biUHsLfM0NNmyE3prxHPXDLIhVxnvaa2qML
+3nhZGnAVIx7bTO2Jkqxmg9k5OA1+smkLIw/aTq+pEEpGR3L37LqOEUh8AP21az2PqW32dq/vBMt
izsShh9Iu0PTPEamdnQIYbFhGj0e3nfc6MeuT6WM0CYF7pknofFlMgXnLEBNAtlWa+XlH5MFKGDq
Qk65bg9y9Quf/hLN0C67pkeOnBhfWsvom2rqNDxciPToOJL9XwFJ1hsxtA65Ysyxlbj96vMVS4Ws
kg3bsUYlkg5/zrqxtXGOxzur9BdHQA75naE3kc6h9py+ewkJg0G5c8tJdv8/EG8Ke+bjauhSZJLQ
c2hmy/RbRQkDCC8QRYiitTMwVWB+qsypv3Y/jDs63N8QZm09YWH37BptOnL27XjbNKpEoBK0ZD34
VYCv25EkGF1sLt9aXUccNdYJXQMunk18QAlykaGOM4fq25t/eIVVnv2493ZNX17pS3gRV8iuthlA
EBlD/9BxAH6f7idFMInUGXNecYZiWaz/adFMjYpD7PQh56oHQt7Z6wJ+mSjiatK/pqLhmaG71mU0
d16JEN6xuCbj/ivqtJt802waMkEUzwU0W5cRLpwwijHGtF8sXsJYsMlxlcdTdEAZ6mJcoui7XVoR
jgcQJAWMU9u/DY2uydZPS+C6qZoUzxsg/sCt1mdNErGqpgXjO6hE1DPZuXOWospob3DQbfHbqXdx
CMWzbc5sK80iLF8+ZThph3F0I+Pz47ZF7P4sD+S1j57tTcH3+kz6LYhBLj0YEKW3+QindssYI1Ba
Aj6A0ACYBBQq/a9w7YB/wwr3BaE8Dp2uJiTUm6NYI1bwq8DsTsUd3HEzrBjaHdmch86qYcWRoa6j
QX3GdWCzqj8gMeIaSLdjbiFl1wXxNwd+agA3qQ/qsTNLaueC1x06+Ia5RWEXrdVKI7J3b6jYbkyq
QTBJfsK8aJhd2q92Phtodeh7Xw2NH2olO/InEwB1bGc9xlaWY9r2PS7ZO/36CNlZzuPSaXSMJxT2
byi3XOjgoLrrTR8uIPv2i5HlG9i3/dqv62DCNLQQYNWBh9vuK1cG2voV/YRJt4NJl1PZXtUHwptL
/MKSpqVM5za7VKYzCp/UzkxjyIiD6aS95rMTqNlcTu/Etv+H7RsKHSj2i5Tlsb2XaENIXSu/fRBM
HKDTFqmGu5/+mu8fzps5tiyd3d26gc1hIEziE4Y8qW3L2Ze8q1NxwVPXYtmOTl4i6AcfGQSRzYFM
WYKYDaMoyqK0BcsUPYoiGB7m44EvC4Ud2v1oBfhiFjNSM43kuJhjOLDb9/SA2DtGtZXArCZuXZPd
WSr3LTjIDTLVyuktlA1CtmzF6XQqeLflGyy/aRjDRRpZImXvBQI4q9BDdc2MNqkF+nenaVj9uvdp
FAxgUSkF24mO5ZNuvxJFJiuM1vGWUf70YlZvyrZoRKN/J0suzeOdLyhMAoJu9mWEnwA7YDAL/0UE
A3hM6HFidOeNmbUExZrOlrmSyFk37J70O6slvmkgtWb/C0C4yf6wIgtRfktbSZ63u7VvMZSMsW8V
Otis/lGQiNt3BdfU3V/UmN5UCECN/t/SX/fqmXnnRq8xVXdcYHsvT5pYvaaMmh1zh3FD0Ua/kYTn
d8MlivbYchwsluByh3u/c9ynew1W2zmUI+bVuZ27tor/R/kzjBzQfNJFL4PvjWDH2UXhalLQvW6R
8BA91/JHilgQ6UDSpKnHQqFAILBYXjcwpZEoWXKzGj9t9BrUtbM9j3coEnQxCDxjeeDNbiKBE9tS
tpd2dDdtb0sXgpgFjLTk6+9Q5NjTy/G8lzBr2mnWE1H+VHQ2PXKvUEqGEgjLzF9BPOt3vpNPugjH
kkC8bLZ+4uoFouSQRlbgMZGFoZP2QwF1C9SZ+klQkfMGdRI+Js1YJbs+SJrfpgTVXeI8Cm1+V01Y
Stn+3tDbAVixu2YWqwU0mslkhX7Qj4FBfLoxKXGxX4zy9ASNBPhAIQykz9zAmQSD0qe3jfsVRhut
p0+h0Ci7p8tIdtIyjlXvKNNytoaKsfxozwMCIgDtIAPGV/zVw7h9nvbi2Y3xCJQGWKPR2WuimZ6t
0K1kbIPZzur7LTzLCFJH/9RN8SfvMLVtxuXc7r+w+opH825DBEzWIxkXmt5n9CzkeKuIMcl+5/kU
BKwcifqODxJlVH8vKhyDnYuu+WfxWkFJaYWO7i7RvjGOz+4TZr3FjWoGWN57hX5j2zr0uX6/zgMI
ln11zWGuY+9geVxy3qWZ+fyVKDvEupacn1cHHe/UzjOSvoBL6EtQ8qH0JKrphId+E5L+fb1eDtSE
S9bvvYxicCbnlCChieVSkzeYgdKofFaEgKR00pBrZFttizqFhNHjaXY7vfgBqFmMNLdvcgKviND1
KH+MfewnPw+o1DCXDiUHiu5IpYNcW+P+ZYoY6a9ANb5B2XSeOe0O6Y2Q1vaP6364GU32lt+dkCnv
PkMVl9la7u5zrMdL2zCkDPAWwCuLgeIGFrhLUDiFR/nJl1ItrXFl8FRbNyJ/sZHnly60/dOuPrvf
04iJm9GTUnGRpowSViqKU4MqiPRhOLahLD9knTFmbfl3aWoUzdHuGqrwNcNIDfBshNxXs3Lt40tG
3J8VnmNTYa9khhXjQGv5cYdO9glAp431GE72dyy32l5As9Web1lgsW2zDZh0qg7NG6Iym4BEzev3
l5W3+yHO7GElTxAqS0IvnTk6SgwiOLPG7lxtDGNpGeWgcerehFWITLF1QPOP4CetGqBmZ7sFUZbQ
ra3cOY48ySCeml70nLXNknxt5evujo3Fo/2cS+oGe6MriVD+H/nnPQgSQmkEtv7RhJcB56cBWnVu
6w61tAc3gavn7qwJCKUWkn8jgjnr2j6RWzjrNiM1f5DAXqzH3X07Ewt7psYmHG2R7quQ8vD0Sg+0
F0nk1MYrKlCAjbtGNw6OvTa8sW8WwvBEXaeE/tecNLZEZ4OhbrLCd0DPpd0MWI4u/24RGr3i8CnQ
k0GwiSLisQxPQ0JavyvUI1iDq6RWLuqPRBV82YmN4A4zA6kWlKl5OJcYYUvCfaeulLDPFlpEB0AI
e1rjXlNSXe0kF2Qsf1Iu7D0v1EzOixcHUkZmm4oox2nkAjFju/FfMCiSWZNmOD8FhBOV/q3cUdZc
ecCyR/bVJ8wTabK51iJT67h8F9pgC8Q2melQh8U4Z+NeB0qRnkTIm1iM7b9CrJFgTt4maunt5A/F
beBS2cBOa6p3ZrpIr2IdqsGBJZy0Vg2pQfQ4Hz/GfruFaHNxwirWexJ4voN8f+OEdO6Zv9Vq2cE6
IlImpVqNPAtBPeTmhwiyGs3YQ12KovixOE4Q5ibQ702BMoAc69PIePPxZDRQWfbE0nZK/Z/nE/nl
9NOngXN9F2mTn4iKjsVDrH1QQma2+2Mdt3ZHdUGTSHiI3UCJRhya71AOhgk60/1Z53Hp7Rk398cG
Nzx1is9Z85ABg5o1chFfKo87hKjRcN/A9It/dXWQMVZZxKlxxbgQL5FahUvrfzFQSDCz+zgT2fB9
HDGGpF7hsom+i3ghPd5bC7YqxGB27iXlnQqCd0U5SxU3RSLYOHjcGTraGnORzfTQo258Q5SMUYwP
csZV094AEQBLuzFtkJ+XJ2sClm/BLs6aAbZ7WlMvd+pg1lE1d4kjHt38V/vy1BR3VfNnPRO/VWo5
L5JyM7BQOGhSYjryhT8t9tFcmgTXpWVR9h3pS1f8qnuIYxyrrZzRebpcokI2PX1MU3OobrXDQ1Ff
dJhenFGff+r5h+PiO1Y9JC+8cbabDR9a/mlPzah8aWKADI5K/MtSd8hE01mWSjQbhcsdmY8t74UF
n+9Zy7/TE3lTgLvEWLR9fIfibe4o4L+b4fdfDsHSGHSNgG+KAVYXrRRMzybGzIwWCX4PpqF7MYDA
X6ZbZ4EeG+jIRkPjJv+xsjJc5V9/EnerHNfqOXBPmo9oiZID+kU38H16LH9kPSAzkCUVHfkBgv9Y
UcIloqFdKmuBB/Qhh1lyHeB+bp0m545hjgFK2aLKCws6/77U019hmDJsakAYGUO3BrfRJr2a0ZyC
DIPm1X8/jYKne/WpiY7gdrRBZqeYtYYPnjp7GB8LfvgwEIKCxuWpezmFdlqQgIEOkDLrkehbeHDZ
B4K+4iH1LVNjmN9hV8CYOxeBZARF44KLwXEDnZXpWBacBxH9nZUDecZKfDczFWVxy/OtVGerLxJI
waK6qPtyJkXpiaIFtnYnE3XFuECsdofI9xyanv1gAm1hqt6IY0l8eSfVjs4gfgzvnDk5MA2zP2OV
ORC5S5StrCMSBxTICBPSvIE0I6RpGlgb9Q2RM/0UE1RIQRg48mkiILeuJA0B4W577bPFPtc/Y66B
VBzI02aGWBQK69s0i7t7th3DT/OaGOjPLHw5kScLEtjNIYjf5osF2FjkzZVgO21apcpkZArDPRl8
EcwR3ZAQh8rIbieta5PWZaZwP9tOaeok65/LueUVivT+IZJZeGnp534AyIXlpEP3B7XpyXoVAkzh
EZ5Ll9v3eBSoLGajne2rS2oRNLMU+0q4Jww3S5a6AKZg0nCiyQP5z6Rk7TH95pmm074s94rh3y+x
sMF7CiR8EHDy3fdudpfyfwkkFKYP8ms9aVd+zbsJHAzpoYWkkA0XS5fR1/eKKT5vzJrEKQF2ZZQf
NTdRS+5b1YvFoOwy8hjmI4CRBSE/1H6iHCtuEF47p5JcwfXq5M3mrbilSXH8xmWxxA2FZepUybVL
NNhoKT9AcpbWaqFtADmJWxHVj09H8OH0V5MG0L8WurrA1Egm9eR7FZXLWiK7liDOfhARu+JTIGLO
j3kqzgFUWYuHzQ5zH+EUFsqGz0IZ008J/ebEf4G0dBe1FGTmdRftxuwao5wxbS72Z+jymQAR2tZU
ZCAhjVkmgygbkD7/jXQlrgh8ZvahewrGzZuhtxHoXWqrAhJEaFsVmMluIqSu1Fvq75N7dVYND5UH
qZUuCh11AfBq/M7EHnK6y0a+n+hb1c+QFb6TM0ZbdWxqNHpKq+tvxYYDKzwXllUFHqRBMmxjY2tW
+9dr3A52N3NOm0FwMugGqm+UEiH3q69rptazDIIWX0g7gxyedx29Vk7wlQB2E3PmBeC7/Hqk49da
1A5PuvjgFSvkBioOnngssy5iytBI11Sg84YLR8foENB1nRB5MR9eM38jypbYsbkKsK2e2ZdKJzu8
5bKCplnpu1vCLGbzRLcGh6m4HjgG/befDVUKJIBtHFZ/AnqPzGCNkfJPV1lX+N4vzqoJ5ltBn0RC
eX3duBWjMsGf76LRK+WbO7MzLoQbugHRivITuEAcxJYYVOotmwh2BbqSahnkzHpFWWAm0qMbvYw+
9zMXScdgi8wLa6Q2mC94SdpBWwbCPX0P6GxiExykfl/exjESq8ZAc9y710XoFfib1VKrGxaU8sQS
6SkOpuO3DMk2LvKZ4/Yfh/KRiNw3QllpCZnEsNFj+W0fv/RvlOdEAMWQ2PN9GJiBOsUToblhmDYg
cq3qjx56isoKhAF1vRoq0MR4VjAs4J0VdrIQN3wsNsJwPv0aaWqIXTREQ2mOk8VNLArzt7FgtMZh
hnY+HzMUJfrCGehNFoLix1X4pyc7bqco0Uxy9OPokFp2yMR55vDTR5XJoy9FDRZCNuiPsPTq+vs9
f6G97JPX34XJnFrFH7VId5D+hzvZv5h920AoO6c0Guggao3ht9V3ql4aoXbbPgKNbBZEogQE3H9a
hAB8mG4YsJdPZ0k3j07USuReIkP5bBvihBP9b0wjr5VDBO4EHkMF2u8UY4Iylilv8TwdLZkbx+LK
+2TIWfhHsblfORWlnN1DPj0VPSiBa31eIoHpkx44qZwi97q0UIB6IzJC25JiEJYvDx025ac+H6z4
HRen9mKcVxG+SqxBi7TDZfDpEuc0/LkTVxJXeJL5MgN7ugp6QR59K0fGbXxGrcMe1fRGNMo33jQ9
PO7UIVNgSCkFGn7BdcwE8NPiAP6XECWQB/jqFb8OI5tRKogaXDZ0Z0vIf49/oDHycoHSzgF/gCEg
kvKahyqTdXDwtMI+J8Y4mTuc0Necz5ytzBpri7lR+4Ri+LI6d9UI3haiQHOVHy44z/NOEAkhcM3+
Dcz6L/b7Y/Ys+xFiJn6a14DK1CjMAlzIYgWjN9MEBaowNFMubUZMDatB14bHo9hJFS1zdHzDIhln
tlzOYWAYFCGJKPu6GnZytiaLRQna2eT0R4/YRBq8C1mN5xLyPOfzwsNvZaH9xU4DRQR8DwcGAf0P
885EISIe4RfQTrQKZTR/kp16uJklcJbP3hXQPX/AGHz2thS6IODvXVpUr6OFu/mjHNPANDRoeCLm
BRxf+E/f0iV8aZrtT2sz5ntdbdWkxw/7kGNs/g87c40M16IFlVYENuVn8wm4Gr97oTdPXpTpz6uD
4H3XBxFrC76qeuK0MNWWGpt0IpDyIjk+wLzqIK+XN1+xZPQwwOvhiSjtxR2IKzZXN0rGGWtJExd7
WvKGeX2VxPxlRKUp2A1feTD8iRT6Qcch0ykTFsI9yChZkOSTvA0anSDpmWpOQdoiDa20JBWiN9yd
8B0PDc4YKzL/JNRZBiXC4glpOpeGkvmTop2HLEaFMGMXoFeuhQlaqxdhW9LiKuKlUKFTFo3eKCUQ
TbBZ4soXyoRwUdSeVOXsTySzb/Zi0DXsZAfP9C4OSKaeVGecSTxCNNvHDQPy1QWBLB1VP5NPuRqe
/7SMja3vi/JEBatQfVHqUGKj34I8lr55fq+Mk/tpJZ4ljNgNem+Wo4E8RZGw8RKwnaxTYIPrQXXh
BBY/KryZo3AfANvssmB1U1YVlJ8zWxXxFBVFzqir6tx1jtfoX6n10S34fSA8uLTN5qGEn1LV4SY2
CFeoGFxttsljmIrkaKGtaw2IC+2S1zewOfD0uB4dCZfABdAR3jf9yOvxN1P7yQvm8Ulr/llHRzep
9IvuJj1J9F+E1omP3ujqg9XGS29qvLxNRiTpOwXtfzXLSczusaWXCvOPs5RFL5m8CqIL9MEcuPHd
DAgNflsRQsukgsY1cHRzmeRQb3PxHS7t/kbxmmetPbDZjE0voqIDfNh1coAq1GNashalvpJkrFPx
RJBMbP/+avMTwmED60MAxnxo/9OUFvY+RgkMMcoddidAeoqL6nWjmekG1dLUeH22p3Dn/8P9nAH+
od/tpPcJhV7HkVAdVvF3YxQNxngiPExCkv8JV2YNcOgSafVos8gXAo8Mzo65UblmP7KIaQH+84M4
Xp7m7Pt62oxMr5bKlNbv78uehpmT7o5R3UuKOLxV19FGoIuBj2fHg5YuNXHnEvu8axa+e2hd2ni+
fZHaKhBpFGF3L29Z1vuHx5FDVrbNE2VMcmsbq78uvWf0rSXyF3wJvJqiq5AFct8dpy6p3vQ2Srat
jcoLNCEDyaYxKKTy0hKEozdzSuUSfvPg3ay6gexuAeQ1Fhb2EoLx3cz/MJE7P3QMV2SQUjIzO/cS
yC61McQTTmh4JDz2mOU1cI7bNmbFevkcaUps1EuJfhNI8TfJ/3nDg3d0lVJ9c3G+ndexwy2G2GhW
WZGw67d2vWrtf2BCFxTnlO56T1jbzzEHYhi+Yxz8O7YO3nhp60qR6ypTxYOb9sdkdc1EbFZ6zZuR
+OOaiI29I3HbnzrQNxgkfFhFw07pc/CluXRTFVllwxxVTtO3xps8/p9MJJ+/HYwrOphQeRxlOQ/x
bGlzZ0eOqha05cvzIquD/PyksIqvaZILgkw46OLjn4cfJsz6gkIVvo+tFJq9SiOugcKxii5xg8eC
ZsKYGyHmELAwUkUjgYwk0ZowJP2xqVSmACgqrhNz+Yp1A5YUrl+R4PIU293AUHQ1I5U3L06kTgCB
daL61hG8bM/zMV01ra8harT9lMo4BuQTZO9CYADv2vi0PECrv5VsPoAov1sZ6HMZD/9QXJvvh1Hi
kVeT0gycOKUN7lR3HN92x7sipnFJmqjw8/y86Hmzq/h4NBy3Snl12n3MxgaKxaE8EbJDetEYwdZ7
OrDL1AR1KYMQlBTvo7CML8oZ70F2bnA9yAL7lzxUMDVKB62j5ycwyBKO4G6wdRf2N+W+4NalOXYy
ljZatXB1vxPAZe0zudmEJRGCsXi8ygp8L7VcFV3nVzmj9SQT8xWmSmddsihdOSy8uaxKbKSCPOqC
PLPW2MgXdrB2NFhPYGQMkqg/+Y0C/Q2s9+Mk1oLEs72n3mMNz+dqW60SZEX50XePgGZaOg12Tj5h
z0YWckSkk85OJMwENvi9R14WOpGXAnzDR2p/tB7qmjO9yS/WHYnQw4ajCSa/7WMvr1aL5hceK7ea
WJNMVhKvuqFqli2CzokDOP5+nnRZbzQOnFUCLyMZ7O7xI5fsxU7yPiUCOS1LxZ4jeuJ5NyolTCRB
UDLJCD47uNebQSBfHk/UZRekeORISqD3lQr2GAP+IRhB2JAJ7zQuN1LYyUD6q+x5Y7txPtrx3hQa
obD3BNZJZVjZ9jcfH2/tZScqvXRvyPokODfDet0vPzMPMF1iplhXbjqhSWJ4Fi1s66s8mmpnaMYn
gcMBIBtW8oEgu0cQtlOjkJd7wLVQPEuxLtByn62MGZBM/cD1lImIpPb5ckrDHjNo4zrkrHYWyXLA
KnXLVhqGyFSNYGNqAPrdEIwcXkjeUW7eBjB1gNVs+1HXDx9fM4h5qfIrksU5Nf/kh5jZx969Ivlt
iZFGOmZ6hcS/Y0jVhGhpa4LBEZx1UmLnBBczLt767z0YmlS0BggbrPVWFgfbzGcyDkb2Xk8YzM0U
Fa/3MFt/f4MEeSH8bmQuAQf6sVEi2ieE25TOCVWqAdAEal+/dYsid2LkFmRFk/ZoEJ8d+SPAiitU
RdUG0M+uu4sip/9UXt1xH9cQJVD8VsuQkiyxktyyHBdYFoLZamd35SjM3as2MkDvw9XOAGftL8ou
JSCkTQbCokqe5/k1//6BBXwGfu5Q+2Hdnk2SZDY78qg1N1FT9Xcx2bLCRBW/HxL4REBHu2Wgs4M+
KXvR5E+f55T3WGKwkGw5wecDf5j6G9qXR1fLpIvBWt4/wTkq8qGZbCYackRKH4tr6QyHXHmYjZNE
XLtHf4EWbixg2hmgIa2fOOSp462KUcXaRILxYmvKvEL38poFtCuHGLmIi4molwMV5ZjYymwIon9Q
fCTMZ1YuZANXgrqgrDLpNcIVwX7yEFfcmPPZolNM3g2iNHL+TqmWPZzElhzj3Et073g6C8GXWIHe
zTnkosBpduAy3ywetvuKU0TpyehIvyY/FGcL/ezLkijzGOez77hrYnlxyFvQVjNxqKcUE8Lt2BHH
l/ph1aLGQ/DNaXTgTrNK0HcpeSp97QnEzzehO2NPwAWGoAkcva3XBLd8wya7qLRLw4O9iCPGC0/T
pfrcsattO9nc/B4+SAYKGsKNStskE/R1epTRD9/q/1CZipgCb2XtBB1FHYcASs0VFrVUD+xBVwDB
6cUN2Ws92r0lue8ZMltkt4ZQJXNYFCifYVv3/dWiH2hjQ5w7gMiLHq4JtxPkN0DSvcJHXp+gsAPC
NIF8jItBJv8BvPDRnOhgw8OYX5F0zgw2/mYNgH0NOwOuXHsuHAAWjsD231bRFhBxyO4rbiKtqpVX
WhzpkNCf97Jk6Z3PmBAKp8NRTooKYs5rgkAQdNi56MvWpSybKvoTSwaUwJR48tOhzUy9hUNR6DY8
jamua64Mfow1dvHOFKBZImnZCvdZ3zzNX9EdCbLQaOVuCiPBYOnxJ7S608f2O0KAl6pLqaH43U+E
xYA+cJ1G1JWXpvTIU1pBDQLK3IP3WyHPIzx3sLbts1l/HYatwKKfX+LHu19ROyM8+u6Y+F1YUgCF
owC1o2IXdwp+orjffEihJi/zXLIAeGzxLPy3ldHTOjg2LqFeq/J0aZQapbhpYyp2tWfcoVYRmm2h
1EfolAplgD6liDoTj5/nffR2x6V42w3hpdy+Zi5gvmrNHlmphRyHgUAtqYC6CcRYJIYPuh8TLMGp
uoqFcqBmsUeaW5TdM8uvrafzVFmz+ZNVH/HoczgNl4wYvPVjiV/AsTklLKQBpByabDt+nHLQ56OS
bP0ad2pWb+0mpObkgukXfEzzucVo0y78uhJiSeXoKFBuulqRrS32QiEDGJbwwVsJolZrdXhEOIPy
kpj3O4R3d8vAqjklV0aHXgALI8m524D6EHFvIr291Vj0nKd6tmSB8kIW6liD73yiLpQy7a9z+XXF
qSIJ9kb8d3bscjwFQDAfqq4D0uUZ+MuQogcTBmlXjhHHQBJ/I672ktKJTlXtInnhCtqIDEP7U5Bi
BrZMHnhP7FnNj3aEIUhU622Cwu3IP0cNhDtb/jUcH+m2onNkainIk+HsrSSSOXG30mteKg6D/wnL
6xV/5RYF8j+tVOnliRQqBvzvLfy1zkoYEufbgaLQZT+OM58xTJxhsdhv/QV8Ya2gyYF1DstJGEsB
G/Hs5RWFK79IuXaFGsS42CzYw2uGDjo7pjtPy4ojnOY4k6mnObO4TRbpY8MsQd3XCIJQ2iPgeKSB
HVl0rrzEdPUYBeiU/BI0yz8rTX7Sfg9SdGl+U7/fPUFkKaF2kV4HNG7gCM2PgBbrwi17MjKcrowt
TZ+u5YmRDnvFN8gmYjWtrmG6L6VGBGpBAPxpGUi4HxIOXBK7lj4TpxvBDI85pRYMzsl5Nsn40nu9
Sh1EHEtbUlmCcTFQEHZvc7cBuPk0aMRRN+9dKMrw9sYYrvNYdKzyO+0ZmkZ+Ez5wVAUDXbsYTcoI
udWD0v/0HdBRowyQG1itr8VKiPNmVyxPBeJy1ycgmLOB/tcmwqfg7bbWsjfoGPMTVirCWglfb2fp
7yKWHFliQ6Xd97ezRTAuBQ/uXz19FM7aNFjOhxwKusQ0OjZWtmziZMf8gpXccGY5sa/toOWl8I73
MaYTPmtqlYBVnUdhldXbtPCM7mBIFwaf0WnjrjuYbBu7Hlx5AkXvPlpGSU++S86d1HLLlpzX9Ou4
U8Cp4CiwfLFHaezlFMbNlJbfNUeX4qkBJLSfFHGZP1ND8oQvTfLYwitmrRqaC4xU5Ab+3U7FqtuK
qg7wUgNBFEtvpmoU6QqpJcRm5DguWm19CJD2DELd5phNQzUnR3gt8Gm22MNh8RS+aPGSSjXz7VDp
V9GjzfoFAwpY4/eVPpT0N4W3k0ZxkgKJLZaT2uMRHZxMMrZW9ifiGpY6PAlMd8yd0JLNU5aZJ+Jd
ikM+ulO2TtTXb19ycRoVIa18RTFYTSBbg/kWlA5ixcYEef8/TvL3WdruBeTlGLvCKg2Dt0qWo/tQ
mvq8EVe5jutxuIZgauciyUcqPqFYdgDuZvW7F66PUpJIz4IC7/vTblZj1yEj77Ur+IYynoWpmyYT
Tx1iFPWGnNEAYOxmQ0UeCz95OF8MxbkohQIg3GFVC6DgnY41ZB+3NlYZ+By2yPG4dmBhbHQ68mVl
y8RLK0o4ttU89jrGmcxSttrm2ERb+n58i9FCBRpP3/PMYOSDXJOGxOuz0Z8G3+R0cWGHs1pD7GPT
h8E/xsCy9OE9ehifyasfcyB1lezQUzcr9pG4KQrZDhkOebhCd7Wc7FiEWNauFEW2l10JJXE/EAuW
OuXN1NJwFcs5ct/EARFIPH3Zd5jE/m0ZHajhC1MYAGJXhUdxKSJrsKoUVuQ+lJKNYxCfH7HDEEC5
SkITXbhz4S/0KL27m4iSFpY1HWQlICkWItsUiN46hkHOFX57dhqCi5rdL3etYfckjnp8z1D7+EFF
9BvD8enEWRzDahSVDZ9FokDrbnEkMQD45wM2XLef9Wq6FR/aXq7swQcjy66WpowPrf9Cd9vQ8GIm
R2kmhbCBnptcIEdNCLC0yKYWZlFRK798ZtaAFDeRcX7norpbfIUs+mrNlJrcT9OjKyNHqjSrdg2V
gAOgb2fRtqEZzxOioEfge4rCm0nclFZrNeIYOJFqfazQzNmqmkSq1YERtATkIZhj4tcAJPHQN2Z4
SYTL5I9bs0ZaLSXeNcat/bAtSxpoYgi/LM5KUsDbv1VGYZRmHzUdWTcnn8fEUp8VPoK6+dx3JL/x
Hq6lfm9AqCH4rHJ1tr+bm1Jgvocek+Ssj8Kdrg3fnCmXeCBgsC8WKW/qCzcXYPU3cssQ2xWU3X6D
nHp73gqkUidzxtWOi19mhWKXhw7YAnHTacYN1CDQ2qxWWJflpnOvQjDRJyQM4F/1d4lamRbUt/63
AJbAwfwuKjASvd8eYLeSfbCL/EJ36R6EQcroh+0mBBjEhyat9+pculgOGAWliDyrPQk97bMCkRAj
oOT2uPhQIKJjm3fwZb5dyvuaj/s/HhiX2NOUk/8bGI4CW3/wlXujorIfPusbsJbbI2Xh7m9wcltD
QiYT4yy77kgG8Tha30/zHbXZt8jaGMzpm1cFYU2lerhSnrGJPtRQu5PYwofQPA7dphl1TajYaM8u
tD4362ceOeXwpHUQseyGYokKkBkead5qOWLhUau4MCZdIfU9StS5H6W7fIn/5LxpGqE+wpmTlghF
qtIPONnObRLbJutM5JbuCopFdjh/nWl4+MH/I3Kgn9tmvdIzRlLtP/ZPcKUmkZXTNr//RK8GNXpm
rEcOi6vZZiOYRiSLu0b2bHRfIDAEIwiWFB3HzBdBLnt9MCyTOhgr0SDSXR6eqyEd3mQWZ8a05w5D
mFUDOaXvoUA0RaZtWdAPwQG5DZSNSLsMbWnjwQI0ai6/WmZZAwELkVZ7RZVFM7U1vI9Tzrgntomh
vtn8P97UJVR6obtqd7pEN/K6LWneYCTtK5fDU5oRPROJZXg05qqbVLonStgfaOhysULkx3MlD+Ku
1COViHX1sQt+6/r7xWGZA24uDErdEQxeGLfTzEc0Y4T1+DkjLS91h1Q33k6bRiUqc6e8Hh6k5iDF
PZ2ZbwllAheKm9Z0CgaAru5/STZRsjImQAQxgjJaCkiEO+NqSLN7z9VlSf4Lw2tr//ZTafnEB4B/
pLH/sE//YF3SH8fAEXZd4z+X+XT6VMtShwbphBURQP3G2Gmd3J/67bEIUD+JKHvqv7xdOa14kEli
hm3Wqx/Qet6et4ePxCzD0ZLEBOBLUQloW0pRfTX/+JRN7J5Obdv56dCg/8atD8gczpeyhbiEPwO2
JApJNR1cgAmuav8Y1FmOTWwt2L+nhxNVEvUJDuTthTJlYaV1bgIGdvRkyeQQ6+3D6SDa1x0Z3PzI
kPSTDFBPqJiWMxaa7LoJYTg528ww8ISWXO9KxPMwetop3cmxcvWKUUIEUv9CSxWD3qmCrguAW18p
aPUI8xkLah5pwScEwkOV5q7/KH1U4zUbYCLfhIpgnft0NBQ0/CqdUYnXUkZJcVtH5z4A/4Q117bb
JutLKEE/IeYnR4Nt9ttAkuF8lgZoigm5yn8pjMI6PZeSIxZofrhh1vJ98XUj8N8i+NG9Qtj10d4j
v4c8g9bgnPc5/OLvMDezfrKS+AW03Zqp6h0zppJ+BxKswTiDlu6CXh68s8cLchso2G5tM4bUkgjx
m/aHMxU8NrdoY6Jh/p/1tCuG5107MpQufG3nmRF7rpGMGSP5BwDpWt9Jdj6c0humOSe6T4uLX1mp
v/lme4SfwG1CKpDbMQ2Ct3/pR4bOBg/4mmD8/xhk9UmSb+T8CAVssEaivXCiVOlsYURPgUR66jFV
G/hkmmK1/Q8e2/GhSoEYGaBJmS2Ud9KqsJnu8F7PRbx+TmJy2NVIN3+2bSCZZpkoLLh4+7Am3IOw
w00/fVYSZauWcitjN8BsAbB1gtm1kXn/icq4O8lU/xXOWJbwM8hnosliwCw/tH3j0YY+P6HLq5R6
+07ai8wfZUhviOWDj5YVHHnPIanCygt/ipwiZ/wEz2oAp6xi03Dr0qAMEEDyOQO2dTSJyn9FJ0f1
lWuBZlcI2aZ8XdB9+A/Z/xifPU6gRBnmEi+Blvvwuo1rijEvS6vPQqgDMQnEGcsh3iB+E0cHA1EQ
ApHuAbQN0bDB5fI5cmqvAxNApF5s+nkRxMUvZfjpOpRPc7Penoy0aSw1oc1OUHjw3jc0ahwLxZO+
dxV+LcrVchGM9nZXGlfHS4W0VWlivibtDYsAaFmaOCSB/xwJ8NgjkGDtoL35wogZJpFWGaqIX1Wh
kuiNcvpXTRXA7rmOQj8t1OOfuT+enquSkYpdy2P4yzF77Cmdn/CTF08Hhph398Sakjf+2kH/9IAp
6VXddQsds5RRoXmXY2gAT8dHThwhwEDjFT5GXvoy0K6YDTzM6ZqW3Endjb0J1IokqyZTRw+zQoR7
XNRZTjs/xFkqEFJVE5W913MgCgoBbqrVQtUgLgFjaQEiimCpE78PuE8I5RzIuTowbVrfUJqXFHUU
6/75gomn1gtZU5FQHyLhklUb5DSEiDxNs5PxJhVfS1CloxvBCNFNAYGVJPXgTCSX2JhARWDq3IS3
gULJAr0+KO2mA0VGzkAYObyJrZjS5jrKIRszb+z/oikNh/m0Zfvn8rDDcDZK+fFcle7X/wb5yNPW
BFRtGvR1cc7ohodmwMXmk5qUDQW4Y/rRrMTrTqknSwqVxZwtpddjLn2KjCrb8SGlm9VNWKadCcLr
McYZtHzwou2KGAvDAqbWHzAl64HdsnMpo3SKxnFzmyjuI8D70qROxpE8Apd2+H4bkFhV+UxucR8s
KrhOqe0fxcEt4zSEXBN7kZ4YwqVoeyipWnylm0zrHdZRA4YrjLjsakuMK06r2JwYTDKaFXJP3q88
h8LZLL+q26oOWHkQLhW8j3N00ShIDj/F6o/RZe6MaFgmoLePk56SdRV9jOtYRlxzjPTU353eNsJn
4LnnT2Wo++e8CbrGm6Qr4Gj79GajsX6uCvy0u2jvt9hok8jGS10Iu9odFyR7Mn+hd9HK3NYAZJrt
ONN2jaR3c7rfOKFQuWav5DMEgr5qHhtvPbKMqxMoZrQ8VGu+kBmd4P4LpguqhhVUKvfQ6Kr8t0uZ
jBHsmxeCRpovYweCMGPDcPmjukg9zjzZ3miodiMOV1OAZINzZ0akqQS0xAMFurwUo31yF27s4HGw
/q2UlQOib7nTw+haT9l8X44cj4MNMZmU/2Am81VyMNxePW3oJrlIgGnQDNSSsmOrd4Kkv1qskn7p
i4dNACS/vt/ON5lmdKGlRjq05c455m6+gSiIzCtK6FLU3hacVb3umGa1eWu/Mx6Ix5ewJ7dcEQaB
MiFiqSKtWzX+KGSEa1oL3sDEW1cqt4cnAA7tLXipD/Brvqom+76yi+MVmWJHoekLF4cYWj93kOWG
cHANILoz7utcLv39iviUfZXKorvECtPenTGH5FM4GUE2GPd62H4rvvxyUjn+venbYq2HYLwfpzIl
E1zRVpKx+Za8XMKkQzIjByx3wv3CNoEYgRhDe7lo3Rb3VjNi3JBTDx4DhD6NdLbYowUQRAyWVizj
W5NkSk3VhDFHGlin0kS5bTbmqKJUPhIDsfrz6Kf0/XLCbEBxmt9Ez80LpoZqb+gBGiCx4tKlO4p3
Jj7w2BOnDpPZXW2aeB+HUExX6BVzdk/IErMH/ZuZHQ0aAtTpeQA1s8TxMIRMd0NGvYZnbBbqet6V
xApAPCe/N8NDYBPHpF4nZu7hb5bKpnsvf0AnQR/x2M4XY3UYRQ6XwUkMqtJ2yShqkoyzA6dJIjnT
8oa4WvxuEr2kmQNcSIVbRYVS0KcHSF0QnXfV5XmdGOwg0lfiuT3ZR9xNx78DblqzOHfxxoaSKYDP
8PIqoSqnO63QKDr9/lRq7JRSQq8n4bPvu7dXPIhq2L2jQsEoDpnEIj5W9Kbb9rkPUskj+kgITPAM
gAawRG9xoFNhkdV3pOYBYhoTg7lyusyFwFskt0EaYbSIA//OAI3KiCmsXrUBIJ+bkm9hNfKmpupS
MwGwszJ/2bsAvB5lLoKaie9sCR0lRCSd5KRGc2ul4qwRN+AAFRAhoAj28RQsjexyP8mpX577fHdY
0j+WkIZ6NdQoKkbvG/L20spWG/CE3QgSCCnDXPf/wHVCUIOouEbMwMWHa8lgVRuzs3MebK/0gG9E
w/xggzcZyhLhpvzsDAmQ0NiB/4u81z/ner1GaLFNlWwCn7FeeZEjDD+WUPPUwoyLzXteamCn1mUz
6cNfVWyQIFXtRnGsVoSFy/uLfPbgc7ud59JmncUrBlCpwmkYoIvvWNTzSiH3uF77Seat335PT0Y7
WdFyuDDAbu2Dm57KWIBQAo7kKwLFReChn1b4rReE2s9pwQteeYykJs3j+Hdi5GM0u/WEAxh3PzO/
ptdI3547dagt4YxMr+UGuzwJzDht+eLebHiJjFNHyN7ewtQCnVJwLtRlru+Un9YD3zPdSZyqIyA7
IJuPm/1SlrLhTJxQEaJ/+TgwfMR9jMIHiXT2zyiGiJPVmJnDO26DUQUlxl/brqONzI12Wf5Ln2PB
wJso2bWsua+/+2nFqO/N8kLrCcphg3f39V3jmUGGEkBOcNl3ai1imdWWC77CcrrX1IcTOMCi03P7
culflszDjqtEyfJ4kcJLyi9DtAnwjDm1mdgZUW9ycZp6cWZc6i7k4UU0+7cEDMXXXAQPZidwQO2s
dJRhjRlVqJo9YB7TUFCGpZ0J7DYOBiDtiLpSPmmkoAS63/VNBMfccE4kuyUeIAKihZqjrC4hZllF
xpsOtKBWRwWpPAkDluW/+q/tdl+Q/ceONZ4+9KOhwLy3AAqiJztVFg5ETw/QBZ+n8TvY4S9xcx2C
+09WMe0SeiZx37Y+HQ0xvj2KMfZix9YuXi7e6Kov3wo3QNhECMzR/BewwKO9yrDQzf8QAShXqpSX
RJYgMlLXIcFauS6gGDY8h55FQujqyGJLJ/jG7JWOR8y9jd+DNQ7ja2myODTzEOw7j94jlg1GyeMa
CPu1cwCKtmfEIbY6ZsPT9Huc3/Uy5za9Wv4IDKeRwJwe789kjmitfUquKhTDNLp0IP0zrVI961rj
RRW1o6BWT+ppvlDH0uFTMigyILLZwin0vVLcuA2Jovmj4WWC8TfoToWRTKsebjfNEDsWNQsRJm5E
9B4AMKBp9m4xB9IIX6I3vFRVPyWGE3gIonLh/GWV2tb0T0Dm726TFEv32DGvUsxlol0WgKHiT9cw
evYOxVNFJC7/vCOp1b3IYZf9a2QIYaMUGsBJlqDgbYvEQ0DGYjdnX5weJBcqXWjM8w9GP5Nf5fij
XBsMnhpfLbjrBl+P0Y1z96btIVnyYG8GJzp94A9I0bEMXtnYDz22eIDpjPsfy0NZ67eVbQMLiCYn
0Wlv58iL82yNZ1XKQCoNQr4e78icMQ/XAbmrh7xS4eqplqWDhA5Ef5S4QDB+yT1bZoNceZIYegUm
m/e8IxytmyyQHPzWc+m3h4QWR6LcAfwsnqGO6CTrVUJJ9RhgJNSN3eLJBHniFmRefuVmqoGo7/z8
rWqRxr1JuG3jRmpH6a+OcFnvgFK19VuqI4fJfU4Wnx03K0AY91x5IFace2t12WMEveYAlWzgDlf3
12OXsmzmxQuBWDpJdOmZ8+e0N2xmGaYLCMy3+eXRSnYw4tAizB3Hxx4Z+p5opJsKLJo1Ajen+R7/
mU37nKK8XHm1SaHDSW2d81tdWFW3lK6SszkiSmP9nk3UCC8X9rWnNRI0FmV0DvXPvhsDNaqsP1T9
SU8FYqwUr9gqXROSvrr5qs0bgNpL+76DDvxt8LzzHgBQV8I0hQ1tIoVvh+oqCmN56ltIiRaJBtsJ
OY3kH7J8JdLtgi34UOwuXpT3Lkt6S9gBjTGb6gefFESqaKma1KemNApG51CRh1qbp0EAchMUvHDr
DtYD2PIwBEE/8TGJoMgUHY+X0RFNmIA+uKiIJ7TtjLB6ckY4e36iBPzeJcplmoP7raE1DM4krie9
Nkp5wiHLsuY2YpAaBq+VQOFfy5+k2mvOEvRp5qK1u0enfwfzxe0MbIbjtw6LftewMF7RQQ2suCt5
IhEQQrlMGLEyTMe9TAVHpThfVBGcjAp+CW71ymSyCV3jII78JbITcC7HG8GxzaAhO5jYg11I9f2i
5lpRAz0vTPuKx/GD7mmpdcS8O+czSn+FNxiMEmIKRDhmX/b0siCShS5AMQeiC8ximZ3/wI8/buAb
qOIU71C+xJ4ODf25A+e6GPAZqs5puaGKhtBeCIneYpjIZh8jjwXAOtqni0FShe4Z2Mdt+LtSRFNJ
B/su6muJq+fFD8MSwrSppEOQC9mqKZp3+Yte0Ro0XqxZcaT9XXzk+NwFD0QI2iAHCRTs39Q649T1
g4PiL2GbVtx/wtC+caH1Z2s2JCgxZWc4nLGbjQ/GdjJ9iUvYAJUmhAwYyywcSgvnESBzKLjkpPcC
t2tD6ARCwFfJXZu5r4jLlYPMp5zXB0EG6F5UrIHFxzwBtLJ8ZITOOKZy5dmDMJImqH834wf0iRXY
WCmM+SiPjD1iPhxXCQC+azgc0tOVSdvjMinE17o2yJZdl4jbbX9SquPHXkG17DhVwQgDf6y5TKju
Z76OVc13jHNHpZpyk1F9cCFPCADJClhwRzbjZKZ05WxrlXohpnQf0XjdSVJ2dTGeOkajKrJCSGGj
Up+RviayErFhtclGv+L0Ez1WE0Pw/LRroCeIkuQ5FYvTP2NmwixtFLiBCjDdFn7sNOFVGYLKD+fE
gf749JZqLi8KTs5Qw9SOxu38OE+oGM4P4YEpmDckm1fu6GA8ttzTA9uVeHiBYmrV3yrtmXPe2pZU
3k4d0Ss+fvLvV62s8O6RL2hVEujjt+swN9brlKshJe9GYPBjVmhXCKv8otknJ7520dsIXjvqV+39
4gej/qCD3e6vQosjP+mocYt6iSunII4ynVOQ4g95w5nb+T/ESh7GT8SxVToDVzJp+hO7x+xzXZmR
uX9d/JrTGQhbDUvt7qHvL3fYbLPWvV8gfWPQJf00BQwdYLXEugXEMfG/wwTCBjjbdHibSuCTdamd
BqoV+L5Ma45FH8B6MBkgukxhiV9wtPHEKLTxlYwR5pFSYCTujrmWNcd/zb6JCmFXaKUkgi+ClDak
opbVT5EwAzKjdH31Lte5T6V//cKMWUmW7MWKLte+8HM5zgDK8L6QqHmlkjU76omPoaz25NI/X6uU
iPXzJ8vwtmJw8UVRs5AA6RSVxBpIRUW13ULhvVeXq4cqWFnb8WJbO9xTK7IfD1bvMCjJTAuZb/z6
Jy3yCa+UD1/e+ZWEBPLthGwPcnpl1lKkzYwWqmqS8RngdWMbwPquNSXWb/Di2ODcvk9efjfXg61n
6aXj5EIiFqFao1Yq0m95DPZD+urlT1SpNgp0HP/WIpbbIqp0FASedQrhZ8Rvpuus7O+/RCSAqZUo
jtZWoEIfN3KHXG93sfSOCW8xxfmftxJZWXrUR8nUR/RliWCAvp1gryTIN3x370kgeBcfHyS58x13
zxej1hBPVhFduNpUIuFU07g7HumSJbBBn9+hA2EIgNesCbs7uh22sRuvjuqgh6aMsmXW1PfeGcaa
CT5ld9+grgDlH8pU4pZV5LeU7qxbNDky2mK5ngy4wQMnaAghLqOlyHb3CajJMJo9VPc2m5uQd2L0
FRLtcaZFODaSzdclBlznYBcktE0Jn7Awe3wnqWI3K1JZe/d3bx4b5IjTsw5mhIDY9/3LqTJ/FZwS
juZKrMFj0jpcQgEgIzgVpaSoI/xkmzi804XyOnTHqQXBvlnC+/Bkb3lnRnOObjRzgGAPuOjB+CLo
uhrhmw39DdegHXEzKbKWyOlCJgFOpQgYddYT7M0OpA4CQwSI1q7CQgX3GcW/Pm1SXDWVphAjUzzS
IeNwJGNorwG1yzTMn6SeOsh3TqMXLuD7ew4RUvuBT9I9fKWt5rkjkHq/NTmK6dYXVxrtAtyiQeFs
4gzvrYt8HI9/2dyogemu6VGg9UDI/RpFQH5r5az3ksQRwr/faO+SpFfNWvsA324tm3S8W1wBgzxf
tCN+QjgbPvPdNJLUWyhxpo2V0aU2MDxdJ5SiNlIdmniBTJ0gIernZOjJDJ8H4kH67P5azd3X3k1E
QgzuIdqkG0s/Q7Dye+XbhBkZCQ19DIISu63yGAASzMCsAzxA0iDx9VVWr4xSrTHsnBwICGHJTpLF
LqGVzHn3E1mXTBHmQeFnVcYmBsUt4d3uqOHUXm4Kza1Ph1XpOzBKUSwFLOVsIxLGq5jIiWA/mNYh
EDKxu3p/6/2r7ZctxQzTG5vTqnFQu1zVMhNLBEiBwR3/bkszG5Bso8EZdzKXH1nO4lJiw1/akm01
TosiFpIw/PETvI63FfxNkbv3kFlSHXZ5vyATqTWw5qbTMmPCJFVBmuKCAP57SXiehGk30ZIbvj57
HNrOCSbXwKZH8a8Ido/beVmYtl0kqmfCJu/bNl7W9QUPgVSuzxM2zlQ4F9ySC3Z5vZLeCDv9cZB/
sok73LaMrpfPBl9gTDuS+r2FJQjyqe1vwO0gwAlgUgSJxtssWydB1ZaW4M215QZGdoggKiqRjIe7
CKGL7L+3s16QhjMP1gOsurVZMDrK4iu3+RJFEyyH5dqhwoIIVye5C2VIKLfb8T+xeNQnt1w7hEym
lJvV0kuqB4k6LVJhe8X6cs7Lt/HsBZbO3mVUlIQBazWH1OqmwxK/WjF+lO+Tc7+25+uQAK6BF+e/
/3B1gRZsdVvDFTVivsRqSg9cwDubXzE1Qj5tVC5lB3TEn5NSfCwpk2SQ6UYoDBTdckmVI8woUhSj
+8ehmOXpaxIe9LcWUpYli0G0yWn7O2WtMPe2rNOHkRae5kMF6rs2qkgesTl733sVUNBDCP8Io7/3
nR5Tkra+NpgaSHyXaTovUI9FXQDTYiqVwyKl8qiGuqmQmpGODr7TZBY25SBN2o2mzXoWhMiRo4bu
hOBQN2l1BnXNioAK64AzE4icOdN94svPtmy+IV6kq1ue2Hr8NkzBuy0humQ7xlYOvK5QoL1mlCSG
DhVy2hin+x7UjM5Paz638jIC6Vqi1ws+agZPGUxnGLA/d5XVOTsPkWmjj39ZcyHYUbqtYit+khqi
y28mfOoCiMggfhIV0RyQiDlELrmlJqR93FNL6Xd5WGDz2B7IDp+PPHrVS24i3RfPSXG7jFaT08J1
K1qMD8FQyq+6hLpxbjb4WhgD68zD899wDTmT1itBrkIDijmRpq72R+jOZik6jzsNjbqZPjB+UusE
aWLvfTQZR+L2/FEAfBUXzoCNXuTVFY3LruF880ZuNSoCmcaWbFB2TgVxZLESZI7GiNi6DybU7BD2
YQE/mrkdwf0FvyvC/P42GbQ8k6aPtsGxqAc7MSd00c7aCEvcj7v9JrPz1bLqOjtiQlDNv1gWeD0G
MeHmMuVGz1q8soWYp1kvSZjQG9HqI3ph7/zQhezHLslXvbr2XZKprX2VM/tiBzsjwCGloh6o1etc
bnFzktIxkv2MjN/Uu0I7XPqlBVEfaQl9T+OxrhULqrrYxRvfb8MlxdgIUreovvqm1EDIGidCg37L
HwJhMOKtkG5r1JPfIfjmEqI7XWEKlGJSe3n9VJltFzRs6woyRURZVxrVuULNuWtCPvWV6X6LPdSS
+0we9sdMej7hzIT4d08u4onh/TNF2o93E3k9pUrFN3/OLvuJ1QGfqKZQGBusnUW8vtiezXwfHXaS
alqwSuA5aYY9sUBtjbHuOOv7LD2SOcT841YVMEkBVdIWYi1Ei28wCKssiev8dFkdCtzFVJXeGfCe
sXjo3tSHHiVad0vjS/s7AB85GgZwrsJeXlyWUzEmtVAjVJPCvT8yaCpHQPPebQK8M7G6bAcPjnYi
HF9+yeoV8sN/aVhi11spDPYcbHL7amToGMaANou9n7JOXqEuJUVFhlpJD1QuzyG9vl4PYzN5JRyO
ZyGBO8E4iR+7187Yd9VF8DvvuHKsrxAqASZm+Q4HzIXaPkU2BV0gPsFj1VE7oE2yOA4g8vtGS4dy
lv0JYSRZUVPBgS0x79egqDjXiXx7zxePWl4zVtxH/yiQndyaSwyKE0PJcIlsgX6XAVHzpgpsPetB
lyKkMscbWqjAZDBFRCBHVIzlzFNvw+GZvwnyZlV3nhLb5Qz41QAx/DpyXJa7POYPPA15quBwgFdh
OwStyQws04clWxIDc1qnusVqYge8vgxEZwSOXI4d1Ur2/8d3CT9ov0ukJH1BoPVJcw3usTI1+GsH
+iZbRhvruvbXEKZidGcexQbDtJYoL/+opNGufN2UZPe+YY4n5h+dzM+QsGkE9BV/HZP02MpI0+s5
dpAaEwpVo8GmXbgTDbc5vPaGJZW4WYuuEahKzNw/wcoNvDjZQotbNwxg6DeG7ClzmYvOzGvBRNWw
9jKs3tArdwkGvhcqEBSvJqc4rtpUZrdaznlTOM9JzM+PMQ2NzevkoSVy9aCreZJ+4OjcZEnX6Y7f
+/LsnicMHQYDC799yRAnvxd4tvqILGEeqXKtAAieCNdc3GgAW+5BMrLq9ARAxscUw9VXvbvzcjoM
hUoRftRHz+NhA70DC1R2GQTOttV/HSfrJdtubyl5YIMP02Gj6H+YZj4MJH5v6OFJr2EQGoDfqaNW
ggwCQ5JKdq7QDWFT7L01+uH4OZnYh87wKVYFx/MX8NJ2g+aypppslWESfweVcQkLKtuv24xlgXR4
4X5yfzfgN+j7gIgiOUwFOdvc/mZbZkdZjEBP9dpWHo+88EoOeCRxzaEvYJedLXgL5EsqcHhLGtRt
P6j1uPdIiFs7WjNY/x+L5IRc8HPSGaTxjVIm4vvPl13fcjS2nmiw0erVNwWRUHIGvkzuMuX5jVj4
l11spF0XjvwRCBXOQw1ntvKcpej1Fy/d4W8K8RUhIFQly41R0l1TKtYe3pHHjUklqos+09Pz+Fhn
FIRDyEMITmsQhlTpJvo2nN8/5p0VnSY9uLqXBWuWDF2ZDRZ/TEIg3GuG3jhAmNGZz1ZDMOZ76Rml
OnC93tT38SzTgEIuHKeJBxJyNf91wTOUJggRLi8GzEPLqSx33W3WVc0X3FMJaVprdHwEzxchZVmJ
3UoaAtSsL+9tszdycsN0HMhNJ3+SnP3BoD1M7ROwuBKa3Y/Ele8ZM7U9iP1gFYnRWM5ILgGCemX+
PZBVRomrMpyHK56FeIFT5eetCK0S2pqGYEIWtlpjA/ZVhTZ6OwtdKcopuGaqbjM8wIccsjQvXELQ
rcPp9iZW+H3Jq+I7e47ccArPjltJNT0QNuffq27eWc/qDjjsDCasqnXgjUO3y65aSbBGHnYonu4B
xp3q1B9E1Nuf2Sw3hoHRp9QSovex948ZlL5NRnWPFrhOHRqCH+ydzR4ASLl3B/yfhxXJQ1xXUVz8
YGP5nHuAr8tFlkO1+sNGFEU81IZ8bd8rxZgT6loZvntfy3YnEa33fhCyx/s/g5bFvV+FN11AFpGn
b6JX8T0Eub0p0U7FOuMEWgAWoUIbYA6kIWff50VK4AQ9JQgsdvkVBZ+haMJGM45tJiwDw88cOLuO
pNqE05RuMlz+1EuYytSKUxdGtEgOaAuMO/heR757MzbE8K48nliOW1IJrX3n2PX2SZCAJp4cByHB
HyoMpgTroAf4pskckSS6pXA6qT+tTw/vMXN4xvdF9vnePshEwiUTaITKuxE92vVR3kL+q/Yncvov
t/QqSJiWeHqE++apmuxcKxj+ijG0PUjooZGAqD6CIMRR0W8fIqE/kZv9EPWbkzDYuJ3r6IR6HTH0
3knvV1wOJv1BlBMMkvDbYPblod6FJQ5ci8PiIFY4y9A2N5fEJdUnML+WEcRScrVx9ZEpC9DtUOKV
IMuPQM/EkmUeffrWnd87+9PSmBNhAj2R3sQ6OY6IMwSr3trPre4QIb7MXClYqGXnBclnO8TEG+d1
Rnqc5Iyt7IsHSUWX2UCzGkutmbSKjypVyDPdita3z3Lf1Q9OyOwZdPmVtuUSOt/xOhjF70vYNgX8
jeH0BtPcbHn2piE9Sk2j53TuK4IxXrquC+oO8wMcm/johzEULx3B9tILWYYGTYumu/k5rJwaXnTb
5fIGVKNVpkf9E3sqwap+Wtw4gvIX+7jq6fo0xaL3PoCovdWEDGxFg0zVzxyV70Yd80nnFAYJnBfM
es0acJFNeFIiLBKUh0zksRytO2ZGDPAWPKhzlDHf7GpS3+KMyU5E0xa3sbSE1uuTmrMsjh5GPSPX
LJvan/0agDh/FY9U6/pTwbCZ06oh7HBiIPTtxuQXPeKTD4BpKAgk+jSoz6AMvAdQCgw+hzz4+PmI
9t3hil1jHIrhVzDJqajTs0f4y9yodg7zUwU9ocBRTMvwl5VvObT6Toh2xUdVj7RHwQHyJM06nYWA
ARficdxfe/smwzT1Vguah7nPRT1hAfKVwNfb7sm3JatA0mMyN1gwTKkHBsreznqP05hVYgBk5+AI
LFg6DEyNBOdIFo2ZQ2UHBlK9h2nS8qcM7h3QBWQh/VbkfgO70vEs0urHBVRZLne1e90ISMOBPDjh
JOFaVZnW1yr3PrAreiheO3l8Cnv9JPTjqOVeZ0rj8F7S4LLU3DuZS7Y4EcuAEKPA/KHEfKPyYwMF
sBi/Iy6OZhDtbl85kcmUUcnmOVKJbVXKDaBaz+uwaL78nSavwzqfsgWi1FQH1He4N3BQW6QLDB/H
apbXHQR3JjETaZ8ZObn5TamIA3mml0TBvHosY1Ler7Xlcg9xqrwbqktvywOVS3VyjAim3PRIsPgd
1TXTyo7n5fYVxtmFrvd1z4w3zSF0ExvJr49i8ijtrOsLJOGwb4ThA8zItAXCWuTk1QSH7EaVkK+K
G0xUo6EVYF7r/nBUEen46q+XBubR4qF1Ml8ary8dMYpGzAYPZzAmHT8gAknVA3O7eOvfcJh4WAAY
w7sJLlxc0ctHmkxFvXenP6emGIpQrdVh+L/SpLb2hLTkTEi+q+HanFZWXjZeLFEhAWCNDGTZFdZX
al1M1gUz7ljQIzluG3cssHjiVJqY9xtumZb3x1a6K/35nUCDo24/fdZEeO/gU/w4S+eNqICjlWof
Xq+qUjcdJV9uuo9SGwN8e2HODagsXLP5e0F4Bm3A2ZbRU1a+ACS9ceE/HyxKBAnn6gBIk105wfUl
mDlVeYSK85rQ5YzjTqEnHnjgO3Nt68Vp1OiJCL5Y9XjlpwaA6MIBPavyIQLZ/PWMs4laEcyoBhrj
Isb/VCbF4LeSXa4GM2eXNJXUDKEJeZTNVI2wVFsvFh0CHl0MFoqWZgCj6n3I7+XhiszX7+mDYuKX
BR6uaea24XDPmLu5079Vz0x6cjocROnlQcZsg3+bPmNjDGw4Bt6HzYJ3ACcHB5dgc3JCNYVAIwwp
rRuESctMVsp5fEECEYcJ0vCOFnzigH5DhI/CJECZXZ+PLL9cPmUCozt+WtCUEJTgtPUWjUSjtE2u
J22HY9ljDNsbOPqGmlHhVEFcYAS5ULPRV9aVn9K33hCXaW7TFF6Cja1Z/Xf+KFKdAvHhx/nyF4UX
9ZLUXe0WtC8KCuuNgdOLQcf2Lx3UzHPfN4B+VqN37mhng3MlFAuGqD9n+qLM6wxcYhsyIK/+xqut
3BP5SJW5/X0fnt+yFnBpMTXjgqOVehb1M2k/ez0U9ZepJpD88SnymyxuKwGNaATdMLE80oe+TfgE
HnbiRyHGgf5pQBVdpO9eb1hsur+i0MlmuB7Cuan3ngpyuUq0sDVo5yczzV72QYjU0udcHYGzCP7J
5o8v3bB327T+HmhEexszubnZh7p6GJnZ71UKT2qgt2N/zvijPwxYKWQKNXtCsnFxZWWzqbqMCgjU
mHAFKYyCw1uWPXaLXF50LlRsl7ynHJoAbPy11js8ROmAnJzaO2J/IsycFI7J9xd64U+lROpAwz1N
dHdXU3mjwOh/SfOi6cmC7NuZkNezeHHHlXoRwyvcgWjulRvB2I6v6e62Zt7sf7auQ8lyKw8VA71C
xUGBznYDUH+0LV/+Mz0QdG7UrWV+XdfLf7bu2zUdgbCtWsQMhH/Im1FlABQA1isdA9p7cgw/hoI6
/Zr5tZ7qAV99wM4Q5/dfLSy8KpQkRMbCv2hF0IC7NBDSwvo4qfHa0cd41Suy7v6ukuesPg7WeWzY
qG7f18/Svd7MWratedzp+BRX1AqFlwKNN0KON/m/VK1OQd6vXMNHnEyQW74t3DenzN1A0UZ4EfgM
3Ie1ZpmWQLcIQ5F82uByS2P7eVH2lcnWd3ZvnykduETC4aTX3QrTZLkY4ea3fPbIqiHR+URVLxVH
qznavqXzmSKzIWnUiSfJ7P625sh0Sow5/6tTpmwTfh59+oYksfUHlNReqQPZRBBLI1OwlSWaj4m1
rAdIbmLmLrocs+cGVKwUxOWbvY8p/H2FUkjh4XNqt8b1uKGT6wcmPJnTKWrLF/FVPejWRLw5GTEZ
kCYSrj5fw0d9a9jyMenTVUHiTvhxLmg/cK+aM4aEGdUFRil22bzpEp3IikHLBQrklPT8SvmdxJFO
LSc4NlkHHk0WyRfrOFtNH06oyW4/K9fkxE8WYJWctXrtEkL0e9+MqlrQ3cEV7YEpsaInh17NNgFN
YCCYtah4YnJXMLazQ+kdPo9tzV2fEQKiGbrFpMqn/is3VLNqH8MFx1y7xUITKDiiQmmMXaZjHYuB
TPHjLN6uvaFJuppwHUcHPqFgFDVPTPEhZBUF9zRuUxCgBJLfNxHzYbXe5U3BUHZoGIHZIXd6PkN6
CoKmOi9tOpA3c59MPfRB+RZfaOhtdgwLnmJiAX6N9g+hqDosHqmIbYw9Vc47IGrbT8cK6MZ/DAYh
nFfe7v3oEwc3Yp6Cy0UPWrZhdgF/xk+MeS+pTV8lIl+iYyD6QwoA5xywBVxFi/1U+9AN3bYTtvrK
y6FO76GaPSMJbk5+CDra1naibVSkWN4l6OPDgzQMTR1JQkdRbrniyrasxrGBhnJPeTNWCyjmEzA3
CryuQzppek/dwxQQEoF6SZ0EVkHYWS2gWW1drcwEHFLzR1Y1GUIutGtb5gfCtcbtDVSTDCfIy1J/
cwLvtoMxQfrhvnQQyDM433ssr2CLsmyx8SB1LPB9w6+25JbufdvY4VEP8zCPAaCrPKCFs5aVNmEi
n12wRoMgim7hSgYtJGV/W4aBVjrEZv000bcSyEmuYJpeD6aqCM/8/kmjkp2vXUDYMrKqvWX/DcEM
47iR84fFhG+l7ynwIPjdKZ+2l+4Ms/vkPei6dQXkspMzQP18UgL5nKXnj9/b4dIkN8e6tIbJ7H8y
N99MQH0Fa1BeZU/gSz54OwpABNKmyRUBlsu1bthoMf0sMXwG5BDigeclh4dO/kXT77fvIuDAQ2Ja
CuvdPnMsUunxMtti2xG4/zmiZvYJEBqf1RJKnvS755ogJuBY77OKaVntS1y2j4MSnka8bA46tXNY
doIQwOqI/xHCZpbNu5zSxlikcA70gY1z/MzWAUELtQQMebroDPRckbzhnSz36fF3rH3SNULhvDzd
qm22O5szMPu3hjlLJeENUvZp8j0UCzxCRGFdQhcyn+EXUhzqJedEZRGJBEJH5R50lKKU8PjDvIrl
QWR4R7mA1f5XTBwC8ShsaU3hFb8gvYzm/CcE41sJ2rG72NW6LNb24jcvpIY6yCVQSr5W3XVlUOE1
Ot0o05XMqivIjPcwt4cQ5aGv6jSs7aHdmUfhj7fhSZvEFE01/9laK6BdqZiLnmjLF4fwQVxjbnZC
NgGU8XIeoUSnGwmb/TlUFPBV0KrTb7LtioIvnWSL/llFKLmWDVl6zoBVMVPMayFOtJKzsUCfu6hQ
inMc8TmdMlSu6zwmQgEorWpelGiWyFEw69Y+MeNfq8qSp+9sJ1mUIYY2LIudZT/NskK5mk0GEvHI
YLjTXbuF+m8KB0vRpQ0BYvm8pO7wLlOBfjlnqraTqJDuXKW02txQcWP+fl8cPMIdy9qMhwukFm+a
A6d46naS1Niego+vzh2Xhy7iTeb6LF9/KLQuC59LAh3DbCZge2Xm40qCyFiB/GksrlEA2GBulpwI
+zxJWqxyiC9wkIOG9TlXqiVrJ+nmBxjZw6ZBYDTZeogTM3Aq2427zKjm0pAb5AlSdEDSJ0tUGgV6
5IF6kOBkhLg80JwCR+QlMJ1MwGDVqQ6BUvUJB+OEyvtaklXmU0FISImkpOAPplV5IESI2WIimVJv
4MEWyeANnGDBm0dmQsgwzu+ax6eQ58Jiim3M2aVZFZk4GrkGykQRf9SQj5lDqAO0K1+RBoDGHNdP
1GSmRcrWbMqiNgUqkJH5Sjzcky+vZUXAwB4whFmFaRbo8Hn5Wp0iQioWatFh0jqsai2Xkm9HjkqM
4OukP+dmvUke0iistHqW9pLR70PBiSviPxC5QoedCp8pAlaBJ6c8IZefOF2TiSuA7yNp3IAcLCxK
3pd22MV26JkFtkRqUtIWl1mbWQpeycADIEIMSUjcFeDSrzMSjcpT5GNV/ygxPp4M/d7WWTLpw7T1
um3owMMsaTrxuceAHWLFyuHgqxaaCk1GeXQ6ragoA4uJWyk9pBNzVBg+9biLZmfAOZQ8QnFk1VFw
OfkGa4AkC5wi5tUxEuNNg3AXoEyk3ALgVUK5FAOErPtaATosFec0UgvSai0cwfbYv5mm3/ls50+6
9ijpbAOdhmxNIoOgBEaIcU92y2C/XoGQ1BU94QGBeG0Ioy4M7I0Wpw7cd6Ba7q3itmlMWx922EVa
Jw6IL+s/SRjm5IHH5XkVrGYV6IJZEP/rWcPogVtZLLz8JYCNLGxythFnTn/RfKuwwXpzKjmcqpgG
/wemqXzWVnlN22qA1MJTqRq52w5RMw6SoSZZQBb0XkYdTwM3iU3NjgQ4U3Pa924IofS4rGNs2mIJ
6r1FraN8alFVxhQCAFVJHK8v1v6FEsp8+4xQmheHAews6p9laaz7r6zz0s7dleWjK/97ufctTgHh
79MlXlLjTzHB7kAwmovSufgdGN+N93p8JLp/k9t+rsQWtZk2Q488ajKBNqzf62+MZ1Wu5A6gFoK6
jippPtP3MIp5kZX5NCCAvLaQZ/FzXCNv+5+5vxQfRWFdQjw4DYQrM0TdOKYojr93unc+tCr4aneK
nTe0HZJclcQ3zjOTvwVB94jqbdQid7lPvC/Dxb9FH4ZGzDH0hXL8Ndb3HqF4ags5t6oNcu2BFv9K
YB84RKmKKwrL3kQ8lThix+xXsaZAGhsk15s5cYyhiIJRjbScgsG7B8H8ddISpLcl5eObQD3F0ZkK
JA5HJAjqffka9xV1C3jwoQ2kjiLTw3NPXZ3ZVETI52k5R46fk3GtZv50qfcRtWvMv//ualXUJhuO
1igezDBwCsBGWJMZBcKgsAFaizLNxmGZ8hT0ZJydPflIC22UWeqhbRv8H3YqjP8/v8Pf6Z6zgOAr
4ui5gVC87KXkIQmUdZtV8wBnQL9oVj724A6kmOu2roEQ5vo/RYKphHwUgUP7erlvX4s7jKn55OBZ
av5GWiQEugde9+0DsBwQMHTNCzpOHZ3FTqSkOnHo06oUEuUW0OiTr2HTz7qE/TGSkGIY/ITcHdvF
3BRqnnx13T0YtKaWLY4ESYN0/+UY7jHUB5ghxPy8ExMt74evwqMh5Hc4QWcph/m8dtYnJmyktKSt
0J/zevL/5xKrgP8TLnqWHlOIGqeh+ME3c6dYwY+WzaiDa2EfQQrnF3YiOir6nLo+qh69Sw1JFG0r
jgMfOY0j1OBHmevOILggANw3bqAz/fBdMg6V5aoMnYkDAM/vrqY4S5pzex2fPvQzsBWnufFzZC2x
ATlZzAZdCSm4o4pwTntf8kaN6yKkTdfvvptmYQo4aCxEdAv3kTD68I6wnLvqaUMO/1gkWKGvlkN8
yLthg/8kGv2e1ZLXuMFFrW7Bz2lK501/zFN0tdBxnWHX8myYwaktnHYbdtLKjWo1rUMT7TCDSlPn
2PTA0DS7LqKiGYjHYjikMmjGEE7Urv6FK73TcTE2T492x/YJSP+Jez8qKQxagdm/YQwJ8+Es/bsL
eBwBjYoS5kcUJ7u76hS8ygBPz9f3em2+2VYjVg0tNbdzUY3DqA9CmIuGWYsV2GHXAssjhVD0rT4f
pYV7QgkHxLNDtG/p9wn/VmrUP0VajlKX+BUIqwfvDtalwwsmwUPUrqXF2rx02+pCmjICO34WyMO7
gNdo8fnW7VaPHmz0H8whjd6I+cCP8dtHaJBustv5tjX4m3Wvscswn6oI5gA+6+rML+DbWxvyctpr
nAN9pPlt8+t2KelgK6/3VMusbbbzrFyx9Tw8dpmf680Ou2RKhN+R5GrBditztkdOuovHvzUAyTki
7pC61g38qmnsnN6ur+RpkD1mB8odB+7Q0BbfMDCp1OxHar5m11BvVYL0oJcAutxLsv8GeFJOWFCF
5ffCuO9L+1atSD6mRPCk8Eb8AT5PiQ+9y4wkpckiQ5rtfFhvHEjLK/WAO6qcvH/VsDIPiY051kl8
r6VuiYOLii6R+BShxXezebHWngB6GTAxX1zBHh+9/s4SrQ4hbXdpyEAwZrWjOim0b+w/dqy1ZVrn
dnGjo0FQ9E2NluVlwnfPbNFm6x5HuVgYqdWLuUCs2lzyOZgj/G9FH9kRvxpVmMdsbH/ZmVNsx63i
rtm0LfSrWbs9+/HVwUhF9wJRtC7ZvuNocBtpYtAfASjQzl1oVpuehOziRMQqAuM/vfEn763ze7WJ
x5o6CcWwzhsOrkvdCimlyyOIPrXxJ31/hP4cj2788rGtX9/sXBx8VhN+BcAarcO2rxk5pD60VMdm
aDl/w2IeQE2orZseglwzoDmorZCp5uxlId1c+cf0YjQc07I0O6RBOVSyf1ZN2TE2jMORlPVpiPdr
xLNS/0F+IVpZHkT1hudAGTV98gM8BcpvjB3xe/lTecBp42EUSWaP++1SL8hBgWLYfBPyHColUwuq
RNGPQ0DAzUYPS8La6GepyTZponYW0fBoGnoURe2L47MKP1X2xNGEugVAQOwS6I0gDGbPrjOuuhGJ
Jchh5LvTb1HvDmSWhInRjawubZXngy+wqecwZidjV7acCRZyFV9n+RooK70AKqDwxRWK5TAxwoNM
cmqndkGRqr0s6OsuiyqQYrqIASlrXpDzHsBlqBtYhxICAPtCjlhIqdbRLXDj4E+smT+AUa88XTK5
9V2lS0Ft0pJzy0SuKDB3LkTMUUW5wY5tjBUzUA5ztXxPfcevD/SR36VAJZOzIE1p9hB2j8lqr4DD
OTBjm+Sq71deTqx7UdmjupnwN3bR0Egf4Aj+RsWkiFUz9dHVC8uJILDjVFwfWd8DCV8U0gQOqhW4
cyjHTajyUseJREVo2Zi7WTv77FNbBFmgo9rv0xmkKjeO1snMurnUBr/RAT0dUaoX8FH1epynxt6z
XFG/JhFbYyq3WmAznxqEox7UCER6o/WjqLo4dfiAsBUBB0wupwBtQESR9+DsnE2RZDM1h9IMmgHV
4HZDqMRzTMUFUHHr8qEKze4YqLdbDJIif8NoZo5YbsPYgs/Tarn3MmN8kEO5SFQaEPSj9NTCI0nj
pHYu+Udg3aJHjWEUExpSdou4F6+48de0GmNRvthdToI6m1gBkCail+ScKeTNmj+lM4SR3RyreyH7
ltnQY+0SFA8+L/K6ttPHQ9rOKHZ8+7IyG5tXrjWRBuS8mByxjJ/zsd2o1ScR80B0Fn3mRA4W45pG
mMArosKc4EY8RIgT1GJ+zNTrg81852qBgJUyZtNwh4eE8qgHkaqyYAzkdC/zx/Q0SVqHhh5aENrs
Yz0ifIF32FdzAdrcwfHUkRRennyaB7MKburOvVwXuPEbJNbNvlOzfqWFa/2GCT+0od1rIV+M96U7
IscH/kxPB/GslbiZLP06ATOZp9CP28GCqz8J54YPIXHRiIqyWNdm+cmQ71HiqWapgGqNSn0doSNu
irMxckxq38abK25aRqyT5V0v5nNHBcmYG9vHWHoZLy4XYB4zBgq7QJxyxqttqzEjZNIKMvS2Melg
50gn8+QIgknpmNcKGdka4IfLTrEob4bMnSLwu1w2C0NMaDvg3dkwvHCHavuCYPu1XA4QJluTz4BC
Ve8caKVo8vmBMxEFPumBDhwAl3Thz6h8KTInmgCwblIqbfCzdNu0BoYI5FicolnBc6KFbvPOJMKv
MfGBicBJ+vO8H6v4LSQgNTNJs4VE2v9yd7zRuG+/c+8N6+qnuiSwAorkS1SieG17m51rC7jOTbgl
Q0OAMBrzNH0isqNEF/46PP8V+6ICVrozibYF7BrgfCCDpC9bH6toPI3DyEm7hf2F/Zc1NaKqnEZM
KcgJCd40Cm9pErP+YiUfKFjGauGn7Sdxq3hBxeJ7zm+u2ySBs9H5jHMxloAVKh0qQqiZoR9I9rM8
PCQXAHIlC1PRMUTPkY9rph2CNoDkt6xmaCHISNyumcswc2Un1CQpUmNDhn2JpBK9CKNJr+RJZEOi
ZT8BZ7vLKrx4pyPPutdvamMQtu//1FC6VZjjJTWZJdmL0Psxgjp+NxiKw+zI9/8eIFDr6eelnDl4
TvZJFSVeFnUqecDTz0cReup9y9MQrF7DBnt7NB2FtPzny5tOHm8u/X4MwRYaycs6z7cxiuDfGyOs
PFfr+xXAX6pieE4Z11g7mg8PUw3993211Q++nLjJNu2c426yUATE0vQJmMGR1Eo0vnYvd06FaVVN
YqQ/yPSKRf2GUaIAQZCOtip3Z/0m6vQ+thukzKD+nJqqV0rL/6hqHioHj4KfXpOQHW6XuqmYXkc8
mYtGzGcSHs30ndlTjLCcKtVU/q4QQZ8kR7brVdAhPlo1xUDRwZzyZLNHYfGigESrm7QGSO7uGL3y
gUzS2jw4I6JNLvsYvXtICYWrR6oct2YnZDI3Pq1T0RW85hL0xaW4YQlqJvhYTZBWSXA4UR+4Njiy
vqgjn7arupNadQzNglSPVS+Wo0eDWi5Qwc62irewMfFoGdQ0jPMvagTPHM/gJlmAyXQwgMEmIUPQ
dwBFQvb2wyGRnB33u81mdpdfG2T7FC5qpj2wk84HV2Ed1/yEmf0u5i83FypgYDhR3OSKfL7RpAQ5
mqbLKrslxeUEcg6oTrBhXzDQD7l0vNJHvtny3QgfZCy/gdwjVARyv3D5yasaUKfNeJ3NYrQic4I3
Hudr96nnUwXVZsCemtgV3Os35L7XFSPxKIgVfbC6MavcnmgNo8A/XRvg1RGKH4/U5mbw1f/dEvqb
3FUdWcwg826OiIwNXmYczKJapHc9ogVt8ztLNO2gb77iKFtUAwpGlbP5ujJy3IZfpH0Qp6xXT+Vg
HxwZpt1VHkuTJjJKXQ3of5biSo4A0PzYciNO9JRN0AEhOBm1eY9dSwaGK5XsLAfFHjU4ALUVr754
fBd/4pufTsGh50ivn/UoZVZ1vFnvfPD78HDQGnaqq8pFYDL52O9DVNIAMJfDCq/dIMB1Fb1m95dj
TvmJU9gCxwTXUT0GawN1G5NB4zJzUUw5xsHcWtQvS4ZNEOXHQACeW60OSYRaTsezghu5PeljnqUc
y7ekkj1+3/+PdtUFuYmpGnuX7/adW+w1ycojj5rdFJxg2bY6zqD+qgROwXmiywZF3A/JmSDXGhCx
dL7IebEdNogj+Cme9a9Xk36/YDmF0+h1pXBU9lNHM9vMIItkLQ/Ze489b2QTyjd46le1L2LcnP7z
BLKt9JK+AyYxL9K0NhwceuTPRv96YxFE7I7WLWnaeb796inbXF5vamzvGC1Ka7pUtbhyrlm/Rmi4
Y1gqZsYjlCPL+IPzmBuMYq78lra0DhqY8Qb1KgwvICjuZt45JKZerznnRb28JObrqteiDIxkD9Y7
P5o1Kl4MTW67J7Bj2hZADIK8zxl2YJ2gpRR9M6uTCIqKkNOevkwoHszCGWQQOIPs2RbgncdlqwhI
QUKL9hwE9cmmvmzEvuE4pcpg9P6uC4lg0ZkVIshQ+9e8Qg6pvn/vuCcriICiXbeFRzsp0+d5pByJ
51BEU67Y9Q1lCkPSh/leNA0syq+amQSCgQtCAHWkc5qhT0hEmBWkSD/VBw5qFMht/zBf0Bp/fxg7
DHk9wYGKV+k6qNCyBThnKkyJsM7N4sEqrJnfxehLHDHhyQlsQV11oPtwCk9X2T8DBf8hp0BZaEQ+
GiM9nCpspax6pqyfBMTwHWKrdvmQNAw0T2z+AC/+mabqRfLxSGcndbTEr/eKvanwFn6vnk/+5nB9
JfyZXiUcM4oX1IeLFgpeRaODYt0hzjmRhWoRnIK9d2jRL/r9GUYk0PG8RemLyYC+ptf47ALq6mUh
zMu++1gOepAnM5VIRLNbCt8K3Eb5Jq1poVWv8W4LSi53UByhLFre+XJ719UzTPgJJ7Vr4UpdOYiv
TH2rUAOPLsNjU6Ka+7/3CW/93zZdpwrDQPcpgR8eymlVfnBWr2m9UlU8h6g6KOWJ3htLVkLJWt4F
z97n/fMoyNHVyn2AJ32QvbRz8JQOmguFQX8oMqS3dygUNmc8Ob69+xKCLaNrN+/e5HScWfKEF6RS
/7IMImTY9QPrzSGsONWFfPJOO0UCNEeDDPvNHd+X1NLJePO6wAziyHMmJonOOLgxOd03gfnhXC52
eDIOE5C2EUcca/3HS2194+lACkLyu4E8N7FVAoZQei0OdueL2MZ2mPJnCTNiNWESa6iEQkBP55et
+Zd+b+N00bEaaD4ucyX5qLU4OHoISVmjQAhCZlF9lGOl0myxMlAAaLkJft2as9RY7VVdNmSBP2/g
AvbkQWX9wuoJ6cLIB1Qr7X4nZQP4Q7Mx5b+h7kGGas+zSwvYUa3ArPFXY1zz4sFjs8nvPIMdFcBY
sukHS/rtICSJZEKkw7eLoj9iUr6kZGNpdbsTp2G3qq0pWNV/Ml3gMKVPSCrLlsl22jILGPq+ZNss
XiJmVIQVoA/VqriAFcyhY5EFgt3BGgG1bEXtFK1eRs52o5lNuka3lqwKCzUt2QLnnn12iYHXWRC+
ZagwEFg9hwosWUKdB8q40Q41VcRlKFPuyV5ysbKpk0cG6HzLFCCfrcO2ZBDkm6emG4imGrExFFDg
WRI4GtJr7r24ft1O9TcBnNG7mk9MsmuEJSmX9rb/0NcaRa7mn9s5SLklrkofvceZXqn8yN9V4vZA
XCEphArkRuXu5A0VeAsVFQHeIVXFguSJaOzSHljjjDnGtrTHX6YFC/2r2cpBdYdNopA/IFoirMBj
Q4nhYMwGdfp+9aI75hhQdYOby3mAeEc6Ta6YZxtRvAzo9hwybltfNV7HjUnVh9cBEvVCnzmBsj40
axzHXRXILvxzWomNraTAlN2rxXSMX9hGx4U6Qrx5jKuEMC2iycGl8Gtq8g4Bop7ZiCrvkn0y284v
SQMz6TA0dJNyV6lu4WJgeqipmzlWqSDJM96dbwNHJWvKXy1rJXOPlcX0yWi7rod28Y+0z3PuCKkt
MpFjne3ZOHdsbo1cIyuqEDenZvsEL5z4VsL7jh5z7DZaSehqWmc/zC9yguQbIOdMUwjBJJaaaQQM
Wcvk52vYk+AwfKvTNdem9p8nrJMbq/qDF2x0rK4Xrzy888vN53z0hWDplHfcKAgod/YzWHlmtF8O
a1gG87VM+mqVPBnSFfZ14qeWPSrWeJpENl4jrcIkPEIP+KbFipFzAoK2caZiEanpxmA1Su3eDywk
Z9ypBfkm8ZY+vdjEFNi9OGKmgm8UtUoQTVKdM1hq2e7ipEgdLzjC5x1ETZUrYowH8m0lvEFRrWnt
MuOzgrVhyv/x8uoRRl/p4ASTQNASybQNqq/c3R7kUt3P/I3v54RoLqpehL2rHz5GWYMpbngwZL+j
/2IHLY5kMz8yhg8ujT54mBH9sIT3zbLtInhr9hVbV2hIHAhC1wy4xmrEJbaWtU8K3CZI6FALmhFK
fB2Of55QtqeXKl/MfQcFScKhb302gejuQ7C5SeUv+WcjYk0K7CP+xV7Cv09v9Naz3WDfjQ0kP1qK
fDyhb08B3xglzDQ8ThuA/vB6k4THYvbXgKnkwyzXm90l9Tg6z757DoGhjlW7basxhpRxPZt2xOEh
yNqJ+TnPKQppfJr0UuYL30rPV8g6C/uBQwaKD6yPgAtljRsMIYN7PDZbRcwB3PW9AikazQLXbtfU
EctUWqQVZ1ecIVBBY7fHqqM+VzeWxTMziwfnjTrHK39g51FzF+4rxBSSALjZowkNwrqhzYtJaq6r
Jl04ygUokjwbl7rolvN/MnPVR87fkmKKElEstx6Qd7PqN4QyJyj2iYKTeGbIZgz2KhWwnI9prgaM
/hRRwDLQ0255iYEEiyntXQwaAoXqtAOkAeuIj7N52YN8fY/EQSgUzwa/SEge92iEctNLYqnXRPk9
8hKULtEKP83V8RQI3r5I4BUIKI2C2Y26x+qc9oc0GPFMZxHU9UdBAnD+dfox6r+AdsHDrtXQBHn0
NAXbmOS9vdJIbFXZL3FaP7b2BQKUgKIDAR/pUNL8GjkgtS45o0+893XnS/JfefHBCQYKXvt9lGEC
WOF1A6ADw5XO7zSQSqGwlgbA5nLpQxRkkKbDG+wgbR/bJIEw78OuO8C4wJAvfdF/DHchyhWVxly7
7DHYY7jFsgUaLBEHrBtAa635obEuBfxCPZbIxeD3OmrHE/5TtEVvk35vqw/bR4yNagcvZ6JnuB0C
vTDq2bilyv3dafZPcnmWxeatG1mWx+OCzjM8AYh5XpendKYdQkwENsxAAtLr/plmUsClKLwsfAKD
Xyusju5ikKZW+fUCazXqdbBe+VCyg4YalCUOIwB/yeJR4VrgqMtDDHawUk8Zn5T8Sj9mptLaXS4F
gKmcMg45feKLqFBX9Li5f56Am/pLhldV1ZsuoI2c9AMWDiiQUhhP4FbNkhQM93d1Jeo+cGuNRdBz
aI08yXv6rkfJgeO2LAzxKtX4Mv+g1rz625fbDRXvs8bIkfQ/tb1qOYYjVmAOYyJOXpQOTHzsX95b
s4rvjxVfDsfAgUyKPQSG1YfrchrmdyeDNAKesQR+xhuFu7sn9J7UaahlMzaeUYhLsj/kNJLI1kZf
pG2Yd6X0Ge4a5Cy7Ab1tl9hDJa4D/eeKKZzp9Dxn0ZNkY8CUbLvmlPIzP1S4HvaLkfImOfbNnqaN
kRkwNLS/eqn3jVE7N60KW+pVlqdySXamwXHJC/eNwnzNlIIuCavbnZDhKMR2DaRrH+DkY9K5a5gB
fbZtjp15MuJZadgXK3H4cJrUC36q26W98PAxcq4es/rLVhXE3FPB7O8Tsr7LCnn17PdA+py5dlu1
rFjmSSKnwCi7Qbr7OHvH0PJYUyxrqj4rSAmYXYHyR5N0nHswSgJkW8ABnnxNsWoE08Js5of8ZGTB
tRhx43VbFZF1+OJgoApkQ50RXiW1t/bIlTJwqeJM+iLKp7NAefzoBwlF5uoiIiKAmZ7hB45ZwFOT
6yhpljcC8TJx86qNhxpLtUo/MY1/HzP1iNgy/ALNnb1xv79+wmycPVirM6SfCotoIBMUKnTDcWUy
T0JqGsJt0YOReyq2TB9He+3J5r8rMBlOHXr3i7ujJaNFnfgprBJmMDSU6Tac71pDxa9q/N7MsmP0
pYy5WfQg0ZJbQpJ7UhSSALoxQ0r2bt3htd8uPvpcfOY0Bn7umm8GVZqusXZ9ZhpCZSdpTU+iasSX
akqyH3LqhW9qbYa7+ZbnT9fPwctHaDaX8BzpXBIRMxv4L5SBTf/BBktyDPXtPmGC5Vhf3oCPu2PH
BtZ8rPBGDf/7tdTVzOTz25hJuFT/2h2OruxtX9bCG2es5ngg3SXYnCI7kQ0YnXOfSZznkMCXuWvm
4S30tWnNBpzMjNSxsWYmG3YQZYhfT3qp2LPd2zQGjWzP8XqtI3/69J808oJskeoFO2uw/JKfFwWR
nlaviktF7A0KlszEpZn3DHYP3PL/4ORI667iRmnY/bZwHYxyG5Xw2wzwICFU1zIgdeC50chKPRhg
wtllCQrAVynsXLOrtSLjfH3mS7Qqur4Fwr68oGX+tjK/Q/W2kzMxLsFcf/6cy/4mvIChMUX58Mcc
2n8Afdzdm/VmICE3JcKatDkEMCUGHuQlPNKlqarW0qsI0Xedb/h+F7EHEdv452bMPBMHuP//qpoW
A30JkNZUX/DUUPjQT2l0NK9zh70SF28mlLiTSj7Vmi/k9M87x4Yj+xQ2TxmSgrA0LRe57I9VEkyT
PGzBjlMVpuRGy7na60UwLIQ0VurA/MeFPMK5mVzEVFwzyk2Fs0ucxw6IIdRk425375lf36nQyK3x
1WET3w7ps73/i6TbSjg8L/arM4m1FNy66QGhl1SVooAPvvfByRmnYPpw5QViUzItlVm1l2Ztud/O
jCUnwtu+02RsTWDXFcu40qEbG5W3VT/PwLYYljZo3znOaNURXPF8Yr5YA4oCfSiwoUc8gc5rKAf1
yLxUCihDHrEWqzM28lzCtLVz89Wd+MVMLVgOmlDEkroyV/Jeb6qqQKUt+3c7dCVZHb3b21cFxF/0
ymi36m3UFqnKQyX7hQK9m74ThdRs0DdL+svCPPRVtz1+1lKYmEZ+KB6Q4AFAWv4y3fBHjwcl0zSr
EtSVEeWVg2Cct9E7+fd9Nb33uzMSVCs3gjGlUkBvLhs/niOPZkNv07PxVsnbvkzDvzAFaDN0NjCZ
0EH6wU0FU/lhAz1LLtdsRhjd4MxSbdSEabW7NOaDgqd85pPaVkVsK4tX95HU27a/TGkqCm2q5mCW
PlnsE8wP31u9/mO6dN0ociJ3pcizrhRxC1oJy/z8jWfIBvn90K+prQ5HtH2vqecP3OyTCH2ieppU
SclHW/HmK78KM0oJP7hTo50FZHo1O6irfk4m+mc1Dgqbk3nXV/983ABJXvoAG1jrr7+5u3lz9roD
MlSt0JKWTWjLqMzZbe4T50PUzG4hYHDwrwg0akAOiZxVDkL+BoC8OAsd7RJ47MR5GyGTt2uSVwDp
aa2dmeP4Uk9hRekO8+eTVa2SbCS0yh7bGtyJAVSd8lx9ZbkL5XF4kk5l5kM42esxplOqrH8Qmy2f
IaFU/ltJjW7JmuHEEpamo0X0+Y076b+bf0VBXHl9aacdR2NW0ui1yzM8l6/R6WbvZ3LWtM8gwut5
1k7I5lujin+8VT5ZohBBLxTYNX1UQ43rg2aw6j97EQd9PbbokSbg7VpuryQzJ7LljlaAx0nFwuK8
/QaJt46L1x7qGZ+hrxW1IYOv+iHuIgCGSrI8P2yA72bEzXme7QB/1ACgS+ufWDsckpMApIOPnOko
tzKaFkYmS2gm7w5A1brngLX1XD8bHeYfW0uUW+jKzhrg4yh2SRQgJvmKjwzpF+K9cDoEZIA4dU9j
gY4u+VUVlIcKKRyDxiO7UtmtxYybQHucvedfzpFtDj31btBUJQ6CP/196EKWMak0dfgdPNFE69h8
tWTvHMmVHei66lhQv6A8SFOLvIhvqlXckGLuHWzGscojErZyp4J3n8Ak/p6WwuKwjwIBlE+f0uom
RCJgyeKrTiuXROypCuJAiflxoXxDM8Or53D2UvtfByTZv1XyE8f7gFxlKq/Kx9ZqF1V1vhRYPvln
ihHmzz06U3S1Lu7tUv0GtKQvhI4Zlp6mpI2rExBTXsWQpQGMmrk6sqvWvf2WxbCk4vmCNC+wTgHS
vxac8Vaykxx4609j20XpAdug0HzMoHA2IRkkcAswWkUXW0QccF5+Euaf9sxZNJldU4RQhUg9QOnm
K4UzJDpM+gduWqPFlFqKu8aWjGpoKwixOoCUV9yWgYTKAZ0GE6juby3+m/3CCvPMGBIm9nL85VEv
mM2wXcLB9z7Az4xcReYYQ09eggJ6ho2+PLcLsevmH7FaI058YYUMMGo5MVGB1AFnWgFSc+nfaEYb
NHndvJmLOeMjpEuyErJyg9l4GA8N2KYBQbo2GDc5kLIMiqsl+9I9uGsB6xNMcZx7rddzSDmNfRWM
zSXmt8M1Adm533gRwFLdBL+CTaFV/zmwQnc533JkJ1h8R1VDLn0CcMFsmPWf6SKmNuHuE5hP4H8M
yePymy/eQUukuN1no72Osk/32eELBholHq16P9ZFUrHnxvKPORqNce3yKGEoiZroO1I8Ogt0AiWg
Nwj9S8+QhEWqi5StRqoyiky28fnIu8tcL6l9zJNRrL84KsOg8dMkuXEtnsJiV+/u5ayaBJ6sXzDf
c4PAHl3vd0wJovrTS9KDPCYRYTByV/+KL++hQ5AfOXzsqPgavYefpzePO1NPTUSWroyuPjk1+19p
H/YgshBY+qJqXRbfS6Z7jWJKkE23OMH5zmkiAC8SvdYODYPug1orDNwCo+GhisInWZt/YVTzcRFj
wJsjZutxnMHaVPsMr1tvg++XQypY/dViQYV8Hi6q4RyKtdS5rP8B96Jz3ZmDUeWPfeKCGTYDhu04
YtUFtsZ/fRtQ/xFnSwe9LwjycITAoHcXklDxDHyXSX+CsFMLmGb9DF3rh+nVMCQNyeKYmE8hjXNT
3UyEsbKtCEmgTxXdwQUEALWnOryoYERk2gsdWJT2dBjzYfboPIqqGE7uUOvsdv7Zb513HLKY8I9y
aXPO8crebqc5Boq6bk+N+xL06SRZhNScyBxl1DrfukshkzTFSHGGHjpNYvuLE5KlImqqBvbv4gKF
MzTi4D4obzkUur5tBV7RNFLv8PvpFYYiRVIm3D+iBaZ4sm8B8X3VNj/XX+uojW3xg4+kwlt/wAWR
RD/kMYJwggBPbKLM6F049UhaOg/w26iPAhGB4SY9ckhh7qAYI/lVcuTWI5iw0TU1xMFT+I5Vg+WN
63iSL7YMYrn34TFWPmNHgLrHAuvi8V7xWhfmEDGOKtcwupuTvLRPkkunM7azPKmimJUbB8WgyyuJ
lWhTSZkJ9zpS7yPbaIFl98ZlKCaKYcGwUaLE979BL6z+fq8olBlZMDrgbc/qJRzKulekBOJob+Te
JZlis0Nqbnk5JanlHPXH3sKG4Q657poiDfYXGNYFJkDlMbUTz231a+P9K2R879+meIVJrxUm89wl
AZY7kUW290hvWMq780THixZaxyNiLhKusX8Gau55ohEhx4A6tAE6WTZLwy81kBsmpJtT5UDOKcwl
E3wk+taJBVohG767a0N31hOEloDhYxXkutrWOkuUhiAruPJN2G13XEU/Bd9BZIWgyEbN6r1IgQ5t
2QsTf+G5rRXrrcfoUJlbkxtzKeyU0namaIwZkhxgMJ+jfRRjO0sDQjJaOfJbO//5qp99XQ8ndOid
dY/246xX4+lvfq1TZFB6Sd/zYg2/30bEDvy/xxHSxMltKL6xwFL8KPcaMfWrOiyDEtlQjK4f41D9
/r7tqQp8fsDKWQSiSf0PQcrUg8iFG5ZSaK2JwKxmObmBpqbkYIqmeIDO2/CUXlpypm/DFbbDAR8f
tjFEFzBj5zYmLiGXEKbjl+rU8Lisdj1j1BwW0lLEwUOjpcCeIR41Evh0kDF/lv8wGwL88rkGQvUO
7QeupfeQMttPoYPWCTR1GHhZZ2wWxyzpvy3RauT3QJp/Tgncc2AclbwapWYXZOozh8pbw5wchGZ+
d3gWYE3lA1Z9ibJVVYygwF1+aLZcwuQc8FGEPilSQFT1qFGe31Zy+vvOjmam5SObDC0R2D+4jrHc
cwGxAFQ+GzSNN0o0qpK7w9M8Wug9THyF5NVcmCeMqJydpl8jXf+iVF/Zdz4CU1Q4DeWUrfCEuAdE
q9k6bn0ZTiSCh6/+5CRIQFGYggnYbY35o8F+qXD1fxEUMDN99j4x1u3g2r0fFlQU3ldg2eoKl66U
wFDXbwX2qAbjKl1DGlt2J6UxfOobCXSz1/d165l3JTqLMwyZBHWMOdCBh0tEpWOL3m91o2MU4t+q
MfJpcGLuq5YVoYZjHBqgE7vPwkgEZqdq6Mq3goE2rua2JiZBBuowrn181nUkpAnnFyktcc5h9F0F
tr+IgEpB4iwbQ9h2vobBBaW+CFhrgirQqTjqvdMaLbO9RvQLK7qVh31qJikPBHKQ+5+fRbjLG53I
2jgzUznlj4pSZAqlxffrOzrNLGhD4bBv+cLPIIUv3FO4a/IEMqPZc41A5Ge+XmHLUCjVbLAOWQLg
YIt7e4GVTsQH0Cb3WOGQi9THtYIigH4Pwjy60KqYYoQ8CC3h3J9dATW7p10OCqcjfxmLK8QmrU04
VQ4OxkuZkMJ03a5wLx1jGivtWjB4E2wpowC2tWdp7f9+6uoQuh+lpMZsYVA2ZX4HllV6fuoX83On
caq9mVGuZXa7Z0t3qOYP04RSDbR1KFgbuxUnczJz+4C/nqTkTl8QWylNQRnJv1Eg1/zpsA8TMM2D
Blyds2gZtaLE4E9TO9Hz6ccBccNoTUGdvngERF0ktSaEctrQ1Q4QOpuXZU8RjyYRpO4RG7yeMFMk
FZDkU8Pv+GzwROTKp51z98oxjGuTgqMwxyfR4JiZxFgkn26qun4eXn13R4OHHHYT7L5D1tsAX81O
SMETtG2w3yS7DylLGq+V6lOnEBgkPJxaAuXPfD5bhu917o14WYNSMhybsznweEt0wcY4LJXh4AWV
jQ1Z6gzHLjsY3KYZQXQJQO00vx3e3hNvMRHjTcJX/RiTHDy5MdbyC0FTnFCOIGM4OrwCBQBKU1mo
tpcFbAB95IOHi1/5/AadBp44FtkJDZ6zwP9EKH/rDjB6abQ75o7BE7N6mN+vponlNd+CeLOJgS7p
qiVP2+/kOrbbFHM8AQqZZWu61annIgxhLRYnFDBorYHfAM3gmvhhoE4GQdhN/hDUtquvOKHX8y8V
HEmqFY18MCUpgVVWijKzr54YPcGhpUlnc8ZqAk6F6j6ulHZ6TrwAG0AW0OPVeeIv5+2tfJQZjuN/
QZm/KsUjD6BRJ7Xl+Yx2y65Rcz7KTFoJLrAnWX2YNJieO8la0qTEkFerJxtbc7JEVtifep91dCxo
GTQ3jkTmBDpClm/hB6DzCXtFDeRqNjfn4kgSft4shfGHS8gCOCL4nafIWAN69Suus9VP882ZTyYB
nMOoJcgRBU/Jn79RcZQcJsospXcNDbsL0YL+77G7avd1P1jNFC19OFb6TiLat+0sSawnHQGjoE0J
E9XdizwnxWPoCbishcuk26Diki+WlVCAsSs86a4mokV2cqmNbc99t4bDYHcQFlFC3C/zBsB/miHX
ZoOK/rjXl0boz6+8EoHnHAUoGgGBFZ+iuVHTyUpvW5HcgYwlCrj1HQMwThV/n47DhJIOPa+9+lfW
VkmYZ7oRXVg24EOV839X+9UI6ui//FhsjiH3nF6Oaap8cXMDj3i5nk20W1ndgqPypvqAMexF1P0q
YRIwQ1tK/nViBMCHN7w5ykKqf1iRqjG6CZUW543Odfh6vvvuBVCJb8pzEP/wFhGGoHYxs91n44Ow
xe7WgmP4zZ5Q2u0Nnr2tFimWEQ9C9dS+huCuO/nKMLvFmNC2vLrpqOVAwms9KFtIvRsAtc1aeT9x
02PM0Zo2P+holFgSbfn4Uqh0WlI+PGmTlzH1aD6fVRK2XMn1M2URP8FHCnuWiN59swMIW33bXlcQ
M+8LjYEmMmgxra6fz7A6eHKDnednTMQjK8Lj1VgzMpomvQgEosfImd+Omsd11Lf4/hsl3OU7kJ6B
ycjJFRkxYCCCmmZqHkAzmnb5bkhmJefgL6G6lbLq2nMJkxp1XIkFT1tmW2PF4r5b/eWXxl8A6gS8
c50IKamwIxKvBXdiTU2AJuS+/e3b7wY8LPfOFPncwf88IdkJxsetOo/gIzCsSMZ4VLQrY6HWWmVw
IbRL1zQoW1OpQPn/yyn0QDk4zOWYDMxGgGOrk/vTZY0p7CyuPTpcLGphRCOir6enkSX+LMU6g761
san1ibKQ0oYorJ+Mkg/3bmdfA6oehZpHqIrmdZlYFAuXorGTNwmhLEU1ilb7tCcV1AhOOVSXaR+A
LBnsrs5NAObfxDIf7dYsdT08LCX/jOPZOiqI5iSRthfyjO+EtUPehk30e5eHLDCPvcXxTbEhh7z9
Qr/9PenWEkesIc4CMmaD5t4cZvpNZTS1JnFLKP980SInLoODN0qnUTH+v7m7Z4/9GbgmMxoZYsBc
rOJ3OJ0LR8ENzTss+Nbgz4zk+v9Fk9Z8o2Kfd3pwXlfnI4+4yp/LPdSIk+IyIcSRlFl2U8g1Ebf0
bUB+/jzMlE/E3l1FMZWAlzeyhZuwR5iEQ5HY6GR9io2wlrdWf44xrCS3vgAbahjmOC0OynrZZp8j
OnR7N3XduBCjKIGZ57LdNkwqG6KPzz3fNMJfEbnltjK/hqe8rWkuL3J2T3GHnfpCT83sRpm9VYg0
rWZSJW/sg2ZIQbehYbWP6p4mnnGONa7xbYIiFn8gGyxjX/plvdWHWLVWOFRghcsD6tb+Z4sMisMX
OGqfkOZ3Y2c5eGQ4fDE3EzdCUDyIy317UI1V+Hrj3YbAO4Ohzn2OuWIzcQV69F15it4yDsRrV5fR
0G/8eozZR8NCXmUDURB16r6dG3hZasxz/g1+CQA40rAqCjkQQ5yo6GEaZNIrlonjJJRPG2SDatLH
KCmHNdWG1XPrJs1sK2l4D2bMzr7TAhLXf5gBaRiS/BUGqJthji0eMHmtBvWLZlB1GYWHfM8iJ7+V
Yle3vYiYkl5kyZyRyjtyW1RvVoeM8OKs+gHOTEmUHO+n6yUNjJF8HOrKTWiFqJ7ygeMnsKFKy2J6
jT1sdHxNk0YdZ8qeZYGEMpeqg8MdRFJpDJChAe/IutBxtmbQp8+43zQcmfyHgAIymujtKFaMpZvM
CBp6ZFeoEwY/6YbOzVjvp4n2xpM3RuYDovioCH4o4bwU707/IGogvrdDkKLmk6z7/0j+Z8TCfAcd
oSm7jcv0ToMIQVcOMrny10OhZARy5R6KHvRUeuaaIaeo8rf6bP2N99Mi5bjsFqR/CXdcaXm1fjI+
+mrcVsVzpP//yaNiXVaLnhwUA3+9FEww5NsTl3I8u1bsU+sa73F3nJVxigTSmw1tGtsJt/MTCHic
ikwPeaK7bdNx4o7sWZBwADUenLPJ0s9pHAU8fe6ktE0oERBPz2xh2cyp+Nb1Ddk+m5ZeMhBieLTE
gwgM6xOXvNCbk3Ma5yHiyV5Kct5mKgQV+nRkhJXLCt+5OPrAnBJI/jKuO10jjZfgOQ1F3DeDeZ+e
w34yZ7YIq+sBiVi2UVsOuxgJWWwOq1GBDL8+PevZKZbTwJZE+eaLKWM1ChHcbY8brlN7kNYYWD5F
KZy7N9nCZbYyo12tRaZEy33aUb0jVb/9i1e3d6J62Z+z1V2BSV6pydKtQTjOymQBWeOn1NBpon+d
sh7c+/Qra6ZVd0Fvfo+XPm7J16Y274HKZpvgNfC0qX/QR0pt78OLCFtQ16msRfgw9K5EHIw0Y80P
b0TO4VzQHCrn6UOTrgCY1iK8BAWqS+afzpUhDQ2nvZuaTOHm0l2pt/nH/AVwr57COhNOPNj2NAP2
ypvqaftrKrVuVoj+B8J4WafCbbsKcuoQ04RUqQRW3F5e3hazX+Svk2Tse1fTwFJ2FZc4wSNKe7m3
J7Hb6xe+ILAxtwdDe+mBQnce9kvOOZPMaR/cdM1WuMdZVe1/HgVLl9GCintRwNlz+XiArdFrBaLa
p+2dtywg4RTEYMvK/9k/yX9CfVsV/ZdaSdOt1yH1nQpN1oesbKknlvpogtBgTdGQR2VSuPcIIp94
P7j8520OJR7VMe82VYYKMWeP+pe8VJ8roVnQMgZg510GVo1iYG9lDXsw7YmZwCRs+9UVkchaVoki
8DMzGQG/1+rOSD+MtwpG4gZMnc3B8prXrDotDeDOopovDWnraEQTwYRFaFbCw62LFYjOo2KyTFfJ
lIZDlG1GvJj86vkckM7cjVOR+RTpQLwtBKxxdZVElJGw5pa5IbXbHrKJaH9LW97unLOdZ1bygpyC
K0iEjUxrLkHmeVOVWsbTXwl0GGGHrWiYVwd7R0qbCXfVnQSGKnUWaJRXyvgHKjnnGZJT2MOUnq65
A1xwP8QWJOyd/KjRsE/YWuo+gxI9VVRnknqM2nIuMxkZ9rbhK/9uIDWV2Y7PM9VS2PsY0osaQu9K
khRw8/5/gRXfB0SIZKsJHjy/c6uD1/mBGpYw2ES0ItwyO/VZXj4w2iqs5PoolER1Iyt//+B347EU
5ICzMQj2BJY33PhZBxmnqdCgR1VZm+E38z51sF6X1rbmZOj3xc0yz0zI9c0foZ6zSf1K0z5dBcpW
zEYmRpCaeI8CyDIKaBsYG7y7zo3zOE4Eevyyz5qwnEFWHRcsC3SzBlUJaa7JINi3EECiLr5PyU6G
5ql6YAqYO/gavKFMtP5EnAXugNwTqeOFf0vCSn8OgAjbLviG1NfGP1ElgmerDqZnlWiSR/W/UqvF
hT/lKxNbHdew1SMqLCyQ8/lK7mHvVVWm5mKa8R5aY9qnnTOXPFTtR+EjmqTWb1mMtVKrd5JxT0rr
x3NNfa++/g/R0ciCr0HxaS0Mv20a7fQrPFJVF4yUKfc0KkqwlJD7znMw5y/jhaNiIYymh9zZpgwk
Q+jOlUPndv+7VpthrhwztulIPbyteDq8NN+dv+DX9esjAsiTq19doIhycDV6eeINklp2DgIxO3C/
2mJLbDZyiCKLCH1LsYiF2NGJ+L6b8vLJrhR+gEtm3jgDVQ6R3yF9FiKplizMmnYQP+ivoQHzhmMb
EhBlssaRCy3aBBTWZN2cLnsRTOClyTIJuv+T6qpO3v4qUWkGJkkzD7NAspAETHTEdmtyoAauK4KE
eU4b9J4YQcGEL3YeU2xuDdAZwRqeHoo4k/GTu0BE/L7r2VWh7BjZ1Iay/3MOE3KQQk8BULq5LVpP
0FI2oV7xhovnC5R0tTLQfjs2SMsfDCi13yQY0TeqdU4Eq4NII6t1/NSMKCuKBkRRiyNp0aM2rMkA
DnhLZ86YE4v8ImUpJ882ZzmjZv0T28suEZfY0VODXNgCkT1CoHRxlVwFG0sLMpKkM/dLj2Zo9gFS
ATeww4PCrrcE3HdmK2RP07ckVvZiyxrGHWHuQunHkyTNZlEztU+IvJPoYRblEebfYkMg1dd2xwOg
zG9eEaXeK+xn4aWLO2NPwGWfJgSrVK6kSAXO5z9IJAEs+qyusn4LkAAhIssYSXHfZXsscHxBmd8J
Sf2MPIKMtTfIEmJV67x3dGJ/7wsmyNiJ97O33Fv4hEOtHi7MJO4SL+2R+OMGsfOGFNbWvru6argH
8PIgG2jNcoGedDQO+pNN11yzYpsTvbi7jbjN6/QLRem7YoAPPxqmSkEFX7wISKkLaiadPEwAtuCj
n5Y1CDlFLFdG4b1MyrULiuHmg9+wrlGnfJJm1z+kdrbbjK1eb0fXnKtNzjCZwoTPPc64M3I+lyhH
GoG/35mDhdvayJFQ5i/UqWQMHCRN8NfflfinZH7T33cWzmJUSPYSxWbzBK9ftdqmbgbIrQ3RYod3
e+Df4we4U7s9yNL3KISgFN7+hy6dc+GppEKELAjOc97ewuqgNG3Zm5UAWwm4CXe0yTtVdULBFUen
ErCT6jb10IoVOOdIkYpEVVa3ETVVlQZyHhHxZdbomcarc6wSBHyzx6eL8oTX2MeFeGPbQ/38TPeF
whSqD4HCrBlscD9+I9TAjIEjRCVArShNRDfeNNstjOyKT1Wihmiaayq1B4dUy/vcCgKLBGnunWat
g2WotHo/anrbpLNL/rEeqYsfHKU8eREE4VccRLHkwMUMcfigjVRh/zQIeuPCwYsJ1pGJsgV/f1+y
uM4eg0MYgvtK3xA4MMsMcqDcbHx8BEzfkFMoF4Hg/3Hzz5m79RJ3/l87gSHSI5/oCXdhKZ+J55h1
FnJSopGAbVjrVkl6X1Y6pYtg/Dik2zQctsteVdQjJQ6UWML061WoIYwpVl0ZzF99qHllD+qFZ7YA
BpH4RXRHvBLfSJRWTJiu6oPggYgPY5NvfMHI7olbx+ZO2Ws0/0DrSyzylxAlv4/gvoT4DDhsCAeK
A9nPmhTUPdLtNnejoPUI/AiDloOJylfY8BfNR+1kXn3CJT2+5pBSp0wRBhG6FDfKDYhsh0BLH7Hb
GnwcOgReV0SA90fHOZPGLE+NhbsQ6HU8w/YFaMTk5VL0CYllK4f47i38xP4d/BapBsf9xsBAiglQ
59AvUhYIhy5vnDLsZWRRm+PVLohfLDDLwqVyRdQPRcLxUXLOwsUI1cEdD7n4QtXUN8oaoZR5MSsL
rIS/tZd4iVggZVjf9ZtTGOP0rUlEUiZvX2Q/llJLA9YBJ1R5sWLLBJMNbKbLcxLck6CUTMDd2grk
iMd5x+WIJd5FlVy1TgS+4vwrmKLDaIK20hFJ9taf35ZCLtmWqB5gN9XdB3VKtxdnKIC28J7tFj3D
JXn/xwFr41LrCO2MViBedbvkoQs0aM0HRZe5SDwNsrQzn9Aj3uS7XCVotiymc02/LvqmCakBXWmJ
VXa7FdfHMPZpl6Ht9l9f7dX5RG00/MPzPdYLHW8l5hlkNDdQ9ZaUaLnhKa0oTBikTpgDacs/mth+
jLfiXU1qCmBCFXyxvwZLhhnkVgmJGgAC44xp+pGVPU57lIhu8kq+RbpjZBVB0yznCuBoIHp1ISUJ
Nh0QfRyWxLrf2GEJt5ISQrBxXzGkLgE5DHhI/qU3+vnpFa1ZGP30cqW1bwZeKvzm1sZuuMfvwle4
q0IqlaWGKvOo2EmYKNZ6Q8yRkccqfA5+FYkaCs8O71cGDbdqyIRsDxq7Xg7XfclaTqCPyBRZ0x2x
1bbeAHpcfIeqlleWrUE0P9cb3E5EMqH5SQee28XVTTEEK/QGyUM8NrIxjQMSIY4v+qtaBhPl6vNv
6iTsAgQ1HCYHoao5mdy1ljDGttusMMFlCogE3O2G3Ba6jFr2qmpeRb7xJlPPtKBUfvCr2gSf3G6n
fIHKwcRWjB03t2EMwUhNUAIfyAp9pcdgvdo7WiaNnOZiLwKAkFkYXJgMg8gWCsv4JHSDSaANXn+j
NshHryhbbptA+rpF8yHCxldhMAZWq1DlKKrXO8S5SbHzWFFITec6YIVQDzr2GpKu7shVtjZR9FEs
EL8JEydG4wBnqx0rHyWRijZ16brRS6hTVAlMwGfc6+uBk8cn2IKp5bPYb6pLEDWZpROjP0yf1x6M
tQNvmwiYlGZCozr5gtPGpryi+OzF8LVVZUXqb8dn3PbrNKwVB26oZe5Uc4/C5Q+3/mN2Flz9uPQp
Zgq4MbmxYwh4mS2zTuRLsEt/doJGiv4f3Px4BY9QrBH0kRMeqgVi1maOS4U56XuOhiTrkQ6IHW/r
P0ZG6U38+k/N1EBxdNIS5cqyo1CJ+pv/4kX3qZGSY9ru5zMIkjqEtwvp4oJ7H9syOKV1oZwervTx
XvDFnOdvKHXaDKHhZwJfCk68re/B3BHq/XW1gzRtYfX6alaQEaaEt5y07XPTRKUbcpD5NkzvESrg
fFjhAL7/EaE7Kig0QOmEJvtcGAg4J7MUWKEQljCsvOi/+0csUUNdEo603nQwmThbUSZybk9yOqSH
gLjH7nIeHBw0AGI4ZAETGaocVwPHAiW2N3/BvMMY2oCxbBS6HiFPhYPmbxcVKS7VW7uCd+T2grfR
FoMuZyUxhKTkCH2DEMwh/ZAzOj479Echauok3wDmCWdnDte+QAsgGiTC6hPIMi/QkXTs6jS8DVJ3
LQXu5mrTyzmclbtgAtVy9OqU0k4r67xPX4/vBeZ1hhz1LoKH0sJ4XmK7EO+h5z/IPKN/DU1dggoj
+WHhuGeI1meC2gKsy2lc4rPvOt7RpM7utDDkitGBrx84JnXqb0WRkSPq5g8TMurbc6Ql1WRHszZZ
V5wcMmoxPVtDdsfVL1oNUXgSAx35l7tKGiv96gUfQnNZUoQqDinVPM1XZoDLSwHOUHOtBYsE5qcy
i3P2CUs7k9SZ0xpUXuTzpxaPWGGUILbsas1PrTQwcZDoUujNx3oQxjjpGCwwLWnQHFJ7Juis5Zq/
PcWBgMXSEQEZbjF6ss8LRcKmL8ISjD6mNcHkkncA/U2TtUX3bWRWkpbuq/s2BvjO3t1t9ZWZxaAe
yQEpSkDs7EPtB/g44kdCaOyoNsYj/NZGdvjoMkmTc64vaBpit8E5zb6a/9CmuL5LIxRMGkJf8V0F
yIKiThNgzwSr3VFB3BqYrWXqcqK0vehu17YLjCIdN4we8YqaPxQds9RdH9OTsFbajujfKrNDyp0v
cpYncKnXbAbtL35Y97xUZTDO8kvb571U0p8H5eZxv5OkmULEwt8G9e5o6KgpmtIHamJSrtfR0e2c
f8Kuq2/8RD8LTcyLYNIj2fnMyM29sB60Yn2x1r8RRAfa7Gsq5tJKw3bsLXcwyx0TfcpCcNoKJPLS
R1uN3BdVrHIrWZE+4I7GI8DgtmtL7SxVHfogmPAM0R9FkMu2zs1+jTURPYKPnXNz92bpdPNHHJhH
yFsYo71SOOnSB0nddBsk2w0+caZCR7ZxOVgGPgGomM0MoADtg7n96k89t9JykZZULk6iD0dOdKX/
qMOZtDTmd6ctO6jK5w4+VrhwWFnky5F3PQ+MwzYv5Kmyvuqb/dmi2A4pRtTvfC25r6Yts+GEg8dE
yDvfYObzKZRx+DhDy8qKfvivi97jw+rbrwW2HHLzODabImZO+bQo+iPHMCBygAg0qWf6lhOcTXJ1
lpNQLqWPCSbeZ+rNvDacHNWXZ8VJQkCHEn5xTXTbwbVE0aHLJqsbxWnESHt00FOdD3TIpQcH/poN
nzl8FpCN78N6VbCt489gbWGWljoJTGCFF844ZuxA9Ymdc/H25WhOiGNJeYzF0INnI07vpgbj+4xz
BL9foybVCW370aAG4S0+7Fq3i7MwkZjEglffQcAxYA684tdq8iW0v2MqXXM3zbo37RhU7Cu4XH2u
tnIwuG19x4ae29UvL+Blc25awdSRHKMtTNoxaC2pLxRzaz4bJqhnVMbL9YDz0Gsqvh7EjrWGAYDq
zVhFBTbdpyEQ8gjCUWO/UnjukNbpXF3PzKmqFn41vPJRA0bwpS4RI+PqzGE2Lvzrd/HTnLUh4cbu
ecii8l18eUE+hHIUS9vsfdONIKs9jqYsS7t/43mwAX+kovxREcn68gfJcDsP82GJ8RTU88OxiuQ9
ue5sBDu0BNYG8su+SIo0bArkwypbV3sA0lI+ELnsGlgqdnATYM6mKJdUD+j5wzG/HsJu3yliT6T7
6kUUgPLhHOfB7jdza5mw3rSxjsIOG+Rq3MZYS+VS4evHZFzMjDWsCy647wQB7JTjh470JvxnPjGJ
W8Ts8OObJpD1KbrpTIAosXg70lUH5ddEjjQ2Q32ZZe+Y40KiXPVYGM3Rdr4XHH4IbgOoTqlgrcTK
neOaSQxMjiTfBv6M5ykqALEyapE981o9OxD3dtjHs1V5t/g4hd7rkv04CNfYcb6tpilZQTxWSmHg
/hlxQY7NFR6exN6l3z5+Hcx9B9ZixtKTEoPISn6uFN4uDldq2AufDgyzcsP9xjHAVx3XFRW7guk7
2ZiBF1TyomoI3YJoxwBKnbqJLVYUfz35PMsBnkRkZUlkGY2q2xCNLwwrnC8MBXC8PtDkTABNQn9Q
7KarQJBJ0Jtkphxil0iyPwYxWH93BnjPhr5+8ZbJgWEUB67xF6BfYJoeKyDscnuDJ2BcML9xAu3J
9QZ2fUFVB7vUvWQBq/dEFx3DoGMzMKNdJHgFE1NUenNtL5Kdeu8I8aWbERBDeTycNPP7o5JSvywf
+2IQE6xMQmmni1JRk+oBJDzu0fg5l724gNYvLgljvfmZn1FaxcU9KT/bgUGq/jrmF3xEEWZY691l
BhYdMH1YBGBqaxs+olm/aV1v+EqzCDUVVx/XcURdNkfyMNeOBUDwhb291oHMQO+Pb8K3FjejpAYk
oRqGdi+svIdZiurVSKdhkk6JluDu5Z5WeBcjpiYeFVf9YVb4aQ4je6O6TmnI8wq4hgbUxFWXzbO0
FpKN7EBqyprTypTixx5CwiLr+dS4yPyVTTea7zk9b0i6MSZ/7c/MCCbRJsnE9S2oqNhX2BWHInK4
jX2ht1Tz6Z5lXbAKpLVcgQQYlAb2SEOu8OiAB8HYS0hgBT3qbkjmMO8cAoSyKZNWxGk9Hpg73lHH
wjz+i2xqGpq1JG8BGZdirteUg2EhZlOGtdNIKA+EY3deCLI04FR7JajqVSXsn2UIAAIjVYfLjini
o6HiEhqjOlovJpfv44W3vL9QnjQsBKtzAiZkxd0r0SFofpKgC00OzIhAsAqRK+wqZNoWimI9aujI
VFrq7fGeJItVdlUG9TwA0U5hA7Lxvs9R0626roVLXlPmueSktnUOSQ1QxmdCE+XgQAqd3AHva5mG
EWSLDDeIqMazb6gZU+lU09KGpYUqT8qpbK1Iy96TSrHNTmLBBK4NPe6C+H2EP8vmjp0lfpf6BJn4
FcuQ9fvD9F3/2Vi7ujwDldjJRvz230WW11rsxNnY/3FJ2sERoOPntN1DPT60FuPoglHSx4MDIMl2
Wmk7psdI1CLhIp2xj46NmO2cq0Pm+wWygBcFL82TabMF9+7FOCWISeRin+O2WbS3PFpOLLR7EMwF
1du4L+2SuWTvK07goKEAsmtocLs+193G/kABNdxkb0RxWOmnvSAo2eXljy5o9RAILbPh43xvssEV
KR7m8B5ATHxb5eJFxwEa1As1/Ak7kHRjnPTprpmxTkLFYw8nXmOGqeO+jl0ojGaEpc3GKmuVXH2+
lPiMukgjvojzJFpH3CDowPUQoiWbKTPBXmsWKa6bJJPIc8Yf/6tUVsfFYeTc+HqCQWxiRWwos/ai
ZNYgRpvAHBxVYNIFjRaR5AKHVf2dAJsxZWhCZvQGNhhEvY0gyY/+AwTnZqmdyS6YJpj6Q6ZGIrPh
kHGfpcNc2OhxqrQQ0VmU6tpEz7Rnm57EO8AIGejpOd1Lp3FVoGfwfrDQZbhdboY/11/F6ewf5hgA
CouiTMZL0KhAPy54xs0D8oMoYt1apbaFEFvi41ODFugKnBLxwoWYH8dDPDTmPQ3x7+yCKmjYHPmZ
CKBz79MGElX4rIYMHi7bde6AB32qF2rwa9ip7X06OalS6wOJu20XLpgwCCc/bec/JzpwrEMYHzUn
aVJAfxEytb/zAYs87cW1xKUGuU5RaUzBczgoxxkH9w3wh/y1dOJG2KQmVDklXSwN0Vz7A4FX72WA
VzS/UVxQdpvInZxL+Exa2/EsOv3mSjvX6pbwLDcfDq01ZPQk4aQXPWw+IrmMLQVqNP2ZZ1sPi8pr
tmaxljR/rzHbORmNJbKQB3MdePCBajvZemiarhYScEr1CNBdP/W/oFfxiGNFDArxQVNzRvAc0wES
XVjKa38oBBFL6i7PMkYj1D7zV+Dodu+K1oOGuwPMXfs1Fiz0Ke3IpimYLNFdxSY6GPIqKVUVax9U
L2KycrDpwdKpmX2i3mbJaTB4viI15CnunMMfR/DxT2A5+UthrTWyggJpNqL77v+4rhG1iwH9RV6+
S1fYAyYCqziyieFzpLFGgOKCbzQB1SUW/X7tfLEI1vTd3Ytebv8b8skJ6mg5hilfkQMRNuQDZnra
rRWoOmZdrsuDcOkm6kkPLpRBxn34/TcwYcnPbfJX/FzmA7wpep/pdmW2QamCbe+ulbAubsN5b5HW
N4r/DF5IqJt783dHUbXN0hmP/DjCJV1tOJpFUP9TH/tdpCV/8QZDSdNHzX60g2cpvP51ktBdvkcp
6rH32jAZBye02j8DjtE9tgwZCQCe4eGjTfFqjeuA/DTjaTna2nSP/qpqqjWKdRpOQVGymHd4jTM+
Ee8ByyPUPw0A8ZFWqVehXf0r8eeMOKurkvOFmCbHFUIGCMnR/MEMTl1ef5ulJ1/PTHDS3ZzRPYdd
4tKrMDH7w0RwWUHH2Ibjjr9xQTZcfscF/zRadCsdp5whSK8xfVKjshvGTYlDv33szIoIC7RgYD5V
m06qRz1jeXGUKSAFIgQsE3AYRKSCGG4g3pvB43YENPj2jOf0Y1lPHneSe4auRj5meVAoPLlO/8vd
yEFVQb1UUIoL6mBwVYWee0Mx5taJCLwBTYzLQSeGrEqyvgEW95EpvbEbHgQHUtN4wSwgnpa3jkra
xCx0D7BlzMEYMLGyZR+01DbUUfD+S/95JmYZndZ8MSsTDX0Qo9ia/Doc8PQm0MuL3Dw+w9UcbIEJ
YaIq5VLNaSXK7LuacO5mE3CciBIcleQX5kD87AIKcZeXWmn67Kp0A4TudkVlEZ1EaoF9dex/9bjK
xEioFQofMLhjRC9tBuC17eEp2l3ddIwmO9j7kC4SSz35+qZn1rFKeYJ6aqPS63M8FDbAZydGNGpq
1d6Rbd912akN6dE5iSnX2umWki59D1VdijELvNt1YKV+fMOci63l5J+GOk30AZq5LCcZ4/e52dig
9JbC+/gKbiwwjUXZdKsujoj5eV90+qTMfU3rAU3kVVco9bIckb8IVLAOAoom8VU3S7uq51CnUuM3
LaFyTTkj1UmMphjepfX6TKjE9725zJYZMXk0QnNyitmFwrd6tB/8rQ1FOsWchdxxhYzqgO507Ffc
Om7Kyfb3BQLjVfRBlsn/DMZAxvb1KmmUjU9iKu9wT0GbtwHt9tQt4H2GUiVYeXqXSzjYaT9UzS1D
dnw/m8CpVJP+WkKG7ivqVZ9miXMc2JPEkdSvLGWvQPEnUxd0dPBTiVnl5XIQNhISi1nNJJ1z7hQU
IVhtZlaii9FjNZKNLcAA/07MT+/t+o9imwPs8gWaBljEiLvOY4RuR3IjsHiOu2DTMZ59XvJ3gRBY
i9BJbr9MlpfBdG9TjocyhkHIezJczlSR+joSzsZj+OBw8OXSKK5+9HL+rTI945w8/rnP5cG8TRBT
DP88pCU0bn7+PBCv5zn3b/gyWiK0N7uJ1pnby1cw9SHRRT9H3kOqMzIk96PhbYjFy5//GHCjdRFg
Yt/NtUKHXA58PRWaYoeb7yVeCG/9VTNFEFBIVCdoDy8d9/Z5SoF7fn7AQDaMWAWKtOzPL+JE8//X
d7JM+uKAgHq4sQLLvzJANz09IeOwB2ZvPGvj9rKrDJ2WZ72C0L7i0TLkUgY/pC52mWiQePQGKfW4
pdgDYZxc6powMRXL7kwzTlVsDFRq90jn8hrKFGza9jV5/9DrTvUWelCsOl6aOoy48Aw2Du3oQ+hZ
6KAzcDdvm4epF6M+ZjE9hPKsb8BpSCdFd8hR4zhS0sbyQVb2EllWTOyBpdCeCRax6FhKRmjWY3n5
ut8bIniKuwXx6WBkac8Z9EgXdnhLTNuMzdSGulixfCifdsHZsKz53fsa4C42nQRBBrfNUR1BVi+Y
a2v0+ZVQrP/qNlJv/elAueKASbjKC8IH6q/OaMs3V/rhUh+segOYtcojufoNNzhsPXG0lfARtRX2
RG/ymT3H/oEkiFRpXDNUjTKQ5dB1JrSPNWruuMCa9pSmcOOQL715XPBtyWPUDJsKFFiqXjpEdf6U
IeFUIJpjW6j5rsT1yHaQzHidrKJ//rg1KNx1Ps3iWOQePot3S5r/yL4BXa+h7VVSOcwut3BFlGz+
yMv2Y9mMZuSHWIao0NhSLowPj0Ut9SdTUGK1E4++8cf0/UvqAGMEMkBeRKNHYZOESEMErLE1aH/J
J0ixwlbjcHIuLP+mEfpPcjW7132KWk15KdGPvRy9pRQjNyzMk4eoYSs2fgAWmKaEyN0HNn+VnN5w
OaPfhohfleXggWZAQB05bBfIuVPI8qS5zbJVCc3iBfZvSdtaEIiKLtw4iZeWKYb52DWTmSXWBGv/
gSvn1KnwIhZpczaqBs40aVa3Pu9tES+KmziJMQQUjfyrS8rMZ2dbm4z+RQSo1n22cz+fFfam+CWq
NlORV+Gc+sOKy+yH78NcLEIEdKbn7O+YStpT9BZ9AUar+e+67++R7s0n6FL51PI7uCdrZI0xnNE7
XfgHm8fUDmJp9z4depDGw2fGtFwX99g7KA+NvVKjhuqEW2NPPNZeE/vpG5Q9c7OXYAwjZ+PGJ0vE
WRjKvgz2eXKMF2rRZ0s8PafYt6bd0E+0D1I5WZqLv/paukBtPUmNIc90DDDv/qNss/acXHWR2Zg4
5HlsePRW6RMG5Z3PUFTbtZwZJ5c3T6evRZYKnDzDW/K1Hyvcz9Bhpv4QwsjY8ZVKMQLJOTQDGD+O
3v/mVAl0gmqqxfUNzSUfANV5sYn3Y5EWXum8xl24vG22tCEdkx78dWIud2sZkmlzXYNxk0ZlUn4P
ZmQhA8yEL1db5PrUbKuiWcKReETLJTkewCRac3mWSf7WIxqieOSYewhmML7rqHk18kCH/SfPzTlC
KWKjj/9apSdCCoEWQdO/R2+4K6H112wPpMh4i89pOXPYZdtkGi/tKNaV/jFVLov7iK4RFqo7+PaE
j77SI3H8p0soAWok7TgBIcNQZnBwoWdAqzhi0zVx3Hdii2VcNVQfkjjEWpvpa0rp+Tvnk10JHpkS
iWYxhM0G5LB101nLiUDqbuFB2uc7pWGIlI+vim1d7Ow4anTFHOjT5Y0VTIbgjo06jP/7VqbWYqV5
x8UCmf1cJlQE005g/AShpqI5+SafFcwOxHqwnRXD8Lpaugb1uoBpBHszm7XKaEM45S106ETQhlOF
aPNokEfJc5OZTPsHurgcajENyqKIGWUbjTm4JXoP2mbk/Ruq/qQLkudUIMYFBktxd9WCjaApaH38
uaEkycbOfbaJysRFEZXbglPHzCdY1QQFBMJ79UR7fCWFe3jqUdx9ZczCeSPudOv+o5DiTJIQSN3c
rGV9RUPKp5BEjwXsUDO2mGIZ/33Sw/2+Snc7lcDjgKLgt1nIk3GiXM1zQ621Ue+gHspWXJ2yetsE
q3SFT/sQIjE5kv4VQNqMuj21mwoQz5FYMChgSRKM3/8mWc0/L5vKS/GovwrmGw6imQzjwUV02URo
VlO0m/AN/YDT+Kwloj9bFYuOT+7QBG2O8VSndBEv2thkElytR1NpW70vntUNcENzbAzTIwjMxxuo
usU73iAgedJ16cvZKMgVuGrrOwVzgN0xA+bz41PG8Y53NImzr1Ba05ZIEAEj3hhRzbO7/6Bx/x5n
xWuK17W8mMGCHvg8Ns+/G9zPl9IrR0NtaqK1ihTXkx9r83Locs+9PE6iVN1Guo/FVqgJOMeCQc7U
BzMkn9TXrnTzp7T47G4ufhBpyry5UyvFwc0LZ4g2MIuVXfU+jFCXeFMvSGyaQf35p9BUJtD+SSZI
aRObw0bdc+aI6eOdQlB/gBUVxF/3C5Q/XS+am4nhgsPa2E3UijEHCfw2jxt6az/L3/r/E3W37Pr6
RQ71gRtGkSWaZpOyWMJKh91urn+llNU+meOjdK0x/0t4QjQTQrRZa1nTsaIjyZhueoJApg8ZODX5
jA3RRJk02s87Y3q7rtJThf98Y16CmQzoJNVA4/yYkDBsc+FWNovHSPakXhHNkKwbjcdyJ2wveaSg
q4fTDYWFJ7LK6abxoSCtVO/8jTj3ZYVb+hugbBVYHJ6ge78px456WxJtnN/jHcCaYdOGle1xhNm/
wv+4bZqhQu2hayq3GFl/ZcFmVYXloNQz+M5ApAdZh3Av8klFfOr5RrQ0j+0L6rENUK8u4aTgmPGh
9gb6ghwJp+JCHHeoIWhcaUvJ4IkDWVAEeGy2oXN5f33NpGvv2Dd3rrT4tZxvbu37zroCnLxhSC01
f+CY00Bgty8Hj8b+FGkIRT77jWjagKOZdql2v94AOp26n2UG0kMCQPf67Ii9HecVImxKZ69wgNHP
DQqufWS82Qu0QpgMMwYZSxvlTJZQ1qW00QzRDszozuumZG1dw1CZrz6LIhiSgOeWOJ9T+xrkr7pj
XI8DRSp19HM0U4xXCwpApkiqv8q9/PHfdungSOoa+K8CG2c2y6USDA/PlkPRfsDhi6s20NEF+mgB
ogR6pyinD954v0lj1jmhQQVD+SX+CA9WJtuL2UP4uWwpC43psBvXGXZDTIpOjZivPpyDXy/BalAX
gNcdrNmwsLeodpHDNGFu59hr0ukMsh0VtMTVwFGhcSZ8KIWoCyBuCNJFR/SkZEWIKuXLtYjoBvVA
BzyIwgqBDtHR8JLC/3CtacHlMg6Doe00jb2EKWBa1VTOAXiwNUUwDk8wI6MT4aPonVTaoWma+yU1
9aL/ymXHK5/UBH6JJKWn27RI0mqlwpp/Fl8EXWlMSmFJoxqgzrPTjkpL0NNkLuoVF56eRmGDjXhT
JIbMaz17HsHb8WOzH+Gj10xotiD82dZetvw6skdrsoSPIHbSO5jgi04x778jOVO0Ep2TT/BASUa2
5o30bgloZ3lZwBUlJe9e41IE5oM38LhqiYMhmvDp+DedBGOt0WNNUiyKjaLh9FiW+kKimYpTqhAX
SkHWnnDMM+3DOxk/FhtGeCwL7SIjoyH/cVrOfztst2S5ZNJ9+MdWfqc+WLoJk7HTIKrkA2KIV/Qh
B87tb2FaeHQi306uXsikguSDizQuG3NZ4arU7PS1AZ6jPtV5hRhvNft5BdwOuLRFym9Yy7ZGLdsX
WNgEfNpoDluGhDBJKU+wH73NobAh9f60AWoJGoyIJHum1HYGSJpUbhWFcYbiFa8lyWCBRwV7uWth
IFWc+UVhm/ElD8xBi+3ek50UqugU0/2dVZ1fv1eLx8lnZiPJvd78vZmLmsdPzCR/oUj8LChZOG38
rWbR6QzlzVtxYBpKihoGu/q7VBYywr1Q7eSINxNGRqYeceJK7/fBvbGiXkcEbFWrdfODnJM3NBJO
8jpVNi3FTzRvljjCiPim6V+rOQwrnIcWpNDnmeYlT+xArhHffvBfgHUILvxKs/1VDlp6rf2PMK8+
hf62T4C7IWCuWybDq4EVKrBt+ooj6oSsh/++ukqkZQOpIi0rQV+hnhh2veqLRRd+4pHnNj/WjTLO
+QFmT4kNxCazbaltAuFv84nl3sF0Oqn9jY5PRvkW2ScQPMjq5XwaQf/77fj3GdKTnBGpp/NJGRKU
uolGZJMjMK1r2lBSft2x8ZrAdjdYa+66F4DC/al4EZOFVirVnLxO3sZgKC8+Ix4TVnlYkfZA+tvR
EH4chWuqXe6rD2DG1G/78CjNqCHt5j8Fj/5AHbqRPplaQIQw+W+2Y6ljnyAalP4Pcr6ZF16hgq0m
GmAva6Lg9k6tbdZZDAOprtSc9criyQxELCmAkLBTig9bIo2RmwsQgl7AnDuFDkkmKMrdV6NKTucY
AsDIrQcHzY4I97lhraHzC0/whSOEfvlemFWBZgRTu4LnsGdUNX/YXwUYn81ML5lGsMoIFPSecSuT
C2HUERlWA/UUYGF1FaWTQ7W7hltDIurwBbwgcqe0cniuCaOL1JtNhTX2MSD6Dl13cGRqVL9T1tut
87972nYpA5JS+6osPtvZicaGamGO3b18isgtrus99HI6EFCi/Vnwkf9W7AqCpE5QE3d3sfYcNXEZ
aNw7/nycJ8xSnChnUVAhad/wl0wl4lQBnRRxtn22+MsRDeJwRtC6BLTeWo3qzy4TcCQ3iPXpdIOc
utKgbWclDQz+fbLRJX+goAl8Kz6vQ+MTFQm6vFYIgH/mkGcSn1Ju7SDFWrSr5aaEjFkiOVdnl+qe
c4FIqdl32xa84C66IVYT+0PIYCNcykV6MW8m26V26TkReD170Hv6ovGomua6YdydmWCgDxxYjI5l
v8KzRgoD0LfBBT2kl0BDJA2RfbXAPFKiiJZGi2X58l9tV4sLAdiY+bJHfxhDDT5bkTPYefxqyEKy
Z6B48j7kGsqj7xNUTIx6GQ3Nv/M2QSW6ayGZanZob+uByKxENIostsdzdyEh5FC8pNdtuJNGe8zb
Ha9AoXGGDzy2f10Be8rE8qZ3EM4HcS7H/mH+sGyBJ2dDntp3LxQawTz0CEnZUQYdLeYVFpmJu7q6
PQh8GBs9Y7vHIsrHIj6tGiRYzn4DtCUkMXoIG8GKnQ71aK3GfxMN3QS+IPUziBTeVc6JaKYTGFCw
1QAvpCrHCCvKn4nsrDKU0f/q5c2FrjAaVePPKg5HbYl3teyDdaAj1M/gLSRefiWEmNLNtOB6Iwto
7fViKR/jmfbeswJ6+AKLBOuOYtWxx50aU7zEMRp2CK/ZFYbQbnwmeZBWqLrA2W+cjlQspyOsy+wx
9bpvTKOu0IxRUMJ4Wo/59ABwIpYr27kRDXJybNbqKgHq3aJethzexOKC3kFTOw0nA8oVk6evEnjl
ZwJT8jd4wi3E+fhzmKQ9uakAlvjHF0X6k33apYNJ5FwQWn2LxSfVVRRZ6yo5tTcE1RL4Nfhbu4Gi
CP3XPG7Xu/2c8MNZ5ox2E4icEZoNavrm4jEyLJmMRVAC7/sE55HjTH95BkkAN1zyWyFXRU7YzAbQ
kKg2977ctbNnSbm7aPk3Dw5Tt91qET7ZOBKFW3cpMvU/gxA1OhsDFPy6l1cGMplHyYhpuKH1UGSX
ZiT4i0CkeGVzurFauN9tbi+GnoYNjsF13Tlt4CZfUgDd1BZVJRQWn/LwY06c6bo/FScJ4LR/vc+E
8EwBh7qd/fbPQAnUnoqLO3AKoOva5260prOJyMYxn1f2KechhcVavUbdJ3/Z2o6jt4Pt9vuL1pou
RT6S14WuSL/Jp1aWTMvK+JS4suy+FKItQMPdIFfO9Kb7S08T9bJOlpJBrx9UboSUTHdZ7gJ5yzPI
8IgJ9seyKy2dnLcOeUOn+4N4CADWwiNfam7GPtMyiQGBTX3+4pGbpNLS85FkSRgzbVI1lShatnsE
Y1AEQr948v6+IgpQj6mmi5BxyCIPrU31aMuIQt3bw5NeIUJ8UawajsdKorm84tPJ6zmCfVNtMi88
+kXy9BAfU8kBrDPzk+5dMlKCoiNNBem6pBHJvBb8Ny0cG/N52OUTvdMbyfDFErcW2x/+l2rJLw6V
terFEce4igvKVUe+BO/GVXxVLUMVRtCZCFmDIcsobqOvTS/Lut7S3w4VmcSRIr6vx3ZljVgWZqTc
vpbFrLrQEabIr/BLeGMPMeR7bnusXhTy01Vdcmwj0yD/E0WkVN2OTVuXNC7Df9bfBQ7xdy+BcUv8
Zu6sruFaDxPmwlAB7LlM9GKP7Jv2SoHsCZr0ffVh2kvukwEudrv5KgmBq5/IqidcNjEuSLSgDU+g
0m6KDP9UypIf21NldIcyjK2aL1YM2A4VckdVoCeP5i3TuAu9O+XtJDqd2az2ZQKdkcMNg96rdPul
MBXMELLiAD46S2dJMT/SnW0NC0n4/rCEe60NSO/8qXwNRKyl9ArUouhSoe/Mt0oZLxl20RrWOaAS
gehGCWj+J70NFg0/48xLzY1Rc/f4krbZF8voRnuE4aRKOpSPh2wumhOvU6xj/X91S3AL/M5qteoa
IOQqJTdYHuhifqICMCDRmB3kUQyzxWYDLYJYItfy9ipHizmBTAiG/BNRl1OroU8h6lVWRG7mK7MK
8eJfUkjz2grywmYYCXqpS4rIZ9LQ4mRLSZNaHGneB1g5+/U1cBThStz7WyBoVjqTXe1iwGgAumud
lv4aSzuz/WBtWXhUZbIlW1bSVvIp8yqV1u2rFs3NDQHLM1b454ApdrjvzQUNh0y8xbOivtDM6xBp
CLq+pivAkhmTVmoTRDUmYYeVUBLC8q5ZWmk/bf6airV0vSfOK0rhYtfAdDCK1PY1PgaZNmpXQ6do
JrHqIltsdE/D1Dl0hilCUlc8KDHwUBdamUUedX/9bM1thqgT4m7OYR6gqMzEs03iF8MDZoX1USFE
YjVOJE3LB0jnpLKU5zbN/RW1GUHjAqQBOvaMIEt9raYXIY3xQFLnanPW3vh/zMCHX0yDM9YYb9o5
TcLTodMlfn1Rnxco78ptxklwtSrjaMIV61IW8rHET09ibLYBbItCX/v8CSNtKq+HNithmRoE+0GP
cmekD1OcxkNz1bpragBVj+kmThmDoqgKBM17Uh9IIe6dtVZ0CF/VxLSYxjASroyQROGrdKimJ2Bk
8kg6AW+NHa/aihekUqPhlkJ1rQ99rFajGQOsHC7MhxT3Q4lKklTgYBeMVC6NBAcqUZyeDV8mUjQp
6zcp+pja6gjh8cicECinPn1a6RABszZGPoUajHkgZ/HhESV/aqDjNrLw815EIK6OawCn4V6T8X19
wbvD/3D5EvYbKhSCveYipUj631ZJ/uzOq6H4q3utIc6Jci/dSSM/oTCggNBX83ysIDHwjJgXg6tJ
m1w3Mw8/jOy5VxJ1wW6ucK8EqXzsm94O0cvogKYZ/uHRXcyGSTQYYmKe6XZ2AXy3qiPYkiaNZMGS
51IhkPcGD8QSy1+YehZ7BUBQnDDXE2i9donkdxWDeQoK3bJVHjabkMa4QoNVlztviTyGqrId+W+y
YprPP59VVbnzruOvJtVdefllGRIenWUFS+VOM63Md7iccvmjY/ksSKIpNCVu8/UNeS80oO30qwLy
Z4wdrLe6jHC6v4u4F5FHy6bH2p7PlrEtJ7CLPgf40Q7oVN3jWk7ElpOBqO8WtnXqI3IS+aSwJEpi
PAkWpeIh6J07/x3E0n2Tm2mDK7id6OHMupED4hgkJ0FQ8tjt7lNNYvBKvuq5Aw7YasU1CpCOktSC
470L7F4fFEmqurl+ax/kkI4797Onygsk9wABuMHmVLyJ2KSPveeoWwNdJwvYxL29Gfop6QHbuYxr
jRgs5DEFdqZksnBBphOitXeU2vBycXzUPFSq23fqSJsTYUYbmOjCTUvEi7CR7takv3ovNwEOWsm8
mlhK9dVr5AywyQaBwFlFJSE6cVwQgCcSosofl5FJRpr8J31n4wJ/lq8zCYIUZ/RBAHeXlfJPZl5p
9TOYil+z7ELgd2+8D6B4Tbd+FJmdXJ/ZknxKEfVMKq+r2QN4C7vC5VZnjyF0DMNZ9o6Lk+mA7UIF
x4QEKrd+PrjJ/JKHoswaGWA1JEmc/vmi09pZoYM3P0T5NsoYvUX216mPq4HeN2C0oLAeM+OSd7cV
c5Bb86eFqD+mC+EBTJlQH0k+ylESDshMHy4svLFk8M6OLvVE11bGyoPqslJgHWnJlltRsUoWXqp0
4h+ZWv5fYTdUMxvNEnX1+TB+e5mj8xubTj7st8DVDHIfi0M6S7LKoLxs7xVtxftzPIb1fViuQGmy
r+HJYvHqrehHV7qb2fQ7xl+caIaa30NP/zZTrBtTCfDk3ktH8naKPxiiQhfbQJIuplA4TlMfq4Dw
4yCSQ85009uGWy5V9WgdHG59x0nMXPme1tzq1VXoQwvr1g4QhpCKSvdlWr/Ts5oo1/mzIM9wMOFa
MVntQXhixLBs8UQncqUVScXeIsx+jib1A9Gq8Jm9Jd7MDFfeuNrsJ9M7fnWbpbXQOkKX/FyJ+c+i
oeHCZLN1DOGJ78KM7P1dgeSjPfDLszcAU4741dd8Jmr0gO9pm8w0ifjtzzHFFeggbofxTcNVElx3
WFCx2cEFs5koO285pruYKQFqip4GBdv5t43OvwSAYmlDaxHZwY4Og5nGNrpQlDLjEkrqA3tGL50L
nMhLfnIhopjUtEv2dXNe0aeJ5zrkHKBuj2dDY0kjf+hu94YLhUOn2tfD2M20HbF9grySTpQeEC/K
QW0+XZ5qbu6/4WzOJd55ay5QWEgDQPC+wb3fPsmvhOijD0LMTg5Hh5guzxk83jUhpMBc7t9jZ97s
6u1X104cPzJybVo8yeyXInVGr0PDsVHcq0uqc/MGVv1YjpKbyq9xcgUbGGIth1rnavvl3fj6zOUL
C+3MR96boMWviB5d3PBxbCIn5baVHPQGzhvCfAvgzCxWVYkSAkCXg200j+0FOr6bxvS8YAMlCL+W
A5Lq7LS4jzjxwfb42HBql2NaPhjiuGTAmObGv4URPACt6tCHv/T21Dw+ASDG915dsrPecmlS+6le
Han+Hr04EQ1s3PvVyle0GZJYOBJiPcK5XCh6XXk9d70JPLnWD/+YgeTYDWvFNN44y/FTNdJ+5OVo
rjPHe3bnqzWZRbGgeJ8WY3tmIv9uvqdSofkKyGIEIxQTrTayw2PPUCWJ04GxFTVz0RBv89FwRwIe
Jb8zFuG6aZTev9t1JLInbVcg7cetaHp7pcXASFGfJMWxKCWJhCbbS54clh4oY0+KvAh6/fTEb1JM
xvVIVbO2I9XU5WgqO0ZGLy5U8FpcrrTIkwb1hXSHIU15FW75YojfIMLDi+8VXLKagZDALH8L/KLS
sZDynHhOIYj72/PUynQ2d8CBTZd0Y6A85P+eFp2w22THKeG8bXQ4QX7UdlzX1D9gCvPaEVaJ9ywP
eFJ0tKcYHDHvufneCPBmZajkzaDxK+0Vooi1Q/r7eFOyZ3t9QAiC79lhaW2pfQQzObwZdGNchPZs
lCUSXaswx0M9Zsoa/ZSAW0S0JBSB3T/dGIlLg0eoIlhxnz2UEfTesiAQ71TVpBKril6MfZdJysd8
NpktpsIdD40DKIeHkZ/MzPpGNn5x+wvhFFxRXwU3ZzZs5L7+m8Fi0FMemyeKNBkBSPcbv5EuOH5j
EE7naH3nhAZT0tdQGIqGvanSnmujqEuSbAuXHQM7EEk=
`protect end_protected
