`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LRH3VeVNPCPx5kjPDdumAP9ph74mfj6E1qr6pOPEh0cXuTuUHTpxnN4RFkIfdtXXl8JtaDrA4bvT
5KxbnqDtcQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D39QkgvBiYnuF/kQWUHq0iJle/uZu6Gy6/iwHytRC/3vPuMxQSD97VBfSWyMqlWIe6OIA57oMW94
7I3Og92/RIOA6pZuE53IJwl3I+6NfMj0LTfjwX+SNonFBbRQt3BMpDmlDZUSjUBJUu0wtdstMDwt
bLVXLoec0Ejup7oegXw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BZ5aW46zoFC5NlXSn9V5uIKlWyVdzlaz/9CONVK77p0Ot1vzw+D9tBMKSmHAvt/kbNqsyqnT78ht
D5ZtOoVP0mPoMm86mo7W3wOzUYJjQT1ygRklyXsqAdFPsa8lw36B+2+QGI0uLTRibIG4kqiHm8c3
tClJSAKUIcM3p+ca2D4e5dCIoGFin2B8y4BkQG24ANLxvH++NwbLIwa/Uy8uaqX8RbTDzCewgJjX
B/bYh3GGlVDSl0aSaoM/Ejy61LKNAFtOFHn+0XKCt0fl1N28ppi1OsbLNX/8R+i6fPtqiH2F07iq
6pZ17cof5/KirFjo0ZyxPAq5FDaJ4AKSVwJvJw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o3TQzkhL07HlfUJgRZ/TIy5XLcY5eSK6+OFHSbzW1tkgNbjyernKF0wl+RKEunM0TmEtmJnFQiq0
RdJeJDod84v3LE5U2yhIiT+RO6Q3tuX5vDgjk7UqemQLN5S4O7wEjr127CjODFhoTuEt+9tguVpJ
hcMJBYEt9uqIkZk4Q3YRLjs6Hhi9TIyFOM/EFvnmHUZXkLS6H+42zs6gptWT/9wGf0bS6wA2m9hB
lBFy09jDVpYehtDfucmLXcqi5lwiimDxgZsXn0WcRm2aB/Vg2F+3Q4UmwNndosv2+lpzmrE5Bka3
W61ShP2z6AOaJnl6sddj9GVPcl3Mfhxii7ELJg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ndmdp83hpFmk41t63yznjvkuqcacZHjLSSE2dHoQjuhXbQYwjsHKNTt7hZ5uiigCGhNeqg2OzsZa
u0xbo2DK/AZHSrzIfpsj0Cvl1rnW0mLKyPg7b8i7NajInBrSOnVvpxUQKlV3CyOzrbBcqmQfl4cQ
oCzJqhz6k/I/DjFmJVEmpHzSxy+TIsdrVTKx7aeAcVVPjQ2xNwBZBup21IsoorO5kaqZPPo3/8KA
B9S8jMFqmA4OeWdbZxGt2RSVN03O8NBS6GGAPTAQ4zQrVCzhpYmCzB0mfgqfKE0kWPqrJbQjGl8Z
jEIg6dgKJzAT0rIiSzlEqcIDYvzi/CrhfRO2dw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SC9At1KBitnCk2bc1BghVxoXP5FU3CiulVRi+L64OgXIyQYf5M3vsCpq/zuJzx1xsLU7JisrGjQ8
Wozjxf2no2XOg5lj4b0B9Eh1L2h1TjVUQ17/EcAzIIzNTfXQZGGH8jAQQF7hs7vKiHTe+4MFBFU6
4RWD0wr71ObF5Q5ElaY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LGD77DZBLmtrJazVimqtbkvF3IezFTo669T6SL0Fcq4OqO1/5MVROwZYgO3CZX+CdQXaXgQW4t59
oVlwYpDkQ1ma1SaBQKkON71Z6tlMY6xDkbTYhi061pVSvSs1gbkRbId3JsLP6H7iZ3RAZxJOIYiN
Rqll+D1LB2HCefEZBKP93uZMtqHtSGoPbSufO2Ivp/jEYLHuorjqqsGDN/JGYJPybaIF09G+QrTI
DqIznmACg6vg4xxt3D5iuJvSMR8OIpxfLZDaEq8NtvZHchR1joETfH/qR19gDSLNKgZtlHo+g54Z
P2PHO/Ep+ZqrOYQqEPLe9yBwB1M6rv7cS4gFng==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296352)
`protect data_block
BUzfmwXZaeQ/5VF4a+jeRuH+2/DUhZ4Hm51VxBS/bUYtPbWo5EXtFMCJI8kZxNZzo/kekMtjFU6Z
CfDlu/sIrwS8dtsLrOwbXxZJKr8oCmNN73ZjQ6d0gm6YdSmUYjMAOh+UINyuIZZ22025KXOGNdKu
IImcYAeHsVZZNxKfCXF3QgQx1w62vPBSmWWE6QxPMNP6aN+1OxD45LOz6ugpY9BOc6Z3oJOZJtyb
HzuF5nCf2t+k433PEwDTiGY9l/J8D9IG47iGBeK8a+wfBr6co2aruJvxkS3s+AWD2z1+lPIMsOgY
lt3p1uGTi5StcPpzT7fCRz+PbSH2aSl5VVbEm+PR+k1hzFd+lNRTWKKVKqVo33R8qAmeOxL4x8F5
fIukYp+gIf+8E25KZTuwMskZE9LuVVwgJ0s6TGk79AeKf+AvI4ptw9xjTZ5ibydsuOOk2Fq5srXt
qUUkTwN0OHkbauBYTlhx5QZDGlwqphQRUNaUiW/GwPw/AGp7MbHuaOuihCSi/v1zXTMe55aKnVpQ
gVB6lT1acegsjgBiy0R0AB+ygZrez1Tkd66wsyW3DLBaPxRvoedLMdvqieilBlorqrB7sIEr7aoY
8PYnxh4YCztxM+LtMfF6g8DfuScc4yRgII89IoMblSWPVGhkk904YvWgr4LK6e661yppcJdmdF4S
U19CZFPoWQdv3/gOAoUppwUCDQ5pF1+PBqPWxnwaCpnV2PVXzGQ5Uaim4FXNwoTdhW8ZkxJYew53
E6UJQIvvO3KwVYvA+sadzgTwmW6RWYGZC8GU0XImZWf5hMYgjhJrDuOa+gymO6rI7PEryIts1FWk
/5wlRQ/NJrJLjRYACgVKYgyw0C/BJ/2zlecs7Kw2euSJ0873Ohoq1GWsmuq7ghWdHwVYnXsMbog9
bKH+oo6p7Lp5bDFQTmOYtKk40vVuzvZecuw5vb/+oIqE6BTuAWN3hb+5cg0vnoTnPUfvo2mIMzfq
Sb27vF7GaDgTJ8/igY5GCAkYLSY5rXRyKAF+bYRqbTpDwCV0d6LZE6mk/7XrSVjiYBGxoasfYnPU
xzMFCv/mmdmZz8AIGxFyJ4zAlVnBN8ItwowWoDe65IS93CPvjx2wagV4xt09l0DjZQX3loQEIC8Z
HFo555JwQjc4Ra5bvSHhU9rQjUrmGk4IrQ0HgCMGiNSVJ8EqAe01DrY0rUnVLX6RO28ZBdU9jL4j
5bZEz2ne9RxSFKLcVINWJzrdfrcezttC2REtlW0FHBugTCKEnpZoHICg4lW7zKjpMPIWsXF/wsAr
5LKKs97jtDsjj8MnNS9B796kE3hOEZdqqhGmnzzC0fYm2JvYwl0r8kYR+7KNR6tydraWMg2FuzL8
r+kD+RnMlL1tcc4JiUuYGDwuSkOFOLFZ2HhSwDla+kjYLohGw61Do1sgzt8MPb2PZ9rULGGhbc1H
SAjWBJjzGi7MgtR5ROuxrg/Htu9s7RaxUg86/0eOkb3q1/jmbV2txTPp5SuMthBn0r8lv5QgcXSJ
1EVqwOWLC9C6ZSA00VgZfklAnRoFbie0MOlNRxKlwN9w5BrrgVsdXuN7KWFKcPnXOdA8YTYDJAwd
RnEvqoGF/+CjM8sKG0wKn/Q/K+Ah1+QPtIw14ZjM5mQftFn0oc9nBpPo33/1Em6+2hw6+bVyotSI
ilWOqpgYIfzgeiaoJynWNCzKIebHMU/GcxneB1Ab78dwxMujLFGEOj9bfyGhZwbdOj+/QL1TGAx7
1DT3ZUysVu05uZfLS/6Fb42sA1Xhcl2Q7a1BWsj/tEWP102LAqgjZHWdZ6eFV1IIvcXUWLBtKgUF
Tm2erT9vy7bWXza6wLXRJd14k+sits0T1pIwkIXuRNVc5fwLYpr7oR0yxfqm6m7vnQrH6zXXLJ8L
Idrtz6grtWc+ZZ/3ZJqUCuZ0wPk3hCB1dyVBOdCK5y7upGQt9xirRPW+yF/dhaAv8v5wJed9hH6o
/Bw2WyyXwthmbsje3SCHwZFFPb9H3DXTlLVUgIEgDPaQqDd7y9lrU+IV48BlXG2sZh4EmeKoRY9S
I0y/1Kek9doFkUdfZiW9Zo6cWXAb1frImTAdouDc6G8GTFdUAelNlPNC9s9jQfJNfJ+wREN2UOXP
OQ86IkYglFRXblfM3NgePzgJa0sd/khnCdF73tMMmHCcoSMQ+wMo3bXinvwnt81KCZEmwxHqmuKa
oLTGIpwnedy8vK0IsuSa52xho4o2frpwhSyHg71fmxApXZfBwd+dk+0AbxZZ4qQZtNRhdSdUXlPM
QfJkKl53iIiqnHINmWNEHXFT3gdjkDzLZLSteskiU6YL7RoVh2LAhf+hlbDtabRUFIeyFMwZK5KQ
oiNtcGr69tjXeGP3R9wKvM0maugYK5vX/uSu7NZr447xvVLdEjhuwbwtzJRLfV8bmpsb3ueKM6eD
6Ombs8HOHe459jQ6ItbFF6iMymwXgbb9dGkA/6FeVOBUKhPWkNo/dMj9DQvUtmb5x5FuKwmlphHs
R47TPTeMtVknPJcF3tcJyduNwLIbSeev2TRdlgh4gU7HxpSRtq1m+tW9kbrPnporLJQ1mdnKzNT5
wubWTKiiRAv/yxZyV2Qwvgj6GJ6YqDQlsnrvxsaKrV+viUE9OdT0xcKbsO9wNTHrSptVuk/Soo8z
eejcgewhJN+z7H0dTkrWZmCb7IuP58X49SMjXpVKERhNHdWwkhgUCJVDpyJNfDFw3qE7EsijTtm5
ULtLZfaBZtviYr7k/8YOOUbZ8znSkGUL14qShC0PDNJUW6FRBQH41StE1y9yn3lteQYJhxkuFwvm
ue9kCN0jzakF/JILsm1kapjp3jgC4PCkLt5FUVVM5qVUaeKUrwbSiE6YQxgzmQn52bnSDNOC1YjV
e+IqKHpPGhziQe24oglyYgSck8I/K3AI9JSPYOCWh6PfC0C2U8PUHeMQvzivYBXg7Jnkxryj0AzR
5qGxdomPdUO013rpy4NGiCHQHA7GwJFlwwktctfFOUGCS7R/8jra2HN28ufGK0OEROfLYCJmTFkk
2ym4NNUUAex6RuPDWAG9QWNYmBkK7q/plxFbJGEvDj6djoW8RDTmHwQKipMomT90cT2UEb/EEiEv
mqLmb94f5WgTPKsrb+BcHcXooKG0ATpAibwHpimAuuWa4Lc+wJ5qjVg0aAaJvDUR7OEnxs4f3eU9
pRUrak/IYmn96lCUcURUVFse/GNsG8CLU1Txg5DzQn9aiTA0itRx0itakqCkJtmwBEkYSNHDEUv+
H/6MSwFnl4BthihlZjQZXQ3yVqW+TdJ1vIMNKijVvj+Y2xn36gUeJPKmRPBWQUxwru9vebE/qf+J
nVv3C3iwONTO8fJlr+uU0o3X36NfPGYV6ExzPXJOqwejpdnpfjtMIvCpEdoPZytlsdjhTO/MqrBW
ccecY0s7IACB91v6q1eVzPFw+yg5op/mUYZUkzaJbYKmzqCtlD/5UQ9EVQrAl+RtNOwOpc0i/liX
PtIRfZQ74XNbqmOtOecpfXqU6ofQ60DJTaiCdijV3aP2sRy5SOQYaTiSyCArHGQZ8I0YwPaJqIEm
Yiz2zpcajnQ8P17eHF06SrSV6GQ5nqgUkfGkMNfAmOePMT0cRixV1KTxgLSponCgwdJ3pLmB/tUd
2DpINs/1nBnfynctl7hRSpTExQrbWbQyMN4qvCJ1WBdGzRkOXLNFtGT2nwsIqdQWMNycEpP+6rzN
oxC27tqXw3Od2adgr5by6O3reBV7MyuRYJZsT7DFWtgvZnYrB40R+Mk3QSXTY8Tk7T9T//CZLz4I
C+eCM0Rw3uyk9VG4RqCDgQohsTGDv+DujxKCov3JLQEJFheyplpKsdmtK0pLVpeuekFdoyS4w9sb
Y2Lac3bVWttkEwGRD5qRAjY5iDJ6PYPtAJe61FmOuS2YjCe8LKWKJl57jo0IhDMjnPoFFgYOJits
iDrtPRYR9Ik0w0F47gCgXeWL30PsHiYr+ZDIe4+yQbaQZpQ/TXJBaobDrzerXmPAhi4J9Gpa5iSa
gf/SLEkcoqi7mgEPZBRtxjnskeQBjmxsUree8JxmfK6kvuDJc/IpYnRpCNGLJZcoywy+XUp/QKEb
Ltmd8aIfFcYR1aDDOh60DyUp1RDFW1Jx+Z5W6XMhPPlvIissUv8kPNekYGmZgRPLn8uqnu4EWP/R
DSYY4OKd3EkA4N1+DWzGSYE5AHYWveu0VmL+qQQvR4/bf+ZQLE5j8VK2OucfkOqeohhiqyuKIXWw
aVwaXBDimWUdWSbQT2GUMWjcqRrr9SMLiCL2WuxW6WQ7jFyKZNt27hqR0BJ3xcyjDAHWyov6VQzq
FBsJ3sTF/Egh9DW6D7OIbzM1AIEXX5rshl9OPush+FB/ixc5NpQUJ7ReqgVRYgwwbOCDK3AVJDPL
n1YT75OwQK/AOiu8gC3IVmXUUZ81CLyW3iWgtA/IOwlKOCwZ/9TfzGQ+X6ZFz/lfcxD9S4JVxrgY
D35+g1wOhZRdNGonW4VpyM3TZbu45v0llRkh3WkBbq5/Z+Zqc5CAwQB76HKF4fg3U9ILwU/CGdYy
J21gPcMlJWD3iv8yuJOCCfK0AFXbsQffxyShvXtshB4XWO5MoGGtbpfsKeVDtYNFMHwmBbbp6o+m
iZ+lnqRiAQYkJ2GEH1RdGO5LldYFHU6uhPDW4NWi4ZuEx3g2Ga1bwR5nQFhQmDUqLbSYjod1SJ5t
7hoy9r08f/kDLnpSPDaahg8sC7Vwyn092ddzpMAbNrSdcI/kxZ+70OW/PvXGHhLwqqJL/SgxyXVU
LtfgEV+9Ip9CjtmeZwrzZT7+K/aV3c/GBDUUpW2m4ZXRAAKMh1mcZtv6k9Hc5clveGszu77S8NVa
+O3tkAqeYnjHDalXlRM49JRMiIme6C/F0/2V0ISQzlXH4he8bEfU+15aEVlbcGVdrkZQy7PbhHwQ
zOsC2XtIB3iQCyhNK4+adk6urJNBV8wrQGcq/hz1HabpMTE9sDwq/6uthhsuzqqM5arOXU8uKm2x
cx/EekHKY6nBCAM/yAlP3zuMOdMMSjOoGrCvPsMDYqiiumcq0jdtHfM5cvIjCQmoRMdRR5DXYKng
DQIaYEE6u3BFGanBt9/E4H35Px5aenG2w+ZnGdATK0WiLeAbHjf5sC2wDuzwxPfVNOAPbBWtMZyZ
0ky1goZied8uz0ikDJLSm9krJY+vXe8zxCLU9Way7SOF089ODqTmuGxXgMBnQhAag3BttrXrhGau
j6Lu0dCblp1cCP8/1ZdVzwW8aHEGnCOclI6ANMnL7HHDpJTOdtzOG2ZGb+K+XkDEuBleLH0OdAH/
YYJwlqujXIJrwOBqVrarQsWFNmxnaZM3imt14/9RrEzjEWXf0dJx0XpjA/wlV2bn/iYUMftLk7eN
iEHPTtYbmG4gT2DKrMcTN3MxztPsYvVUAT/+Vz6QrrBfZYAyQQ7qXBATV9Rag60ABKKTFebJuzTC
nOEDnKjk3ZVaYFpTCl7/8oSvNuHgddJNHFupYj04COcgNER47usLobBO9+mI8PbxYLgYuBjPhnSO
IoUPqeqa9OWtSXs2ZgvCJZClhIrU2+9AUrf3fHq0flooV2fjTDehduvlfp1tGODtQXJl66TJV1PA
ALckkZrs52UjrmIFIF9+4tApOCn5JAeLyGHmeCZSM4danTdUu0S1pGtKlFkuptJcpxS7DU+iNGtN
A0CqG0PCQ298FB2nlNgEppHXBESzTBnGNTXsCIq5JbTVoe+wCt/R4cjj92IibUgo2yBo6n7f44Fc
NMuX5g7vknCOI/llaaAxACg0aVx8z4b88MeF0FFpOy9cT9jmacs5B32iQ5/g8N6jv4ln04iUWYoD
6wPIKEk1ZijSyOMosZR4rtBcOohbCXrwegvQeCbIglT5sPBdIjZeBRi+PdQ/CfEVXoSTkAG4iPfg
73nVVOBAbXE0atXuoRDFY1kRtHa7dbFXTRd7yMLCwU7wcIeMP37pLr1dd15QuzUeY48KEGITmlDg
BtW+JW43S1a5VHFjtTubKieCkdYeAyItXPdkY+Dua8X9dyX4T9N3euigRRflUI2FcVSsrX/76YNO
gggfzJtZ8u9oakmJ2I3SNa0nxBEOJeTmHbn0KcfH6DCo6nXTNF2gdnk8/Yt6AZvnP3vYgZ1wgk8D
VrTCOqSKwmWrdiyVHFgyzq3MS+kln4WYeXiJ+G0prH4oyMfTua1Ou9S8sC0FG3qzVcMqfwE27Ky8
cX+uGlpwWFrVlnmgtmY/tG6OWsS6pYGXjJoRft3tPjDAo+XqHJ/zm4xW5p+D78s24cZ5ln0C5ncR
8p97/QEUJXAcKV2Ow4feUVhtqzurra7CzsJHgyt1a0JI5nfNgBfDmW7YF0WPh6mW+pzyxaAUTgYv
yc1f9dniblzyjZhf8iq/yo9cCZOhS7ezNWpjS3cy5jzQOBN+8QTJb9wFpo1A7lwWWB1wDWGrsM/u
iuEMgRlOa+TKP+UelPt2ADj9umqgDEuQWu07aRZMpAd4r4RaxkLmv+mJxaHdZ3UeRjT9pD/R6DeT
LbpmNDToPDmPYdnoZlqIVSZH4xG+UStvpulVrLx4WgdemPV5ZdMsziPcYZawRECOoiHsAt59NS5+
wc+OZWHgIU6o3GYMR3dt1OorwBwP5Kr66mc7SPIDeVC1TcgVT5YiKHDNTbNBjUGmvp+399B4K6Zy
j11yYfJ5H007gxtau/mrAywycr1I5n/7KG+Vrh0Z8wJOaRYyIOsQugUgZT/kyipLN9GkDBxG4eYb
NjJmZtZXt7FiRbAQrhRKufI/gM8NJbt0iy4na9OBYlkICK+cakIyZSrwjWS0dD8CLt4lYzE8bwiz
UKYQXmQIkGjuxnXuJIX00RyZrzLYG9VkpcWpDjhJ1d653btrAbp420UgOkdoCUAV3BFohGnuzIGC
zh8PhnkZ812Hza2/HpTf1mdt0JPw5BkrCn+Z2w6JQ0a8GriuV8Kd/7jn/C4EeAJVhLjxZuBQ9oHO
92nlkG+5n+u0+KyYusrIGGeoZ4vi3DNE4VthYY3snLAlY2a+zQ4Z0w1m0TAh34NpBPCEO5Gjmx6e
oy/WhNLY7USsHTtZAu6m+vU8VuZXbOmMczCvVC3tNqqU4YolvWyqTuQhh6+tR2xc6npm4i/DNKf1
FdNQa8ismwLRHSmr2vbZPdZ/17TjbBlMYypLexQslR3XHgIecsymWuWNFcAkc+8FH0MA3N91Bedz
E5ZzB+IkRdqDSbMnCE8YhHeSH3pJIQsf5WRlbFWly9wWnUPX4zqVYMBbM9nMnHzjBLjT2/TRUnBi
zPusPxvmtNZ104CumY6umKY+bu/kRSw5QhhSDd1PAC2Sp0oY34aYPcdiV11rlZZAkHlDNgtPOHtE
FOw94UOIrhDc6YMgg+j/onLJbRZc6Nco63TOp3Hn3/0vdZv7teFB0gvvF93rYcj4u8c4hSBmVhvS
19Fq8HxkZ2eOASmYAQTzoZljBFa22i7XeHPfgoF5eONAwTBeSgbBJo00ST29a3MRI87WPIQvD5A2
saUSn3ljEu+CB8dEHvgYVAXR7oyWvUXkbU7tNrJPferE5UxfC8QTscdLrKa6fjoPn0K5PnrF4ElG
HHImT3iHTxI6/T4QzJ1wQZyoltfsasiDZIE/z19n9BPl9L55zEaLWiy4S8hR9oMMplv7HS9FpJf9
kKH9WfJZs8O4hDRI0ZgVGkwBaQ9OVodiayAefvNkDZuXbdkV04UZyuzkZChcBkefgUpfdAqtRbdx
71qes6Weun6D07eumL+rBCArPAgxRqsgouzvz1e2hUswq3BBmM7sYRdjoo6gXaowJGArVdiV3IFP
s6gOFRyEScAd6jIv39s+m+OHLTWikwSIHLyFGzIybRjO6w9h2ZPJ+Nb65V2Hxl8JVvyHDES/yhIy
m7pbAa/jjizfcl6i68rgsc/HCLg7DCREZfT3BoSl31JM9vfxwF9AcW3fz86+bXF7UZ+s3UwZSF/O
1VXrVoUcgkONnMGIuWQ00Ec2MGxUmWU7yikBR5M+ePEYKN3YpJj5tnldH7rTOQy+PrSfzCmVkfcW
PVmQEiLxPho9iFN4/kpZQEYavOZoa2Wb8pTvfojkPDyB5pCIDv9VD6qB4xFAjffGi2wsm7NsFlAa
x7HSZ8cIZ3ixhI3XnvYIjm1yY1wSq6jjL0GqmniYZewWTsW0CuIgd0Wg4+4aPtltx4c4uOk/BnaS
1+rp8QmVEcmjFp+/sf5qV/Vk84ILXDoZ7SuWRAdtQ2Pr54Kwa+uGq58k5JXCz0DFL92c8JryZPJj
pg/vKyHZrLroBZqvICy8aQq0Vse4LddJxjSbKO/9Y73ssRmmqa+iOdlRys7uHz9v5NPjnDuXUE4C
jtX4qXGiz4TzhxQ5VyyMLb65vIQPHC9I3tI7Oh4s8ASIfaNtqNuvB24KqcNJGpAHcKmDu4zuiYmk
borik6+jK2Wy8dAcbYWJp/WOf4KwQaBMGWFMDV+K3TuobdO1hUDKPfwLLVMFbdZTSChKoZIybd0W
0DJopmkHsVqUuJs7VsEPyec2hGPs8WExr6WodlEZrTmV4orfVbE+IZk3sF725I6qGJhqWZMmiEnr
KMK0inBQYvhnh2V1C+ldgaBJSxl2/cpjqNy734tcEXbugHtMUdMBMZJWdoGI4bK+86CCVOEmJCq4
znarVU5b7YKVUl7HBJmy4I17Y37JhyROlA2g422sQKw028lgmtdwSFDKH/0NG15vsMaqU6Z9R1po
HaNtE3a4y1NPWVJp2F8POUch7qNCtiP5Bc5dSKJuFkd+THqu67DFKbAbmsYB+pePktATBU8GLfXs
MjmTUbc6ztaGdtS85qeEqttHnbHfg8GHXuRuuEFw32zrYycEceqwHfffje2U8iIi/DkXDdoSH8Wq
ZNNcbm5ejInzQ/vI35Yw9slQhgqwN87NF3IscMtBPVovLlOy2Wc2hjk58TZlshAJSaWAm9QE0c2W
hQnr3A7skBlAGU9EoziVFrWhQu2wzl+0XVuaA3XOeVsMuNJZW726jfqHiZhlpzM8QFcUERS+Nqsk
LRm/Gtr2zYqBbGFI0KBR4TNchJpXHjUANb8n76T8itOPXojxzJo4k5FPg+EGm9Oi0dS2oYLloDEg
Qvp6u//dPdLFbqAMZb1y7QZByxC9JqlkZfKClRUUyG8pyQExkhDo3z88G6nOySafZWpn+8PBi/mN
6Snor3Gq9SiOL2lm2kRaHWbN8xl/wGlJgYab8VAYaEyad/7+sWRw97tVR+L/XhIQ2A+UfPJVF3wg
hoUjoFM2piWfz6AizFYKi7PkdSg6vC1riAOaDnRn+/3b7xmwE2sBxgr3UsLbY4g1nvbvao7m+Jv/
nqdWQgB8iAyfzkUYJ+Gr7lf4sQRZ/naxt1NNPeLm7W3tSD5bRrXjgZf23K8pJBqSFlSLMPl1AVaS
9ca3g1/v8hzYCH4FqFxUXqwWp97E/2bsTI+OT/039CmGQHt6PtEOtd+pH60XSZDBcZ8+evWmXWvo
hs6vmS3bxoD4i3nlK6KEtLoMDJgEmVuNLDTR956XfH9zSHbEigqRm5duHhCaG1vp5Glq6dYXoZxw
wNd5/0t95Pw91v4HIv8fEW0oyBHy4rtZ4aQMb90Q+hRV38SN6kA2ZNgxgxwuMySvTFKZhtLcIojj
AmnsyZ1iGNUr//BtGkQ1bxtHRlQJdIFqJp/lh6TC1/JucW83nHPmG/8Cy4XAM5KMZHEc+7PntOLZ
KAu/5uQnb9HmRelB4Gjro/3lW5o2AVsY+sHKx/QiQpohWE13vJJwhZ7RoziEe+nD+VPLXw2YWpQY
MGc8w0uDENnl5001zgM/NS1KYmXIH+7D1mklqvDyR95RQXADC/Wkn9ic/ZOsTMdrCbzilWM5iCZj
D6GZRhwZQqmnMkm4R9MEapExqGuOvj5GtiDtHFyvx7orCOVchjQ90uSvl40biU6e2/e0gjenSyeM
QZkbDwkVzTNloHKWWlaeQz4gFb0SxAwhKe8IQqc+AvBb4I3wxsxl3pGONv+oVplrjrOOCvH2SHEO
MJCGg/pA+r072/jExl6pAYOVWAdxHosYYDo8zNGxBGQirc6Sy/uipWiT83ftTgvW1uT+jNOH6K/K
7/Laj0xc7ghe+whgyLBgl90LJz+aZSYQI/h+ye55iUFpCf+ciRNUPzMe+VMTXMXKVoGbWbHqCMkd
Qc6cKatpXH8zFRAMP+gIF09SwbidGXSvGP5RyTdce6Zr+4ewFRJEbcLYN4XgFHCQajNoPvCp1cVD
c+WkF3IUcYGTUKkB4BIwMQEioykPwBWdbyLnkf3WPYin3/hrpdUrlJ8DX5f2Q7J0RCP+jFaoslIH
wrjUxzUSsf1VCjjVbVdVWug63nBo+jAvfE1HFfVoRkr4wm5mYK0r2JwdKtF8K9Q8u9FCucK5IU3h
NmpSPVLcR6Uw+9bIBSMKzTUKcnysFu/1kDF8Te6M4swoRsxZigg0hdb44OJOYN4rdu0+n7v+TiTs
GZHyl0Xk8PdJAidHLdcL28ArynhbJkJW7J1PJSSg0kyoYFbWm8FYJT3HVlxVW4fwunF4f977n/MX
wn5cD3tB8KPZ+7HR5Iyqgj1iMy5sc2uboXzHY+fTiLu3ndC+vqnACbJ2q7I7lkIinTZafZYlswx2
yw0CFhqxAcebdq7AIqQ+EDFOKzQmU+ok2YRKuXfgv82fBbwjtk8S0VdgfIDSFqrxgTvcM8OX3ogF
mI59p6UBUKqpfHbNnassrGInNE49c6A6/cWLdZq7McCtdp3xHV74yV0iHM430she/nztlrxrsxsl
MFjCpy/9ll3mtogDUdyIqz4qPl2MHO0/wDSYYXwGMCa4JSqu3szV6UnN3uCIZw3UYyRYqs+BCpxJ
DPHmNClNxkwaSntZrkEeR19XeYWX0xDNXd37nXs3BVLcgiZJZplAl1aH2+DkCkrMsjTtZrcXcppA
MHablHWtLZaD90qAdxhP8MrMJjQXvndyEuc9wIJWBBMq/OVLc+ol2rp5xlp/HBUteGUwOnG7zvLQ
TD090aENY8mfU247OF///MlZExpqKh9JXZbDdHl0F4Ie45c7KTg739Imwmfm7Q8xDZu+GAqsFzLu
/567j2Ju4TNtTvrtQo373tdSK9TmA6K49kepJ5IT5nFnw5NTLA+L3Eiho5VuCTpKOoJ++MQe0xbX
IAA+eqvBK4tZFgrfHznwiV6tSkR5QHT0Cvyk/VYAZ0KXA44dPspFCqY5evlTltdsZkyisxSNHTG9
KS4mdoM1xmGdylbv00fhasrfGDD/7LnVtVr1H2CNb36srjEqXn7kQqvU1ZlnSJfm6G/B9dgKzB1P
xtBfZyqA/PoG8/aueul9bOx4C24aICJZ3kY7tRIcdMk6YLcZOWs/H2fz010Sr/3n1TmsRAzMKhuL
4RyVdLd0EF5uOSM60bMoXI7uGhSSuQhfA8KUyJZQ+HE0QdZqpTtAgECGSXq8cWPoBec+er3AJVS7
QEbtGI7wrEys9qS0UpM5P5nF2E7/reWQl9T5f+AoZlakd5coR1PcvE9jWEpziBV/OMaaqvZtNox/
YtNSB6Q0shKxtckx9kZhyOgd7oM6+OIl0Xj7WFweRNjsnjM3/zRrJgvelamH7vk72XJW2xiZC4/E
saaR/wpIkbnijCtVRKfEy8sJiUBoxAQk70ft93U2QZXKVlUNugjgQUrY3xVGkJ95bGQLqKYZDRt+
wMq10o9ZLKg7quWNk2iafdOO3WO3WSh8GI7BmuzEhUh6PS7Gdt7VkgEX8+45+M3RMrA6LvsUn1gj
wm9TEA1y70Toa3zzp8L75BN5DjStwEl9G0RSD5c6lrPmLupwxYOKVfycUQ1CL+NWfZQInRkYqLjD
ZoTgPPletqVtkM6tbtpKlAoXVcqq7+/nLljTf5UNwTm5mYRWLDqfGaV9VdP1ySvX4AXBHh5L3Ye3
H+3CGB8FznqCKr7ePXjt64JFoMh3kfeXZSB0zZ991Yt/V9Z4RvJH8ySIeb7+5M8alCLmpRT/IBog
JsqRWvQvTD51ZyqzEH8+5+ck5MReWWwMc3L1oPc/7d4yQO1D/JCeksnYLCjlKX45EjRTPPylR242
ieSf1XIu5zTCkuEPTU7oJyTIjN5Nsl987uoIg5es9EZUWNE50inv8uGbZiVauWHKz8XzRseCIa8Y
F/mBFDRHP1cubs3Z1osUbwbJnfIyjQP2RVGGKIxL8fGi9KOprVC/7GkDB49lCL+nwUj92jqy8DEQ
/6Y7R4+7cLD0M1SYyYcqVTj0eu2v7eWJQmM/7xgs3UgpCoOZmyX4RXwRPuykcpzT1h/EFhXLWngp
pU+oAGECkrwtyX2ij/y6PyJwGsSnsjyOb7T9hsEF0VWArEzXrT/A9Oj8yU4uXu89vx3ejZ3TQqRK
nHnRMCpLQJkkX5qgvpzgebTMBz6bIYLB3f7i+rOmOeZqYnMygtGyq5lh8eJTI/xwlIbDC+wRQUiM
RhKoYx6noTh3ihKpuV08x6WJNS/FsGed4nrA2PwTGO0QOUQ/u5SAR8/NvHHclVmbqhaZx+OR/oTJ
yUAQiOzq6tJtanqOqjedP/8SpmxsJJvbNFGS/7USY4EzzXPLjSFf8DRUptzk/NJ3ugX+s0wLRnGR
GdEQ2dVcrymDoOWpcv42BmHk3Fej2Ks7yXNCp8x6oMZW2gtZazguZ7OonGYD9+m6lIsPRKkXEu15
FQr4K5qsWT6RD67nqruHQReiRGRIJddpMX3OyDoI41GK6twSchTbv8lZeHqkTwFg9xZvh9n+5eJ2
NrzXQLU2P5oS4WgdSPDNhgMi7ZFqfKIu+HR79MueRb3+aywK5mOUMmQUfFos+1TfiZUmkodp8OlF
Au6i1Fl1Nnh8GHtrrXSd9ClvEj6u5W2p+SDWyvdnaGfP7aB9mvS+6t0BL/bOthmFoAt+vzQ9O8QA
5eXhxlZ9FbBCc+oifmm9iZZlOnx6qgR0ggT1rtERupq0WP6FvmBcKB4Acri6E/UkQkqQ8WyW/aRD
usPBdrwZMHO+GCY5ENeXh8jtqxT1AQFiXKlS/w0KCDjoG4Yp5ZHF5IatkbxDHl8N5+zfiy3qxy6o
XCHYfXMw39cT92diEgi4RVRqPqVhYUhedbEmFSkhtuGi6WNPXCoeGokjqhKLM6jI6MZtCkGtee5k
CqeIon5E6IwMUhlxT4cLyyL69KxWTfBHgve8VZJd16HuwWtrlHgpS3y5UgJwgnfHU17CVBouKZJN
x1oGW/7PbmJOeBquvaP0+qADtGTAfqtuNlLSEgIHR54twtOuyu/gBOVU2ooPAp1PeiVKRWjz5HfQ
QwGvmJWIKtbDMo9WqX54LlepppNhjGbOCFfA+OJFgfRx6hRiFNbDHx/yzGGcftDRIXDQCgTzQe68
7z8Rk+TRoIRXba/NHudv0Lg4oeh0Os2OoxoXo4ws38AGZT4cTYlhccjjU6JelqFAoy8xdM8jYdPx
ujVAz7a4VTgEVnBGKe2ouS/C5zrBKkyaPDOkEVCvA4mq/easevC2Ge45nkHjEPa/nebdSvRA2Hhc
YspJ3fJSjU84KCutdXTfcR0lhbLcx/o8zYxrWvJNPayPXFUulEtR737smJ+nklWcZJ5gsMpsrw42
c2Ok6hTV21UtqharvtH3wJGDJ8Sn+HEqKzzRyA9PwZxM3VHEfFOPWOm59pZQqcWsrFsllMQrJxu7
Qi/FD2ixqv9UeGHH1qUXnywFR4ouWjF3CZRlsv1ChCR+uCC3kedgpBqHe4X1uECZxJ5twBZPXM2m
/X5CC265INBhlDg/5l8/gJs+VgUH29cHPBU0NKwExCVuSIQN67RWy2Wm0GGen2rTCpkkbQt0AOxo
qHp07a/f3A+sIzOj1YJHxaGf2wBUf6FtXgHLL1ZPlIVzzCOOoqCcnDCm8ZoJp7jD9quAYG5eR5QC
0igMBSoJvmGFf+E0DEehW48OF1OnJr2dHN3IwnvwOFs5Z4Q2d9ylFi+UX+HmEdKUsZOmN3BYxbyH
EdLumGWTZFlWae4r5MCiuKjuHZCWz7nLvSm0QaHCF8Uj81szLMpjN+hK6JwrLgP9mGGPS5DH0aRu
OaeSk00JIEzXpve9Yak2BVOlHvZMOI2y26epgiSdeK417T45KuOT0sX98vIzlKcvSqvYjV+LglRD
m5jFYzryTHy9PhkbXtlN3vk7X4QLIuXl1w/fTmQi0/08A/ITViff3AWxM3EfiZwO9HP0+M+EYFqQ
hyRSpEmnRxqgb8vBdh1Q6NqdAtiXJw91xfY2tB69cZegMx6PJaq2abkVyvau4Z6YtIXkBJogUG1h
JFEIr2JqLWyjEHKZEqMEdjdeHmbDBlBPqK9OF6GKiLhOUDckhLqCre2yN1IQcCMoW3TE/sC7oRVO
NLOJFQeDn2+rkNKjhmT6pXBMqFkUE3zbb6NmJdzvrqOyHVcwLBptKhZyAgnsDK4Km13muMEwj4zT
ckXBbHr/fAAz/4q3/UapIRZBQJeg3ncPe371r/SECHWY7wFXnv/SaxS1Azhwjz/NhRZ5N6LearMV
kW77G1RfRb/ZMnjUIyBvbHwesIdN5QRXDCyUxglspbRVX6HxGOFwnu6RVHjGLJdnpSUIQNbG/137
RuiqazILMASl7DV+FKv3elNUID4ueJMevJmywm2fIyJ7dcrE3vONniIUq+tMliterPmfxgl34S3J
xB1EQ1JBeczwlA7De6k6SqaWFqyUcRKP1H1raCogwRnwTJMY9DB2YriN0X2KyVhhnkTcIXqokoWO
/Yqev79xC08c/4auJKu3sfEXPiLR1Tw6sJVFnF0zrbCDNOTE06B6T298QCVSBo9n4bNGRGx4382a
5cGNtOPdnTnDsjHJSPKR+3Y03PbHEoeZB0ebWYtMo2dCwY2lItMbImcJlrtfJ6tNPMieHN38iDKO
3X4EA1UzTpTxnTidakw7jWoGiObsQYxTSz1mi9xdJxMnPaX1f51Km4XLFSRoNAnk+Xfi2GLfxmfM
OIsV/WV8/ulmM82fYKzFhTqjuhRZnVuL+5DYgvdWNoKMs4Z2hxWjeJ6yfBCkaSMczkm7zrCXzpG7
g24OcEDR69yo+YT8kEcdgfi5tKfTM6Wpxj4nPiMI0OIs7/Es5oPUiNEi83sYi2ORmxA/1foaNw+R
FEwiXBEmqBrRjsuzm6+wQxX8KA96UqBkGsQ1ucEZecvGNRaXOtJfTBeHKBx/tZb9T7LC0EhXRLU7
l89Oa/o0RMog44RpFk7+OL96N9gec5arXNdppVSuTIQKOgkb/gcwyooo9PIjuBAJqR0kLDVkh82x
2iks3gZ1XfkHnsh+9B6FHje/T72qjUM8mq0ljUJEIhSZaNmFd6KKCl0FwRvJOeg9AOJvcOoI2HJT
tK+ScDsGZjdPBVm5ybx4sa8HDF+30oW2wVOIAwOql9N+JDpz+2pApjBemsikHLLHjhcm5KFdSeKO
JFma7mHpHrzeGzpTFYHWNzmxKZXE/Gr7JFjcFDjiRPXjIYQVvWhLmHCUP9lLofdwzP6FPnFKVZ8f
0rUthKn9b5uaBhMmyhF2wOfUrSqpCWom++uq4u5jKO3w+tWvJ0pPCJGM9aPY1bKKArppj7oikgn3
myqhtkb19ulFrhCk8cN4Z0Va3wbXdTbwDUEDPN2FZqKAVgeeMK12L2rblGBp8aEeeSvTxwY7wtOK
BPW3jf5lUZDQdB8WX0Qq5VD0W/NeHgVbrwBTjALFSURFaR6esJpMrRVrcG41o7u+c4Tpy68eGmcz
upMWGcdS3tlPug5tfVGr9Glim/f1F2I6pyTjfnth96xUz229RxyDbBJ+JdqSMH4jsfAm6WGGcncN
6A9OLQqpZvV1zX21hFj7BFsEmv8vNrnSOKQuBpknTmHsCgurCqoAdpZmqNJpSj2Z7fHwW/QD0j8g
ZzKg/AUplEXQhGRUwJT1Fhw1YRoNuwE0t5vH2m6MadyatgD3jhATS9DcxnV+2Rks6DlfowfuBBMo
I0heZc68rXeZsfsbgLuzU/YKJBIMIRel5HsRXTpd/KUPvx2edbpHxbrd7YmlV8FFqb1R23b+GNId
J7NF2r0raOORN/EbfVX+oW5oY7F0+02BQochMKlDefua2y2jC8z9EiPyXFcQpnN0SJVxtfi3NLjv
GloG+s9QvpN47+5FDG+OMyL8C0xFTfFWC8oOmCEgAFs7GWme1IQxKkWDkxZAr3bRxUjKHiRK2fkn
wYkke3Jvmh3kaf/8yXRIrpvsz1LIuAC+uID5K8BnvqCmp2zyIAeYrZP+p9lpRlIUN2kk9jBo6N4B
QbRQ3/23ubWvEdHH/6QnZR9pHXX3KjMDnu7cAvbCjexPNfxwFnAgroHc1ru7rFExTBxls6IAcumB
yPS0A6jYDKlhMQE82nS75Bn1nZMplPFJqtaVEm5/HMFm+ZRjOjn9e5uU4zPlIymFepA8SNha1E3D
/+i0y+7B4DskEMusgwKR4wjp1ro6Zir6pul9+o31EbzKB4OLbzyvVnkH9f+ErHCv/Wft0BbU7Xcb
eO3tP8b2N5SzdtZtOLAaLkGw8ZWwgq6RDgnF6vla2oSeGql7o4ufyVXTuFtyLhHw5jX85GN35Q6s
mdOj3jMoDWXAkFM2H2tSVZ1KrpYaB/QqRckz82sqZ6eiirOrYzoyAlmHhUVzdAjIw/87Ya+6Biwj
eNYsrrcchVhHd6fxFVqw3WaYvuS8asDXaDyYJXQpO7NySS1Y9zzxZ4+OgzOcAuXPFVHwJJo83RnJ
gZ4oGMVtVNMqKxchs8GKqkRNfzGMBfDLw8RxQ1TsbzPWQFTHjqrn4TuF8sqldcwmmPcqvDVg0h+T
85xwfeNsfYfOZy1JOcjHjE4d4RuY6TpCbn4jdmiwa+tSJbaFnAX10JhWWk5ATjEBWin0X0SKsh9N
jKxw5S7eHVBMviRvntrUSeqfiq9x3OW281LYA6QAGNew8HQduLtRPqHO+52DYfqCEfWou/EUp+EH
4C6nZC4XNLIqalJ0orUqtve9TsnsQddZnG6Embtan6oYhMr+c2k7omavGTYlToJo+mCymOZLIKEk
oFJriis63zNS/k/nfus1WPL0J12vuaAjZP9f8sEP4hB4vpF6uBC65eeUJMYpTgBjmABH40I+tN2P
uDFv3q1pIvqV1aAll4C+ZQafFsVajLMA2fufApZrFEVvypnoCmQvaZpv+xPGFB7fQzzS4Am41Jds
sjP5WFtz+ei8M7SKQA+nUbR2DojDZw8k5hqeuY6vV0VhxWk1J0oj6ptPYFE9izQFTv64QTxFj9v1
AZdcvAWe8sNSTzLY30BPCJ3tI+DbIzvwEk0xOQVLg0FisGcb59463MZ3A0tm0KBHdaI841REr/h9
BWJ5VlWyH6y3NJrUeKrImvgBDnR42L8Nv52qpM7NL8mYD3QKL/hhEZ/NCOj7SQ5OGxeGu7cSYt9w
JuB4+tbKLvQAwbuA7UJm3FB0rXd+vFnW7AKsU0oplmNJga2BFy0XWjwoS1OVWQ29xi11EksTrugg
5qg3GPMv1oTCOj7kKGNRZQ6w+qdoxrIDG0TugPGfOqUnCveqdHCrR43ZU+9J5oyDuycy6FQYNV37
L7tGpTPnGllBGJ78b8H/LDTI7hhLeZL1yk2w084peubTsE6N/T4LCKw6YK9qOW93Cu9NBpLkei+x
lLELigslbiFfbFt6XbvvOX0V/T1AstaTHFflPLaZe6rvWqwmtR5QvbZAwNI6aSY2Z8DHAnMDj1s/
SWarmYnn1ut3Kxbrc+q6kCWPZ1qR51fkBEv6Ow75eUAIIjP3VeofJ6QfGqO7dJcrXOQG1/X3lJ4J
Pyqn1rpVhC63rK4x4HXjtVZJwOS+QG8vIQMKnMNHUCutdUK8wUXO8E7PxHH8Qn3HZyAenG1wXSaY
75AHvrxjX1Y2CEOKpXXirwDq0INcvSiEDb03WWl68Qm6HNVpNi+HeEHi+tkHSoCq60lgElHM0heE
MWQme9iAANmuohGiiFrHKLVeR1XGCrzO9cqcZl1H4bjbnzLUFhneW32GIZnxM1zskGu4RgI3WlZP
x0OzSz+ZuzGlHkOh7rABpurb3lREos8L5p7UlP0o6lCPYWU0eP12Bvw5Cx4USSYQmKwO98kFknm9
NBWeX3bnL5trRMZL2/+p3gV8X64Zo7DF5TE9IBNHL8U/Zhzj3RoCRmtGtKv2/5iHbD4AB1bjojCk
jsYhvFK5L/TnqAY9pIvnz0v9rZynfMfsPRJIIqEDXpxhXm5SVT8xKLxdwEBZd1Z15z9AvI7edg+O
qRrKC2yHkTyev/nQp/VINCrCKY0wayyHjvHcjPE0Rl08+h5mOzqetMglmLu4FuGRrewx33P/veq0
o8uyGng9dNRTVGlKycAaasZo4r+s/wyHYEms5pvqcs6CKvLpDkVE1IS7zJYNoOsrLYHh12kqChbM
sGDVTYVrRGpb6JUsVzVVTu164bvgbvnbGms0iFVO9jIiup6vjFx5s48OzZanzcaByWU1Imhjul6F
4IevybgFz0S8Cf6iC3e1BWNoIG4dAfzC/uCae5PL+f1i0jqhvoOW51Sgcx0jdd4Sunb/epFV7a3g
4AJgirc6xz4yTHi+wdSsY4/Ups5sT8FV6kHuhRVrHAMnqL9fLmpV4yt9bvOOCNg8ItF1QKl0bpJZ
Yk2nczfb7LDWImNegShu7sdeZqdiyz7etS+28YS3+FVle17WSYc7XZLatgEsyGdALoby6TVRso9E
K7OSyw5MPfyjpY2DLINs59C1Dm6gDlaipKLevXxMkNTsQdMGngvOXHDHBoc5FCDIft1hdMr1ji3S
qoO5kyQPvfYB9cbYkGPXLHMG6cMXwOd4gq5/C5xZ1qT1Wkq1RYBYeIVAhn6wb1bl746XCEpe4gBS
JLD8aMChfiFBDYo6M6MUs9bkiyXlQGyHaZcbUisuNBG0JE6EvgTWjIDPMaPf0LBL0SXNuHKBbV/1
lTiHVrPZBn9AqIdwlJCEvGtnQtQ31OrGnK/HmjBAR+Jc9gCL4zuX094PWAMqz5692ACmF5G6qTag
7mTJmUtR8T99rFQGDG9d7OLo1SgpymfYzlH/RKHGsk1ZgW9hTumnmooE6gS+FLOoUREo9slVXpfx
baqv7lnTkWF2sLscFl1yjo+uzUf3f1bGZMTqVL+iTn5JlPgWtuw2m/llO5qjFAkti62xWzPwqZxM
d4LZ/N0nws1uK9cYrpBneIL06tItzLLbimt+miozfrRj4Aj8JFNt4h7HIzLf1HyUPIGLwJ2aM9LW
Nxk/0NhsuMWqg0QWpMmLuWvI6qOyQudbKKUJroLt6mNit/nAPUfE/2DyOVkB7Y9rlJtbs0i6aiQi
65ZbiO9LbOTmFueSq+qFDhiG/ioaPimhrSq5q+20+xEOwoR1fsElGjTqUCudCU/1gUuhs4fHFUI7
h7cPwXzvQoFoyzV4+5/iuLD3Nv+8SDhTgIDQ3hmgf+fXAiYDW6K4Bk7Ly9GgP589dVIoKbnOJY2z
o0Zxh4Ch+1GKAsyHyEDXIhhnedhrD2RARKQgM0Amxx5Lyf2SwV5ELwKh5OKWuhk08wwDYfETBE+G
KaO1KGaMP14BA2OcWYTAHdwJKVyVZAkQRmM2SlWnWIohug5IAul6v8LU3YqLK5QBIk9YYdyqa5kr
fbm4stbMpVUBTxWEf6r2rjWQP0s1jTF8sdMj60Ztx4AyMCU0RIaTdILF+PPzSctvCPAHsCxHnqrs
GgmG9MzpxWTZIoyzVtYpVVJKtjpCRLn4ZS2x4Nty2XrKLS3PgsyTKBokKpaSy3lw1I1vL9SUIb7a
NBscotPz4Pp/popcScBH90TgjTG9rL6WqApntKrN9O8hQKqC8hbfi3bspRLSgF3biG2rE1iwgZoV
ZopuXIbNfv84I0ot+yZOsjBjAEH9hiunV2h6ox8ZFrNma8S9n4HDFJh292mXmnd+9R4vFxaTOIq5
BYrYUGhPVR+XkySuJWL9+DgG455DYki2tQcEs81sDRDr1sSQyRSkHWbXJA1/vluSjkeGsIyGV4RO
FfyTlyIGytubcU0QTA6tQWDkLce3BC/gd0Kaiezl+Bs0OzlNpKjks2zwMw1OXKBK7oPguaszaBHc
1iVLciElElTVUvpuzxejrNV6MgptArE6WT8l83ny9Ogq+zpc5w9e08JTfD5ZQKpdpLCEKKz0bxoq
KOTQv2dmFo4q9p8npvh9MO5CDR64M3MSzQzmsLUG2wh0OG8P6GrbBi/wbk05N5s5A1kxDIGzxE4j
VyyGYv7bhMltCrezAFudzKcZr7an8G/foPP0/roMupv8hjnFB42q6yC7deABW64QmxZYTzWs3m5H
MS4OUmD04TXGHPn5s+6DnmKtddjVHYBhqA09lYeioAdIwl1+56rhkSf6km2WzSvFoN3lZKORpuVg
g8L4aYd4s3BE6HZTJ2Wi6sR9tmbM8XgL/qd4id7gWW3VvhOYYMZCVd9qmBGDk2H6Qr3az52hLxJm
v32kXJnlNAjEvz8C/SgidUMsUvzDgdUn9rOoQ6jVUCFJX00yIBbE+as33wiss1Q5fD6FJw64d58Y
bYk16lm0KMnWVBIGWkwj8UkTjt/2MUvl+rzYIsw+9PBX3jVQlLhd8FMBZfuyj9N7HJvXotC6sEkx
SrPfjYOlmWpxf+qpjT8F3rcaWFyMT/4xUG5TnkE6xG0U6tdtHEHgzEqykWZCmvHmiYe57Ehrr0Zz
ySbwIrqjbtcFJyI01eksNi2Px2OgJcORwVLmlgsvAxYmgag0n0nJGELQposzGb4ol+8s2vhJhedx
5E3HccmVXAsV9DEI+qLm/+OH5HG7/265NBhhmx8cfP3Oo7cvJ01D9Tx+vGQnUesvmi90Gxihfkn5
hKvTeDAOwxiOjVUBkDIEuZz6L8C/9mKYjIbnPTaRdk3Vb73BHp4cSn1tg8TdfbHnSggDK2wCtre7
axJ3n2uzphjexjahRQiRdeiAskCsmPDoO5LHY9SH6FgcttW8fyhLtOXIPL1dPwtILmAYR3lMVYPG
thqvf2PjbugyEdTMCoJ4Tkq4VdoBMnPB02B4xVrEIhW7MMqQTwUAdf0fH6LxJdCEx59hhYQjeXlT
mk5PYTL/16oRiHmYMjGomIMgAWZuVaEv7xk/CpbWnPbGh1SMFefSCVnjtVVjNulm7jP67RbczXRX
tUtkMZaUU3Pt6ErMqcgTdPfZoEFzbVLm7XMlWifELBfIxliAnqzZPZ3RVw+wViDZvWDjIC/+PVdD
OYGHoEnc/X7XPSnnOVQUpWy4cPve77p/xTy35ct6ANhMMQ4UTL8C6kIdhGjBB+IRi9UV618h5z4L
X3Oy2lbFpkw24Y/IMKqGciDIE+xMkVO15NqcGiOBx1IIF3ldQBpzzCLYcwcLXYSvagVM6mSktOvu
E9J0ohY5y5cRW2d5u3mnHGixRJvY4A4n44lST7KZjt3KuXFbMI2dRy8uUDXwWT1Q/8shJh48liG9
OW2AfMH0eTDVXYHbrDLbXJkHKn8wyBsbcPUzb40hvGV+CroTrUwtmSZVE1DQFH+s0gWqAELhzwK7
OHAHz0Gy25hl1gfnVNGy97dQo9bA88p7Lq2vYyOE5uuuptsi0ALx+7zfcmYIbzjd9RcIzgHFILQF
1MzIbf7Z20WA6Vv8O7o6cMqS/pXwowXbYRsJQSOt4f8PJVC82JtaOYE04PGNPbfsklz6bHKkCNa4
7keuFDM5hl9dMQQc6+gwGXxPznT+IMPF9KTd76txwq6l6lwLrsW2kP+3z3ibrvso8PF7bnT69oQF
JzpoJPpnXJMkR4HCDn23beCbdTCph5549KI/XRzzreC4OmGXxZcJcbKiqbyexqdH+XrEYC3FQ0jN
WNRbEuzU4x662C3EexJfZzHIbmhHhDiXikuy2XTYfyB6/6qvQwpPNUPuFW3KiX97Q4sd7YtOTNGk
g2QkdGMLfTeiFuwvudPiNvabowIExL9GL/ZvuLwhceEdtF14QsCVUm2Xin3jDjVD+b05Mf2JK8BI
XyFt4wMoxMhVNPy4D4LhYMY3hezdG042juYIOpCxdsVhyMFGfP5Ai42NX4y/ZoCogkktxElt107d
QAtiTmZIyr35J6Cw4DEghA7sKpdYjveUaLm2TZWPngYtArjIQ+Z/DTibNHHLtbRLL0l7P3+DSzv4
Ba79MhMLFanpfcHS27nLkXulLrDXSr5Ut6LAfB+1YPwu4oTog20VwRBFIZFFobQziuF2mjc+mGOK
BuHsms1kwcfdlsxg69kQjwLhMCRHe7Dk00eCI7rP4SQVLVRfGm/AvpTAcLDSHSeJsaAM81RNER2t
8VSy6atAkkKYxD3LjRR5rI/QXwzravFSHiKOkV3r7ACLl6/4utUYf5LCzT3bvr2qj1utoMqt33Wx
0caMJUHmzPUN3+odKe0O3dEWPS+Vr5uQ/3bXzpSXjCzz/CEqRWXQhIkeqcZwrDTk/3pcrbzuOizl
Itdj+ALr+N6J/WeseOKbsNotvQv9YNncwRJ3inJXX8RSWbSAbzTLnjYhz53AojKuowhgaRf9f4Uv
tdQImgbdg4BAtTlyWy5KwyjR90SbKHx1c1ESEfBwAbMMcjM1nKW5ILeHR+65icyFZWiY8C43SOis
QofUxKOUS2kZTaBxNgqw9yCZ521DSDNPgcsXp/lKqO7Jtiko6IpqzawuvhkV4WQ63kcz1makHK0N
sj7IDo1nVt7iHz6rfrbStzVwYDuS3P1A2hbSqrnNmPXzZaKabtw2ZCS+vnzCPP91RABahhIgeHao
zs2NPM9Krq9kvRM0jjHtJizkQ52bj/4WJoX91o3z80dysJLYoGKApEslowtsEBViiKIpGQC1QjWJ
cWWW3XQzLzLd8U5tt7vRGt+oBzdqcghgY5vLYeq3Mltuf6MudSKFzV6YmOv0OGFaxl/8Mb+FAhkH
Y6SOdwaklhb5Tg1/aVjepOyqK/ZjIIT1bqCRgYB/FUoZcVK2NlXkljP0Ge2MbIzU20SHer1LHhkV
y1pciyh0b7JyH+nwPbMq2bXS2b639yLz5eD1fd/zT7qT4msVE7Y4ZlHe+Hy68NXTlP1e9NvyBHAr
VEoymw5s6SNmfvYdPCwRgOCBpMu8fttP0Lmu1zmdBTADqFf8YvD94kEhslCIZhBNhTodFFuZ8316
x7agkbLGnJkAin1gPG8mIxnEbUm5yp4k2OWylPNiHn722yCcxy4HDZQqQPu+2VDRK2LkPsw/U5CD
GPP8ZJl5ulRxE77a5YXNFfwGt7TEmiKgRJC9ZqdbkyGlFzhD+3PQbLgYtYBLbvnIKT6KrYl1naRO
BTTNV14usR0COm+xRDrFsBRQkifn0Qci73/4XpWiNl0nJp1cX0et0iFjwRqoZ/xwzRhlfQXD2YRk
cpkrCk1PP6gGfCbkT7DfoZrpCuhtI0lClAPFAAZMd9OwhU6qTLKJR3nB/ggQN5sk2XhxzyPkMPxG
T+IbXfcx5uoBGErk9NzlnnhG7NuYToazPODiWqbjf8WmM5p7pCKWzCncFHqOW2cFMLiT9bSePPea
HOVJRmdyVfpls7sK6uTAbaFfdARax8bWEI6OHOYbcUOkQsK5AqCqdCOyOjiIIWNRwEK47Fiof7P/
CVm3rT1Qynz4OTdxV8aWPbkHpf5b2xGYaoVwZIdKAFHnFcZ5aSEmNua7eAoJw17Th4spUG7cTdPU
/i3kTmFzniVjKbxxYRhIN+iBQ8pzGJnwypheeqyFRkbc7gdiGFTt9YsDYY+RDum8zrIVH+pKdujm
1t0QDCB56faXHnbB/gS3SEF+8a1mb7eT5pXuCBeoZV/mSuPmbaEgkyGMu6FZMpCLcsZsxjkOv7C+
egSvE0iNQqpXlYsScVTZl1JnfNVjPflndNPxvfAI9dr4ifmXfMn5UOpa9kn+9Ln5BcytnNlBg8dQ
pyyu4IaF4W9+ewQz36LdQPPfU1seReFXOy/D9WEzYha5EWUHUCajHZB75r7W65Xc7tSX0O50+dRY
TOZQQiWcW/JYZIwqCpZfa9mR48o6l4GwYJ+oKIRfkTG/sMyZGZP2RYVpHUW7O5BKK3oulB4TEQNl
ppkYr5AbfrZ5qTAXDUSEOA9EV67XzU3OpBeUBynBuYTg4C6015BbOM3VgEz3HB8GCAbVZvt7xRR+
QHJ5EKHXa0ZMlxVd8I+uKKWr1vIsuiDGhwz+HMOw+n7f07uHDXvqY3fIB9keqeRdgIpvnk1VqXHT
VLeWY4kDGp7mkXNVUIPRX8/nXTZv68XwX9gzFskIGsrBjD9pSRT682HXVZMlomZ9ZdBeZtpvCxHn
l299bONL0i/+9bRYW3GMdlrz+sHl/q2Y4bfZEanIxnzfH3a0vG0SVejw15ayBPNpVzChpqWGrFBl
FSVFYs4hnfsdlOastP2njt6QWJjnAG4ygbndw6OGI+xX5yFNugxJMacnUtlYAXxBCJwHKPZEv5Xp
iZYejznlA0zem0oZASTTohOrL0c2TsCRK31VI1h+ilqPwFY16RfoF8mFqnG9mLUrNO6zRnYlHbu5
FPk77KkttlCu8fEHVeJrnUrCsBEWXRaS/+7K/tgYvJOXKfy1NN4e6AZ9HUV+R0GVmCk49/RGGERc
y+ukoegm1HEvAToujcW59ePr+tiOCd/tbCYiGoH4jt8cmMN6VzSQfjiukxQ1ZAyCql1Vt0UiDn7n
5tC+G0gOwNpXjliA2wXUMh3jmzFJgH1VEWXn+ybiVfyHg8uHZTULc1M9K4uQuZQlwh+uBROk0BFU
Mwguew2YvShojjB3KgRpFNfBinO54Jvh5yEHl/v1u9vTJJmSEkKNPKQFLUijOjPOc3B+48em17TJ
y611nN0hrmMmuy1UsHI0yetWPSrqZHQYK5EjXPPWCzVAPFT7VcalXuovC+4A0ZQSVXgdIgVzN9qR
YFkxvL0V3mpEPtylGyNEZhcJXYrdGf6MKvCwHTI++3gnApHVYHAJQklQiIx6uxh09DA841juVQnV
jGFCIT56XxkyCpT/2a5mH16QuJhMXdVUXN+JQAC6Xq4Pa8lCw2VnvurpZ8+Y0HQhZQ7ZL2XBEO3H
hauleXUrXx8R0mc3RNDdlWKuniu35o4cYKZq90h4QGeLGu88kdorc1C9tnwpTSdWspa3m2BZH88W
4b01NgTctUzbt0sRdEGDTuZf/xpAVwwqD8YKnXhTyW20nv2gM1kBwv4ldZEe4hmKxtS0lWTxXQ5V
TBUbgVA1ABP2IbqCZsQOYe4War7P6HPXsYEhwRZWm9Vrv2QfY9ykaakBlFTEISK8k0i3TbcPg/Rj
UWD1KkY/gtgIYWdLPFB3TiiVCVbWRaDFpzh/kqoTDq8ck885j56gWlfozM6dYkntFSvrpN0/AcEf
JAG8dcnUKYM8TlUzMtTnOAmTMVklAyunnhbT4Y8Qnsa0hYQ3zHdqJSgBN1LXWhjrfwgm5zE5vonM
DfStw4wfzP47SUIiDsyNf3apx1iP5OcDOpGHiYRBE0K07HtHf5EfkQ2S+2bxg2+fcES9yOj2URmX
o0YONFnINxraL8rrm77gJplO/sdFjSWzqJPngt3Dx8fejf6zLtMy9KJ3O5RbmIGXZJ5gGuZW/qyi
NrpMop45/e9IQPPcSsw5Ng9xFn+kNhRUNBpM0MTjS7XexFH8WyHZ7YlcI3Wyj58Wwk1fL4FaXMD/
t9v8Uq3/09xzkRQGkQwpWVD0hZsN5osPpOQ3S110fDxKg00VW9CGWxtJYJGTb8WPy9uQbdcKaCwx
yFOFu3FtcOMLmvAhO7aLtoQwaYNmgMYkadgEbWVh1kJKvzfUsFd22Em/zWTLtMamr8WdZ4J2AABH
0c5425iPDbZMqDtluhz5DAwwPojQMOYE0cWASKuzzLZxtydsfmyiCPybRMF2GFAUTvTMbLDJ0m/7
5s/lJAoBZQf6K+BTEuZPGsXObXYbtRU5HkKLBVBXAr5WCQ1MZphQx4dtFb2+zoHuZ68N8wxtHtwm
lBR/h4zJevQLDpa2wOuX2Sq9WN8QdU3XApZQz7qvmKcZyXRVly/D7/Px4NsrxhgOssPalB657UxY
nwf3CYSuEgEtm+34MMN3bct6DwFdvsiY83R6tBaHL+dpUzgjcZhZBzNpe+yZMdHcyIUWhsBx2TJn
1Vo6uVUCINi4vUQG0I61LFLp9LNpi2ELfm3stB7Iez6o13GdKrrfgyvYbe40iGZouY1KwM/6WcbL
BIZ6iPruTvi/3xdcBl1VZyxuPPc0mo1faYd7tBcoPq1o6RSvjtVM1lX8D2gcxn4JTZ7pGE13xtVV
Zus553FOtxPZHMvLZxAj+gLH6scHfh5m98zX4RXpj29xbH8FDpif3mNdypO3SXWhOROnlzetGdGe
2ub1jUSrQmN8uwO5r3M2br4mB5UKZhCygB33mq4VzukZT3I0r3S7CMd1gUiMGivo4Pya1SHEqNnf
NHV6G2N9xUOBapI+1wqIYM+ok3xbRNKeB2wbPaQdWLVlfdzPWjLBP+R581pT5XUsIxcTiOY4Xn34
SV8IkYNTY45WUUqYges2UIXwAgVdMNKx9nPfstVlDFL5lEmciO67h6C4LAtsk2Whns6MaWd9N0zf
yKzCM+adqfjoAEoIa/5woABx5Lsn74N7kfR58dNUsJXsSnqifaiXKzA+LC6gE44qjmXs6qitqlRH
uQpJe3v5MXpH2A4WxUMlqTQl0U9AKmIL5vgly0iqa4cAu9gYq1P8LYptyAMr/EqL6O5VwjnEVDHY
FZXO/IKyNASk0LfE5Zdjr/LussLpr8vOt5z0YQREbRAWaW53qWg/G1mhRtVGcX3Ye9Dz60zZmVSJ
cmfXasg+w7NxokFaCMq9sUUm7BmorKF06ELsnNOU0WScck/706WVKov1PZlWPyL2YZsnsGrV5m0O
XTMCYypccAIPgDejcwOPJraXSQjT9ptUCesOY1hewaxfS/5D3p0yGZRluCGmJfSzqxN0BfjmxGZl
50mRta5/U2M0QSHPjaRtofBJpWUHrSmu8oXXIz4Fo9a4lYtho4hLDYSbWuehF5wOaJm7R8zWIJys
TxkTXtxRew+iLNUasQcC6EsRGYnM7DeBiqbeERuos/S1AVKK3CtSV23URIpZH60JZJ85H5xQYCRt
v4LXo9SecaQ47qzstViosh0wA442kS4XgR8U3MCPjsUynZoNjGyAFmsAiftwXLmJkk3urQvXv9V5
QiOpvePjhaefkD10l2UVxPlyNdlvjuwr502jlTtPZIp5Jluez6Wzgf+l1KUgNflUxUrg4T98XsTz
tnJNm6RMDXSRWFRCGebXWbF/k1V8nRu1sPqRGAWTL6i/1kBMQwH4qnfZHMrdPT3oPXR4+01Khq0J
HkOxPXkMnqHuIeE9IlSpPZYZ8Ac9dsf4y0+002u6poEPeD1Vyd+EXllafqyQd+FX6pQ3Ca3VnIUJ
+898lIFlfRDd77kUyd67PMyC093vujjpRwl8hPcpDgPjL4riq0Yhnh7QI5xNP6E97CfLokfyj5IW
WqnyUwdbjeEIALfLnpUiAuiHoa/vbUT6iWoOu3ysX1lTiN3FDBkVQWjmLL6F68Yp3bFjM4jIUPzU
O63vqI+snO4KOfVV4g4xYSr9rKtVEhlm4yZvtq3d9/rD86KHghwf2gV6A2q8QAnNztLTluYheitP
vwzQw7AYXlrNW/JUxTPC/wqY773ba5TYo6cJRAp2CXB5CSzk6L/YThBGeQ9T50oBJwL0B9mWicrj
mq6CLp3SrR0xlD8iYTDsGD6vrgkW+eeP88OE0rxAe3pjDc6hg2VhlZCFzNDVAzjFca2AvE0xTKKM
aj3RyzLB/o0yRz/OUqpem6RzTWsp1leqKgAwqK9ktWpdb54bzFy7w9VML6SPnFeuW9g12n3vbnJp
vXYmzsaj9xBnz3v1T6nL8l+svJtQpJpHO2heaj71H46rYj67avrx/d2gAO+SqSFEdnFzbHX/gcsH
l8JVr4dwxjJHo2eRMbXsQmHxg8hkn38iZt4rabOCLEKG9I7FDW9OCByw4zzIEJsnte9LKtc7D1hF
WkRMfFZGz0mqWix1Dr8kULI0Fs+lOQtTutl8Hw2K+Y3nAbTtjnLO6ARp8nGbLk4ksDyUhtopliam
/M+i6l1RyK+hHPILxN3jnptk0Hw+U4ZCQeMbAFYgPzotHvqvIkr+cpXxKvg0mfunfiPpewqP/lEb
o5RTQV7Fkgqj/UyJ9JY8C/9f+fABLKvcgqhIzT3xn/mA6fVze66P/AG4dODaopVLAHFwQw/dSaLt
7Cm9n1DQk8QRiOHgOlVGywW+d/1c/K/74+ph4yHUdVMSuEXFXRSdcgLXXluoQxNgNmNFQXrs3ozJ
MlFU08lOioU2NOg7Z72gNftQ+APOfmDwMhd0frJR/Zrf0fSwhPwF19wrzNg7xvNBWO5u4vjCapWH
O27Hhju7XBY290bOkq4DI+4ZyV0MPi2kOeaXwmta9QeD7F5GJ3rX+N2LoRK+6g9pP8pPmO11YhD4
8tJHKLsDrEAftbzpshfgsNRNJG3Zo6Y7itTA8Oav3nJgcnTkf8EE/JyBkGRw2vi8zSqjA59FgQgJ
s9crHq5x+ZwmINNGBIdDqpFab5Y5uirSBn4UIt8MBNi0sxnyAPv0fdxddkQ9bqYp0EzQt3XbvL9R
SgKGOpAfkuTngE3Moj7LOUUuCw6uWy26BvNqpsDvrS/36hrywWceSXrQ0gZKR7VzaIsJmbNgje/n
BGqeQ5HwsIewZ8UgFPZBI1SAIEdnA4MrXSJfMWb1/ds2hKfbPNK7jzjIWkjZfpV/wWNYYARvFZy4
9+WJbQyFYVNhoUTuu/anO14VqzXdElMADppuugiV7N4sG0Kt1AWWjHfCJJEF5iulezELIpILyn/O
2G4DPN8ZwwHDyg+lSI12IdnXRSIXwiCmBKK7zXf6/nE6vPzF7Lqws8tWHG7WSxfgtzOZ+ZshNLBC
QdBACbOgas+QREcfyu1tLydEeHBkdCtXPA66KJtWpUJZRt9AJfF++jBSDFcAQMP6Zcd/SKpEUVtS
uXam+gGPU3HIeCmuOKWsHy9bd9gpIp4fTDTwMGufSab+ISdNfWEWiB5vu/6Tf+hzp2tan2an1h03
sZZmFle+nSR4G/V43ZEEMs/543NSSiHwhcZephkd9CrZOp7UgUCEUEqH4PxFjdT4U3etmEV3h8pr
WbAt4EgRhd/mUhxtUjARbmWYOMIplcVA/lJINCwxmyW4Dg6lG0n9ObVjA05CwU7h40qbCkk6L7hp
lNf3jQoxGQIml9a9xctcuJ5HxVjT0pIqQbF2/QvYQ80E/VN3qhyfOOq3VRT9khXyyjtZ5EvZzIRn
XS4Z63yzKBsWW0kq/dcaKDFn67yFB7QvGD24mHVTKoVFkvRuEDxdCKPBPDUtjhWSJDgeH3GbyrZo
SQ5ehALwzGhkd+tYOacyJ1r3o///MKc5BER3fQEFMypfg1fGIbtkhzLA3Vg4jeL8/Qi/nf15Zm1f
BiG+V5FcQ7irBULvzdxk84GyKgaYlNhHph2DlD19nklJmO77FqtZKUT8QxFgF2kW6mOUFh4PTB/K
nR2KEjJFq+3sNx+S2mw9MQGsDM/RADS4lsewAONxA+jzz76p18QWbnlKMM13EGcLp5+Sngwfjr2V
zgPTq/D/NKvG2zVTK8pTY9xMeMBk//S1UH+RMMnW/YnmjiOT1lTp0n7bK7ko8NML56264QBXFlyN
pVCh8I2ncvkznnDr+nSgMSGr80I1uZ6JVecXVrFMt2W+ruDStNbFsvpvbOIyOcCo9OwwAG8Ok42n
zZWvCHN/vyIsTMo7qvEDPXeSnYvYAyEUiCHWEe0ZVhNg/oUliYrcjEDRjVqvMqNIohje/7y1d6mH
0gm4qY8mV2w7UJ/RyFZ0Z1rysfMZXwmB8mE/YYAI5SDb39h2xJ/IZxNcOOMpD5iB50VfQyripknT
iMYAzp4GEJuiLReUMPNQLKp3LlOLMrntLRoj1wWht0lHx4l2Tm4a2u9o84RgKfv7sIh/4EzRxF3p
fV3S3Q4wAG3h+ZBY1pgCY7aefF9OPnMyB0YvLvOL8FwDXOZaWHIwScqmQY/TwB0yvntlZ1RPuv8L
SWSQJ6s9wWOfqh9CHTvWU1my+YHQ3id5ETSKQdyfL2/2QEwnxHZo4mXnF9f3Fp6Ikf8ZWBysuwaS
MH9drrv2q2R1ytcIV/WNxUfLkQEkfe/xj2fVNymcmyyIbb/C08YaApu0Rh0nortwT4HJz5sIryuw
4ZEVaBN/i+DZMtRnGFHlYIpoyivWD03oc2reIi9qLGuQy4i9iKkcwNspfiFkrhPkXvj+TDakJnTs
J+LlScOBwwIqaOFgHRbDwQmRWJo/F5EI60ehz3RqvzCprwh/fHgaeDT+P8RBZQG9vgaGqMK+QH0t
6PsXCqyDP8VSYEQ5xNhg33tUfcMbmdeXUolX4IMX3FFsdwE2zltwV9QqNQXZ8GvyhvtYb/vhiS/Q
3RL4RJacymiBcYRL2q08BewEm6H7qu3Rdf1At0VhkRSCqvr/hwvwAtXELfKLBhlq/0aqktd+lvyz
k54BzO8c57zFSvWE7wGjZcGZ9IfkHDwI2rkZi2xvgLIn+PmQjVX6ZKREKVPJmBdpKvP2/hIjouI0
M+UsBfeLMSq9Q7sccHyzYss4PsQP3rOVDYafLTVtGubSN4WGBV+yXeKGIUUUzONknUb+ot2MoCl9
bqK4S99NSw9j/oiX3oIq86rLTgKnYesutGEMZgc5pcVFSyEE8TmOPYY9L++8t8dTscL5MtHldSsz
yd8yxLH2agmBAjJ1pCfEuyH2DTU4ReVp8CkA0OZOhkMe1uz+q7GV+ZcTFqeaDvGyAxlLEo06bxRq
5eJn8bw9caQnV8cx9ibFPiV8AEK3vSwtd9+uVAsAGNo46Sy5GOBLW/s4PbhLa5zCI54pq078g3rF
rGPz70Te9692tfMnhU+NHt0jYUbZop+D8f4e8wG45fZtMmODb3wTLdEgT2yWOXLqdVU8XQn+ygEy
b3j2wusGmECE0kMzDZzKiYL/MiPV6+Bc/DQgFWl7IASrXHqipsyqXNJa3ujqaOQAIeN9nczKB/2l
+NJUDwtG7Xa+BRW6L3Ntsw2Ss6TT+xLZGlSGYH26dbaT88+wqpZbh+IFgu45VEf/eyoa12FwBIhb
tDNd9MT9SHY0G5w8MRn3Ib0/C0HCb+1NitKZ4GFjmuFzr231AMCyPZF5ngU1fGqjRa+vtMcnNlBi
RN3dZjN4YaKkOrclT4RTThaG7NXfYALTgyeVqp1EbrNCMDoSA1wxPVQFQ4p0v41OIkqJnUYCDlcB
PACpuQKgJlqo87qe0ygUx2GPD7efHo8F2xQzjbDteakwrvuGW0IizD2WN7Ta+22ACB+Sgv9Cb2cN
8CGU4rGxQaIfxeIUfMrM82704co8VvVhC623Xqr7+FrRn61doziFvPF92uF7iOX2cQCAJlS+3xw5
S8/BAuVGT6a1SQLMxSGKWSmF2KJm+1SwrtbSpIE/DBXI4+oiTImMy/nzbYOwoM8kjFsbBYmN9bD8
KEdOjRCGXVv9M1e2CnjXOPcB9wemWLKpCHAP4YqaG2w79kJpSrDkpxvnV/xSaAT9PBY+FO/cJDrp
Pz352RJzxrpT7dQIOGTqk016btCpBx7T4TF4paeLzbfxjaSLiFz3eMcesQ2FiOgrgE8us44Jens/
ZeYPQSM5P43bmyRQX7prfe+Rk2++IMTKrzje7ObgNSCqeYNCzeuZ484Fk0RqBuHWwvD5vIpaUA8O
fEXAFPjFo7k6ojoTTu2gG94eSZ/T6TMMTqm1iUudmhs9QcitzG3l5kYHi+Xfh38ij2jDecIboOWH
nMdKsWFMVOMFqf3539noj5GQ2Cz3fWwRHKrSFuD1tzLP5pHcztR7BLnDSSfDJKF7sFxahAfxh0tX
XUCuBYlUIcpaf7PyeHKdmNcv4nECSJ1NNHj+aI2xossFVV0iOuvMdj7YeZlPpAFcNgwBvHvtisR3
RnXmqtc01+lF6Poo0CftW4IYywcNy4bxbWQHGcJ/coeM+nua5vOoz7eFSRkp+SDy8SdZEFI1Cb3G
F9ZHbuzrhpgKof2YKVIcFTz/ea9vRh/FfDUEC4c0nHBkpYi6jhgUsYBEAA+Oo5cuJhbKZnii1MR3
elyz/qdXGhyzOD6CTQo+UfaDaBfr0rIsvKFaMBu/f6ft2e6GsPFEkIjqbUOqmqQnHuh6ojgRXxDc
SG4dFo1pj5wRO9FcsXmh42guvWNacHs5caZ6lSR0R4ql/oQ0PLuhSUzSPypOFu0+ZEswOCGpfgJm
W6j4VqTejqtZEOaqPnFoNsXsoAYj+hAEuiKk4wCa+c8vTGctJ0f4V0bpOfL5bTi8LmF1uyrw+2ku
1WkSo0mqqdhQxYehMHYrj31B8VWrT3qy9L0JMMF58ODFLKyTnrGd5yq+rflRuuv3fXFhLTMXOipn
wvN2HwG8YmuikVoxjc2NYL9neBujL1LjBqboh9ZBcxqHAHaxobaSwFRXHieVBgD65yWEiWSTGXXV
LZx6p1ah7Sipt/jGNH/8i5q8pTCVDDiXyS7fgHg70z56fqTykZ5Jvc2RcrJ0fsPxhtxsePTZ7k2P
HINiJikw0aKnr5x0g3b7qaa8SPaA4Tk+EEonREKf0iCUvc7iSCM+C18U+VplgLosJHHdwWbvNDTk
LL6ZbEHWMAdAVLpfHpRhhH8NquIN6od7J4XrIu0WAZ0Sb3dCJm8LwVX5yeJcEvGDA6VAz6L+k6IA
LWxRklNBxd9ML6iHGt2KbA9T6MsWP4c48BkY1yMi+9SgftPA1s3PnC6od5cxsDyPWSAyiNrYzjuj
ynR3OUi11cFiYP/Ix2U50qRQPcgKQipG0uMQTc/Bk1xrwNQj1uHmZa5js41p7UYem/zyozhx9QYx
6waYupoIeAwzQhP9iXKG3k2e9c5E0r1ao8NHdYmyb5mC9JvYFh6rhktXVLdoRx5F5KT7p4J6fRAc
7RUwnZzeEBitlqhgNe4Q7T0TB84T3JRignTwrvb+LXLezA2zZBUR6RabmRy0k34g0HgXGg1GueeP
Jic7r7ghUlR74CLhNPI3nLMBc02j6IKcoaS88+WzrxLY8ibtD1+HQYGDSch797CDBuo9QDiHQqzP
cETiPb8XN1ei/5NJQuqFKAQ11B93k8FiysOtC2q2EPTCDSKVdddRCtn8bzKU0phUPU+KShE9DJpr
8KFgneRgnuJKsBPXhIy+a7UKQTDqqIPMfbrQXRC3cGUWdJaJ4C5vkryRRsuXo75NZG5Phvel3BZH
wTF1aUdJI/CWl78kc6OluuhD0r8UG3ZXQ8MtnakoTJurOc7stxHrVaq7mfoVBx8A5x9OflTBV+Ko
lEKf0FeuiB4XDcx8eWiSZqifdUO1+K0Gd9Bdv09PLDSwETez5Vzf25QhJhPnjr0wFXtqNgMp8IVf
2Vb3VnbclkynHvEhSJsKjPNeIKt58avf41umMiVLYNg5LXtbEVbiVr0w7Y+2zfV5w4q0gXwJUfXd
cJ9nx/HylzgBcg+8hHnbybHjYZrjPqCd8I6z+QtmsQT1HPL+0n2OiDsNVXe9LtXc0vwWLdhB3PyA
uYF0HmDMU/975whsKkS4K978eK/V+kmxbALkoRsw0MaIRnsBzmXHUJNqlOmhlk/vV/a2a1oS/Uqi
S7E/bAqmA14/mLRCSrd11MPqbBOS/XWmwn67Cd6v4UlskbRZNu9DaEzFXs/da/FI4Uz4cwOaSHyH
3sxi2rihYvpKlhUUrY3IJT8pYzHhVPBCHY3NECVAh9E5rVDcGVhnhXs8lAOvkRZIBTWOZSPykkju
KTaSyAdROxqdNzwilD51fvBIbJnherL/BAaAbgjj4nQE9BVeTy2ehjzjT8lIyLZx+2Ammu8DHrna
HUIekt2De6OCjQd5CN/ii50jrXa3oV4QxiPBDTTjGb8pNa4Dnb7yvvIB3b2rImS6H4TDvge8JIJd
s2q/mvUMO8QetAVq9njEog16y6Gk3p8R+MP8dFnTW/n4wPLSlNJ4A1J9C/6GCWjd77BNe+AFJFRH
X3KAKf0tcCw8+N7UuhucQPSkRynJS0AtV2Zt50yDVytjlD12ujv5GxQMRU6ATIhu2AHC75p4DhQk
N16xjgH1N5Vozl9cEUNbSGt+TNTSq90Q0GE+JFuCfTZWVFsUiGHYkOno/CCfgIAxJlk+C/epb762
6nCEkFko+iL2v9Ncnv4McgBe+ZmX3ypiIkeYR18urInzn5sA7+1Jnf5ju5vLqNsb2uMEOq4+QZnn
VZ+7MWR1Jrpp7FckR76RjDmGz5FKwtoCO7rAHkYZW2OLC3+Mz7FmtEKk+juFombMNK8kkXsnqoEl
rEwVmfr4j1NW5k8D6oJ6A+rZazb0wJ6n1KWAx1JdIGIPGzITrBGJAqwAP1ivzfsiLFdoF20fM0RV
qb1slYym/cSnZh63mouhomUYQLLK+GAmskHyAIfflt199vFIUO5nnkC3GooTPMuFHKMMnoK+c9jG
/Av9+wut6/hYnd1unLN+ucDB8yI86ilKcXArxGo0pjzFo5splMWmVsQ8eT/KJPRupQUPDvqx837K
JulXz/J1fCLWvqu4nM9TcSiFkwdUpNLIkdIMAgh+DmEND/znVNXDPHifJkUARs6Ywy8wO1Zd+h5A
saGQA3e2fMnaW0WN4uMo81MkREjGI05RzUQxYN+G9YEFjlri/xJT78e4sZBRxiRa41aUyWt8oePO
7sJ1+NHOlFRYlR+5lutSRfkBduiqYxvZkQhN3ZGFe3bU8tKH2XVNgQME3NPMa+XZDnq0Ydbutes5
G8dguC4Mzlx3qRy5FIcPyzH25Kv35xkIVD6TxRD+JL1FXZsDDZ/bM6QI/+tduBfnEw9u4333YfMW
Weo38hc9oMyB3EqGik0pwNsorcHvLFyZoL2fK0xs2tnSKzSBIQ5jDbaAvtMiNiBQ5K4eDbZC6UBL
tsWJMpvt7IpPhpdT2qjWdN8Goa4rz+dAEeiQA9akuubh/ahHmGXOey9jbQANGHXkMefErpdTVbxS
20GIn8cdSMcG9bYx2lIIRV0t4bLT1/0/O2wqIj7cJSHIj6u5KXc1xBEm9D1lTXAoVjB9XFbFLSve
OVsip4gu6ZgU5UnSYzMVLKO+fPIOi39FOWsfvQvPcJe1rEqg8kmEWO5R6NIcGpo8WUqkhRz2LeWZ
izeygL6B60Y/NdD0cBH/MFX/kW82qCgPqEq4+dFaIBnQrpZuaeBWLcyLLXGD3qikZC7aRhvoBSwM
K0TFUDS9kKDGR5rNl+P+ZCz9668aQmIcJsaDkEt7ji4gNghU8JiJDpgGKHvzuMiYBLtrSH/K0EDb
wcIFi+WH6Rb6pUMIWFx0hGTAhZVh0Gw2IkwYkrdv0m9Kn4fxEwIYVAmfnNzpMgC23KtXy8wg2Xa3
GIzjTgbEwpKgCoEPTPREqU0IyGElzWET4Ev/eI4TIUIRLKa3W2XJ9tn8torXxqJJArOxVMIrtuq2
uGJIa023aJwZb+0Lg2mmX74GIQ7OOtyemLY3vdGTAkGoHbqRJ9e4XZhy6ZfVH8P0pIyBRIFB5w9t
Vn08y0u5CSpWOW6z634MSxolccifexiMvmPYqatznLy2dVvkxg51BBn+DgcW+62epHqzBkbK80Mx
ukvK2h3rfOAPQf2C5+kx89x79M94AyEzZn9F0TeqK6bIXos3Xkje3Fc+UDqJzYA8iwopmvxPf04X
WA8yltcesC4rNjU0v9KwSzpgXJZXAy91ZjSL7QsnY3JV92ll4NzPiZOj73qe6kcG3Bn33myiotdt
ccfclXrT0qIFRjGZE7IYiBRjzm+aQUXyEM4A5f4oLHdmjtwptS8Se2SPPCESsZtvjBTv1AGQmN4h
tkhzRvRXoHut68nhzb0t7U1gI0CTcWhbY5zsOmjgeqTst6UwH2iyQSW2i8oYq1zyTeTWRq2eA+Nv
XcfbwZPdDBra6hua1OcgwR8u/eAw7vTGCJojUmK7FZoigtGCyENuX/J1FLNVatB2JwQnfFqCZfgT
ICZ+qL6b0HypFgeKxry1EdOkAqbJTpaQ95jjqw/2MST/zz1ZGqIeDo4JbGqTYu8nE0vFjkvRZudz
Rv2YckczS3iArXJsFY1n+11Kniuz0MFALRshTKfEFjpiCr2FjWECmE/CfQhIUW9SleGCGOJckNSU
c0E8/cUzE18c7QvRKaywp4IFbyy9SwyxN4MzlFGT5L5BMs53D6TW0byRn0RsYoWS7i41DcbHU8MR
ywXXhblDTN7P6SYXv3HtEerQoOZbWonUQWr22VS9F6rpt7qxAUNwAqjRiqO8rLBZiZ7co3AyiDCv
mGRMQT1fNvfi/iGd0bNSCJmMqQKA1qYFTVhfAu8jb3Graa5Alyxbp1AqgHHs4nVkSOVUkgMZyQgJ
W/NmO1cLm8EMopvLIhPxA28yXckKAeRDo4qlzCjvuULnYqGXMuVdbcTkTMs9Gbv8SNT1ylrL+VSR
xWNlOQvXHWd/VjyK/HuqLH/jQLr5Os+VUGbJqso3NKel7CmYwYJgp9OP+XROd1k55IXiCEZAEKuv
Ek2A3JBtm4egQSiQl3/Prvmcz+aYHF3REPZapF7PNe0/g9AT39FD3Ln8l0bDYLP3jkKkAtLhI2KZ
YN/aOP6e6cEsxwcpE4u1rvWFwhZLVaPs/5iDxOORWDXQOq4k4IfG5vShNP4CZS46eTE3Dt/y7KXc
40eq7jwjLcMrlZr9A14K878EMfKPNZIGyhCe/wQrzVJyQiAwNhAHSdjk5QvKybAOi+v+eNbLZAnK
zHilbMQFMEe7ldCdZegbozB1W8q1ZsJC8ON52coKr+Y+vXZsaF8btLb4DOAw5CW4yDMbfnbnMs9j
WHHBQLeR/svohG7cSdaYZ+TLhsBBDjqz122pczJcSiHlr+5Gr/Lhr7mFaoE5Eze4GboI+4yf5WAA
zc1q9lW8R365NfjhwXyN3nZfqhPVp5srg4cKCIWdiDKMfVqIGI7F4gNeBJLpIg7ysbwjyco23PNT
jiUHptgQitEch/Ii1mRmKWG+1Q/bN1VMYqEvgd0ygxeo9Jm/5CrC9DFuSJfqqbgsfSA6gBf9161j
D9HYHVcEhWDzhjxPz+DsVbCP2kpIocNeUEfrct4kcIs+R/ycdWOdvbAM1lFZl/rmABEFQAGynPCC
guXlRiBemlH77j10oYM13491YGj7Gl3U8Py1jNgEn+Qnc71/4F41YgIwXOLKKryLtxoLfzjGGRbl
CG7NqoZunry3hsaGyWky3HxllJ23A+hL0GeG173y3P7Evrl12lz921UeNMxdBcKuNgbNiXOKe7PJ
LNXjO8yRT6xgXzkLaU/NMX/igAl0s/Eaz+YlisKXs/q5C/JLakUTVIFmCX+kCfpqQ4trfKXCs3Rs
NT1Zg7gMLBEfpqWe9R2kB7ZkJTPnxtZNscA1hWhvTO2Edh6KMS+Hr1gszRHyCSO4+FvgGaqlS0ag
clZg1WdAz+GA0TigBwBmGqIeola+sT6drRDBfE/6s9LxT9JZ0opTuw52g3DQMI9PWs+IcdyRPlNZ
AHUE463dWxYieWGFw5nBmjM2RI41gZeLcT/5ovn/bHPHSZlUDZBoSG1wO6kesQM0Z7EGIxxeH8M0
66X0Lxz/KAOncxYqKmpHvMTuhbA2x7FsDlrmnSHTpdfqKjU2IVsYwRvd6IbCM8nAmIO8ie5QzmZE
QE0XoZk+pHvMGtD9ovVIhhaMqoPk5OmMBHPInWeRAHQkV1C46dwiYanBkJymUkdQomGodrs2xZQp
cpsDiBtKR4KfO1+7wVFzb5WTQ5rfAxuBnTPWFdjfxqkwtcpNSfQY5QXDUScgtRoq7J4WqbDcKgtv
S5lR0xCQ0ELPXMzqaqvOkAUckVs7MltBSnOaJzYElZpeUrx4PKSBdz5YmZ6gbE23NBZE1cf254AK
aDDgVXRuH99W1FTrvWpQ6om7CIp5/5brB3wa4BQeF3xUDsyuWa7l4aHK/BuoL3i7OhC33H8BviT/
6iLZsbULNVE4vcOFG0Xg2+TsVGpGhULMoqzq6j4y9LRZNPNQqHDX8MsnWfICp58uonFwBkRFPaSJ
15UlKu5+1y4Y8i+UhlzuWe2qDY+v6H8TEfWAc9ViYFSlU9+Fi96eFehN4n7FgrurL5rFgheFSjW4
hnEKJHzXbrmn9J10IwjAu2509e0VzCq8++RMHsYeTfLFjxK9uW0AweAlT7BbNCttCb3bmbx6O9VO
vQ5Fd0RGtsnnQoNnyQqCQBkbCIrCiaqOce4CK4lkkXvXsKM+YUNFxbAeMAUqCX6OqbvkCT6OHss2
mbi0vQ77qlisKsQ6BpMworkLFZAHDyNx+utESHZroDSLipK+SvXDoe0aVaq8v1xZissYKvV9H052
xX3cPpTnME//iPBPFxkljPejsd56rJjolxQweLq8CLASZwFlD2yWZQR/kPcwJd5/DPHszNk/OR17
a//r8mnW8D3gofSiHfzovpnzWaljUSrtBVmm0z0mweZXm2vKgeTm8hUQE7r8XZNCGnsQHlIj+lLf
Qs6AOYIsU31NfhxlonDONrURnYWOGeIz+6AWfaArrWBbyHmwlxUiIs9ysILDUyg1e07+TpTTylBL
mE+iLO34gk71eAmKZN5f27sCnYNgdy+eYaeSummEPTUV8bvQYL3B/DmmdGvGgz56AZ0mq7LR3KUT
X8VVnhm7cXAtAiU8CVpLwohQ/Yql80D65BYTbZTWs7Tgh9t4XckaturcD6WhFniPBDqbbmeJEbKR
SPC8M4OzpQ3oIPbNfjDR5/m8wLU8fNZdMIaqcZIkk4/UlzZ3aiw6QseEYeBYPZCJXJbNF9CERhm5
KHP5NbzL30DE7sGMQXJMqr2GMt3CskJguwRQQKF0snK269UbENOorCLdzHFh5vg3r7DpIJ6xhNc3
C47tjayk5ZExNK3+I9M3/M65/ySVAu7Cy8DXe39RZZ1cA+GmBhNzxCBGFF2OJ8vjrMP1YqphymlS
wBgjroCuKmYAp9u3k8TZdIle4FVw95uCJmVxz28snl/Gl16V+BeRD+2UhC2z3Sqlq+9L+wsGZRbi
y2yL6RKOwZ1WUpxmcZHXmgpAk62ioYiF7wYXtgcm7X22MVzIipmceFLL+f3M3Tmjv6Q8sdKlTUO3
Fm2sTw1Kl0U3bcriptm/zAdzVxU5rQ/pBRWTu7MqI8On2htFryWAko1A9RqDpLTkeIPB5Ef0PPXb
gFyewoD3nTeSQ3BNnqyohPB315CN0RvpQ1exVUQKYnkbsKGSvBh38jLZGx+XZ8AWlgI/EM5JFabT
JHmk31+UO6xQefmGT8t4WSHmdy+aH2KPfPWntG65CPf/8MIvgwflqZ/KKg7n2fIZCzlyeW99q8KH
Iew6hnAgFhkpw2DAY5ewSmpFEzo2fKd4TYd0u3CV3wAGCMCPJc8VB+as0Hu22nvFJnE7ZnW/HyCj
SGESorfnWlAOAEVZFWYHEzP26U+7rTN01abM2AxKJR8AE9CuV9cSer3YxVuEjrkJqXRCrgc8ofSV
dypAZlzuDCYDNKJ2p+EbOFj9TQ/KK6o347dROlGabcjhZn+Gi5XuWBfg2glpQCzk8K2B+sdZ9dTK
Ah9lhzY6LWg+61l0WRy6Us3APSbW5I6RAz8Vh9mWeUJmHlV732li8SHm0qAmwFslZM0QYZ/k6HTi
wu9OChL46BCfHmelV1IfrZe8xKi+qygcDoKxrUHQE06iUpvoshPOZLKRUkfIylwKuNUns0S+V5ft
ZHrhrjFxqE7MdOXUJfuVAQxye8avXktD7bI36m4Cx9L5M0znWg7rbJthx7wpbYCkUa7ujy1Xc0BA
Bhmgii8tH2ddavB+Ssx+VrHLYGfi8xCOcGB/+zZgPu/5DZ0PpINcZzf3GwuWM8N8TeQrqDr/L1ZK
4d8erqiQr+12rWXvc7LBEigBSAWfFPgUo1PThIRUlF3yJ/bJ6WDWhjYjQsNMmNTq9x6bWu0N37Nr
0oLXgtSaUSffIpqlVUgsWFaurU/mMaRJj9pjbpqtmdpjmUtrOTY/YbM44U+sVYDcwPv3W+inJ+Ln
6vQtj4l2ivVky7CZ0af3PkzLAb65essfrSzNV9n0A3SIWqHXRt/XHH3MXIDYb4rBv2uvFIxHavnW
zhznsptllCN0aYu2KA1TyW0PZRwpwKjO+zwDfx+pUDzFPxkqQnP6natErL7nLX1U6s0X95MAogZI
0EiYSR0Ahcxjh970u+74ycOdsFR4c9+1yZJBqz7oFd0a+IbSSVeeKZFOgTSxjw8cNwH6CcJhR9tC
X4bOFy7+HtQjThqVQsu68eCtGHcC3OSHsT3txjTcUDssFtykEjwz42ITBBIIuMSwT7UpFA5ncFll
KfMG62l4Rm6boYvfv9+VwrnXacoi3WGOf1f2WslupkWLLFB1DEM7dBhkx7DcjDjmM704R/eyCyqh
kO3qa4Bd5uoqI+E5fRITHCps3Dox9MF0wgFE8cM2YaUb4h3XgH6na7I/5bhWoq+1yZXVj2VjNQwa
rchEhTOej41f3SMhbIpJGCzU7NMMYMbf4yeaVyQ0s/w+n+gKjwEUS/uayUkqN0TXg6EAFtfpOqwD
jT6Faylf4hHlKpp3UoEMiigQcYQBXaSQHDfmd9X/rqPMhtjsu7zK4c95Cdyuv+lWhPC9x4a9vbPk
thsYWGOzhJNn+kFZ3pR+5FtUHk7lWfbMSlEqGSZDN1E8mofLd5t1fB97ay6H5UmUnOKEnTGuDqpS
7ShAjke9azq695FAChl4HA5Ox5iEuh+y1MYjPcUr85t0qDZmGr2X5QuEmfGOv5HPOFfONBpxZJQF
tBoSu2IlwP0HysLMzBXXl10yIFbKLGDbJsqEp+rR7qWUih4YTR6B+zJY5s30LTjLVcQy9MNZbYjN
Zbk16L2/zK1NArLJ5WoqwxOREG7pHaT3w179mf2hhhlx21jFfLfvc98ShW0YHUJFc1u6w+bijrS+
tXp4iEz54pUMAHZRTM/Yn5kFkeq/1SSN5FfUhQ6r87sGHJBcy3r/cvPpzilUcMSALW/Rl7DsNQLi
8xvf4nbzLuCiety9OLCRUZFDgwruiQ7m5zamgN8Dkhgm/E3X6tRw02qndC/cSPH6PUr127QdfOMH
OfXfH4Dns0/Hua2r5hY4LV+g1VDlG+PFPAnTlgu/8vcrS/A82qeCt/MzJkes2yGZU7jIXRt/YEps
4Of+S7jwLz442BG2Ce9mkSAFFAenbhFINpR8JtWUF5WCk9NB9AXbaFSpznarl1bZboHYXaF2COfq
IiJYGNGotK4+xuq1AFAjCVFdsXaaSR/vJVlumEat7+4GGOCllLwfoa34ykZBLJqwR5EudkCb12J5
t7ZmjUB0+aTgRj85SnuoHMrzbMSt/aYd992i72HE6H930iYarjoTFQRAbq7/DqB+9SQKwD17LvFT
K17oYleg4WiFpmZsLfjppbmuNjNMbDq+EJcEh9j8Cd00dYXNLw8NpX3HYLwkN6UpKekTHMy6Az/Z
/uCwGcQMnI9rT4SjO2oXCDDrd/86/i4VrFVCrX4lAJug2HW/kAh6lrE/GT4vVrF/o3jaPuUmhKoW
e7gcDurNo/S8Wqo+vgUOp05k3li97i0TTDQKKE3Vr+HN9W66bQmhC4gGwuSmLGZi19an7nvegzmf
2WUMBdQZyY6ePjOcNFjw8fzMDaBaGEGEQblKF8DuoVTETb96WwT0na95bjJQLMppa7zNMKwBmsLe
3BQ8FgWcS03eMO7aPW8O1ZCKeMvJts9p8963sbVnQcESYgCXamrLnOrS2wfbGgpF6LjFdw1oQ26C
0uEdfSU/UPSdj/ITJAF0I2IyaVR6di5LyDSL1bhNmvsZlBUtjCHav4zYjx7WPSC0MIiaw//DyyzB
APerEabVf+rFpPnxmuQ5ULAHEYq4nN8SKzzExz2U2gcc/6pCl+ibjDN89BTySPZYKMFNeNXTS4GX
P++08aKlNEnDpCJB4butd8l9Nd4ZXoqQk70HBIaz4UHTpkwmBq89DB3/eJ8OL1I3vbCJGtwM3oYz
CnwMi5K0nQftgYiuPrwSZhnUfOwcY4Vj6NuHKPmaBa7nAJVIoJaAGyHnY0JaetZFJoqJE+tYqOHZ
wmg++KvZcaIr25EmDZ45Creb+1CoGJaSkP7Q5cNNQ5W5Hqagn4uK6tfikwFl1RNqj3/0xcTVxBGp
XZd+D9sti/8XTEa4XkOq/zLcJ+jPCP1Z/S0OJhUaSg18AvyBQjZuap9fqNtaNqNGBYl+MQsKMQ74
qj7/aB4lXxk3fXBXib+QdXUJys/zv1P+NgtT2LjqGKWbIbRsCxjLmdgEnLTD/YXnQK8wQmqh8GDd
+YCbxNn3cOaViFUDnEXYlh2atvl2gnJyCF3RPEqvlphFClgRBAb9XnMm/CQI0lE2Bw/yS/+3twx1
geqsVCEn5E9sa6ATb7k2/4JhS1Jnxj/yhr/gh6XYrCoJS6yF/aEEv6SqatLqZYyUMn3KmDQgWinr
rESLVzBN6kKC5OIu4wrp0hMe1Qa3WfA4J+DbLYGfC7t4FSzqN0FoLvYupfr4YfMoF6RmJZYq1WzF
lny+/9EfjeyjEfR876P/LmtIN9xx0Y6i88NVhugvpxJ8GBMY+fA+tL6jOZbFwuxOUVOJSRcfdKFX
FgbEPBf0hibSEit51j0yQZPt4nLDnsPvH/Ew6AVXp2tKeFcSsgjNZvrv8rpzXgHCGjKgO2vDEPDR
BxRXi0wjrgYeq4xQ94MQ4u/QaMwTc3Kun3IjyKQUsJPBvSHM5hWFf6HiBPttLPKW8DDptrbDPj2r
8uQvTLYTpDEC0YrtpRL8pzmN3dSZr3VPnVIe9dhCjVTc6ESml4e1lbbxCgHmicXhYTKU2wbGmD0z
P8fg6uaTp7yvAn0yuqdBTRPK0jzTiRpeK1djHX7qzBouB9NudBu9z0X6xkqU3KIzZwYjjRyXfI6f
uDZ2kcwZCCZ+Xb5HoR+eBm0Bl+5SGyLWhCwHVqpnTlfi2IOX4bEJyGod905wZA/26OXYtWaQm246
+JnC+FLonIMcjEcrftjbk9grFjDoS0XfxTSgCvRuZQIpbY7dRN+9fOabm3fagtAemMdIFzEDpdr0
wiVoAlAtvMeQ2Dgn54Alb1IDDrWdnz9sZ93DXdvPCcyAtLb7INNhxGvq+qC24n0lW1g6iewuzrsZ
dq5r5uE1MSpMqXw6pF9zYd96oSxKA/Ggu8U2PTcO0jSFlrXo5pgfXHpxMjXqi3kYWj8S8mqNU6UH
/qYED8Hsw12GcVa1Xf/4c1CUoUmCkDkDi0MOEpp+u8RBU6X3+zLXaSlmLuIxnsxrEuotrSfCwboU
UD4aMseCmnzcMaiq6M1NqV8mZq1G4QwMhM+ArXSuVhGGui3KJxySxVyJga4taRcB0cmqKH9bwvqB
KnuxJDZE/PyVwz00jrD15qnSjwZOqwATGSt7MZv8mZv4LgYmAUXfDa0VTjORLNQYxp9CSgeklvq4
vbhsFI8LQc+Jt3jgZh1IxI9M9oPrRAxOtc8ZtZNXzbaMUMkekvj4s2Z28jKPy9q8mYm9wsq2+BNk
PwRB5AmTw97qAdFXZzab/r2rVUXNbec5NbTDGkHZs+1GhYFaYbkhRZPuiBg74blblYVd9LLsbzrp
R+J48ZO9bn4uE6ll4X9xbJtn5TdZmf5DnxeFC62XUXClJY12QZZ3X7lcTceJ9EcnHKP7aplAuKOp
bORqXSNB40XBvTu53QwRgUGsypN9scVpAiDrYLwx5iLlSTjhq5DBk+QGJqAK4nb2ixzZPOOHC2NW
1OkWTNXECOA9P5GCA5D/k/Hipd7GDexz19ESNt7g5wihfUwa0u9X1s586tGQbiDsTXtoN7U08s4w
FyaeXNChcGToOH56Io6EkwC5XwhwWzQ1xaVjEF52era70Wwk8ejj43rVa3M4FSgAKsHqyl2y1JLo
Ush1CbzsP5dfkp1hPRJidEGACyuViPfpwXHavBLYmqoDIhiy3bW8iT+HBndSGMnnEQ/yUf0q16d1
bUXQFpAl/qEh2nqiBrZpsRF4zCyG5ycOz/agNNS5boZyknHuQxi0FYevcg5R+xj2N3LXtBS/mbB+
/NHy0OoTLUH9l/puA4/KwJg0iBs40CKBVlKr1rLXBv7DlWGD+mNDAP1dKeyGxIeCzIHEnbt7GoH9
zjZ/PZT+ADbHdWLWlQ1GABn4CL2eLrBkv2jb2MzfS8e9qw5S0vdP1Lldx8+mvyzQe3VU2GkLQZIO
ga8nVyMZQ5p/AYKenJHocsC+iQGtKFUYaalO5mbo/9tNXD2PAoK0gp3clPmxkk9bHbxNWr1DTokv
d9XkdL1KgGAVIuSE9Q8mXRwcj3kCYXDArTnnE61USFSByRS/IDIGJsUM6jPAv5HiP/RYrXDsOI3t
oLInPWElErY7lh6OjUHIBytoo87iMGKiz13M76AArkwWorbhkNgelpXjybqJaQrIl31daj/fCnQ6
S1or2NLJOk8BkYwPVI3f/ZuKb5xu19az/5oESiQRYmWe/LRjxIwfq5unKJMM2OQR5hMRwQT7taQC
Cu5MP4A01m3lkJooK5eQ3Phz5oL/Zpd4XjzKn/0/Q6/5CLA7ha+aqjzvyuBinuyQV2xCsFPuGss0
q/xYnp6tkOPqV1sWMb9inzNoFrTKxVW6/uXnScg28ClExNpsakFd1IIQn3X3Iw6IEtU/dnp05guV
MUYFk9Tj+eZlYQULKuxRuVnJfntYz1dnAATlmKqhBlo+Ioo81eRYv5UjYW0pBJSWWqCunv33+6X9
ihgbWsra+GLme8QdR1OPNxu7rD9nLFC9p+Hl5C2dOClPV+SN+WCStaAwm9C45pDgrO6Nhi1gocFe
N6J6xtkHPj7P1uYmg+Rdu4hcanxKgyatpGWUnoRtUPeHhcaFtBe2WoGwHGTEYy256+avfk0Nfnfx
RlwOkwcBW5cWMRvXCa0d3IOryeHdiW5TTTVbtpBkDZEo8Uh8PQKWEa6j/+RIRbXI+6oYv+MKYyMX
oAKZlyTgpE9z5aow+htlUnE8NlurOnJXuBDMButouhB22aS8urNOEJx2eX1FwnQugxvQB6070uhU
whN3z1Gr6lCtSetieezQl3bMU0sjhgMRuxuXchFSJ+tGcoBHbCzu6+maknZXRDv6iKWpmkMzMdph
lTxYCz7oeaGjvW/ELsLSndjJUt8Wt4R1gFw/+xmKvsbmkRKaWH7pABDsUzTm66A+vf/drBdHuu7I
dSvzxm31nerkM3q377Dl4fqdVNpnPo9agJB5KkJ6RRmOLCeuCdTAaEo64xWbl+H/BdCu/bmORg91
Me6ULX5FUdbuET9Q3DPNd1JaqBCJRreuIaqmhIguF+IS9JpVcXq07XGQ5nLfPxhiKU9jF/26n7rR
GWYVxKNRQrEoRA2lR0YlqeYBOdvBdczzf9r7cY8+lrDuWuEGKxJ3xQdZLg0D6OQ9TihamfgSxtwN
5O0h1uWUn0IzciGwEk9pIU2DrFdZ6H2XXVYNEu8p90sX5seIX+b9s94vBtH/X0gZGGR3NIOGzYHt
dNdhM+dmR+0zbYBtY1PipXs8I8VcivKkx7idMNUVqmDvEBwHf+whEtJAIBtj1pfTwwzQ1bLtDs0p
H0SAlxRNXBF3Q8fDxdEiO6qzKfVjhReB++k1Ak2Fttyod+q1fvF61AavVOxfyBwmzj297rpRcE9V
kmUQxan3kWT6GPeTDtGEBuqsLKNB45cdbmPKzBheJw1mISohP1AMJQArIvPxm7+5Hwjrhv/jkcSE
dXFIXMy3QXxYIedgFI9WC6rjQQi5DNlM39PGhcbJztUT6prvIRUiznJTGNv9uO85sJuJMY4uRkDK
pOmXIId+MurlFGIBg/nB/J0elPVSxTLi8xmXT0zV8a7I/IaeVvcg4lIfYFRRfKemhtBupcg49Vt5
lWrx3sfCHvMC4MhhrBxNdnXyB1tdJQ+4zKiTgz7IN8quvxAeuAof8jcBnP3eYLBZB9D7FxRJjeyk
fNs1mJduxlzkf4CMg5ruh2yaPUwg1oyqKNensXq+YQRP5PDkuWPSgEdIcvlKPWkGXVg0zx7DgJqJ
9125ryVN7kx8PiSwSVc6BNguECba1ktGARNlKmTKxYi4iR49z2Ic2Rdo/cpWOsQQjGrcbEt4LyqJ
pJSkbklpV1UoSp8ihioZHFaDpXIyZaFjl5nyaBhmpVvrCZCBx8Ow7EDCTX03Zf4pZxzU2q6Zw40Y
8pkcdzYRPhHIivDDfPvAaAFrFO9a1hu12yDI2Typ0isAPaHdJPz+zVKhmlnVQa7zrADaB9Y+fyTo
9Id+G4+xtboyZImUATm8LLtdgIFwOFmJfqZMRSa0ua9hs7nTnUhgXZcacVdBmhIlq8jA2ElCZGtG
sLfYP/0Jg3coTuRWcW0QINnxQh+OwYf4mUMIhxBmSj/QjKCzrbPOSfVNj9nl/6r3JPCGpnetD8Wj
uTfsOAWd71y86RaKvvgNXLbOMPD0rmxqfhbmS+uV3O11JfnRsZAs1+BMJnXh/XbPkIghXcmpIopu
MCikfCNAmc06JIqLKFhysk1sUmqgw2Z17KbIrZ17+kzjRhyePH73qgPu3yhO9Hfvo2dEi3JvBMpx
6078cJKfp7eSi0qY5+v+g1mSYwrXLO+ZqfHf47GFyuG0lsJp63jyIpDuMNzx+QwJmPzbuSbvjBOJ
+IpklGM7KUbXCjlVLNi828iXzK2nQZA0eRwGJLUtFwV01QsDWZssx6Q19zoHzcaIrJ92VIwl8wW/
S3kZeIbnS2lwcQ59Fc0GRxoRitwelGNxxnr7Z8uWq3aOYRI4Vjh6JjSwtEQw7bhcndLMwyvorQUs
6C2u3/tMtHpRXR0dgA4/b1fGIs5OAHc9dJ/PZ9ebJqJDN/bXY04JOkF+uHSa74tu9/6o7BNkhcQG
N/CLW9RX/fzAjKcnYS/OFOGv6hK7Lv3lqyBp0Doz45fmA/XK4G7AAHE38cGwqAWmrOph9BLddEBD
VaIqyPOdolJCHM1sKb5Zf8JnHg0Uzxqb0MvSwT9ogp/aBKsStrm7VBp4lJarbcQZE8xMd4pKyMDh
Q6K/YZ2leeKeR4lwLFqzdeb77dxxReauAZoIzAzhpOZnhDOCDchKhUrR0rxgM4w/5iP/ye5Xgpx6
7dmt8omL0fLN8moGiglnv0/xv36GtLH8qQkFVPSm+rYWWZtmzHGZv7DMRmDQ2ZwXH++NVCDw1kNv
NDRemZlA1oB4s/3HGtchlDowM6Qo8NZqdWWXWnaR3MLLvJl2Gn1hdq8eYhGfBTMO48QtI1e1+MLa
UAbJY+k3wibbEk84vuQmlm686j8fo1eTaH0++9+1sg9FFprNnxHZJderFPP9p2Qq7v+nIHwe+LLv
E1xn91UdxcUs/FQrHUKKzhPFA3OT/8+eJjnRIQEfzc4fSRcONuZLANLUul/nOnFqDVJrkhaaMA2b
NW1mhmILC1xW8m/Uz7w/ln/YcER5GsVED/LuI6J5TQhQJNesNNO+GMHpqivmwH3Zw9u91qm1N5oz
GrkUCNFGOyuJIJgjtdTgcC5LMEKUJzFD0qJfZqYLCemNmvkn5YfS0xEZfE7ZJ0PM4ssKp810pEcx
J+wj8jInoOfMfi5tLnzev2UG93xihq1+ZhpDFH3vHhOnKHEPKf93or3h6Ky2VrMNaA9JCuIYbe68
YbWwr2WGcO+jZj+LEGHORdqwFuPAkjDHzs+KdpGizxRJtooGS9Kx7Rh+/bfsWZ9G+xMECq9r2AZF
vM57QpGBcZSqY08E5U1UNVWDH+/laCY6HtV/f8U9I46JNFGztgua6osX7fJ9Wdu4RTiKrpeXMYYx
VLeoBxjmAQMePiMKPb/gKF4/1a/zbQuzxnkbt7cjyin8v2DnVz3DVrRez+ermu26kZ9Mej2IzzKw
GMuUxiLPXWPqEb3Dl1hvpSyWYpaXF61mX2cK0xEYUnIC1p0CYKsoszS3DbUeNSTUjf+zF/HpT8am
44xnzf93D/cu3Kcja/d5S8Qd+7tlRm9IzJaqilA3IrcfD8QT6WTSk/TNgUmF3aZlSwt45n8kCXtg
1Doyu08UKdf+UxGB1IwXIEAA35ANqfnhZTg6XKxMVpo+syRO60ko7oIjPbH+ONNmt9EQ0l1GFfg1
m2nUzOM8HtyXlwgYviyr2s44FKLTFRql4Dcngvmarn8LyndWT68C2oGxnhYnqKp2dR8YqyOfEhY2
5vHt0T4MHwz75M5adpqJUseKnyejLwr+h55xNHjCbNy9K61dZ6xmYUtE9Z6Lk71wYQJbchws+MaU
ti0Uujtz9+kky49sQ1Pa0ypb4I03uHiehvShDSrl2WicSIOeGgS+VrDPNY98LV1EDucO9VwYzPEz
1c0eIYYryT8KM/agv5Qz9uUfvO6I8TkYi8tTX1j9NBDLHucaZnu0B+DOU6dJUikcbYQW+eiOePhE
LQA6GpbSa+BTyO2tRn0TgFCrKHamowFsRywXjhaxWjaJg4L8aPTbHBaOZpyHHxtjGNMNwrikFBIj
8KqvnoIUCq8JKBRl4TWhNgf3QKJUOD+ECLvA0pjEO/nwJfD2DJVuDeqyKf3DtyggimVfuGpu7wDz
l8j48OMJCoEmY1WuRnkzVs8fHubXLOkoQ1CawMACzD05p/QoEn8Mc5s/rRziLlIsP89Yh4+Rtahx
fpeHcrCSO+joZWmzV+Sm5FNVNbSecGOGcJWdnETcCaOxTn1TeibJ5i6c0BUo2iQM16y/bpy0KtLz
7qF6yEYzKBcvLSsCKKxD9ay+9MJLFLmmdMbBOpuxxg+8umpvQerHBYq/7b4F9QSHt9fIZO2tn76H
3i1JbE7a3CpvDDOVY53pwvsy+PP/Dq3hvG4tLFIqKIiExS8YAgOUyi6kEzcvDjaVfuto9ptR2KEO
nIC1QL33XxR+ssYFegfB7tue+y6sULzUR3oHHKu9quAnW4n5odgfVqT+BKH3XK6al3jQfK1txE67
/TgGEF4mMiPp6vMR+BaWQXZ6VtS4wcSD1ywn0fpox4/T4fHO1IC4ioYfJ0pnNIt7Nhpb0IW/sn8Q
vwwuVzTbJf9Bb8A0Mc9cNTkV3Qfg4OOANQ3YSkOb6enKHc/iSgfiS4l+f2xaWqGF7xJU1GKS/rx6
3RNggQvAuRb0OsOD1tqUyCKlkTSjXZmNu82DlqH8ThqusLQDiXbv6LE5iCyR7mZqD8yw+BCzGhM2
2YNovLYE15UcdfFjoQGaPg3XqUmUWF4jRc2dV1nq9pVd9X7j9p3C3PViMOSfzjgdcOoN+J9H5gQn
Bt2YzLrAUNqIoedkOKdt3wXEBWqjImAosQzEr9OCw7O7OxCJYwzs278d+7I7q6jexKqDGNk1aj3g
caF2gOykKJxGYutZLz+Qp515Eo4jBi8q2aoxQ8OVXc5RN+cA4NuRbni9XMzaOR0yNJRpDtuPjCfw
xLsopbCiIMR/eRXZ9k4we3c2i1g9Y/tWtlbydTH7bd1oUNJjAV31/Jy7jKA7/9Nv0C9/pzGMHFxj
b5iNBi+4+HPjiapuVgfcMNiC8jIS6GdYmGQsPs3pKC7cijXkUJFr9rrhnpFyKx37hTfQwG/T0jAU
rX9w/FcCDfj5tRo1wRMhwUhZg/ud06QK/xKQ4oFbkC+zCT+RSKbgsYO43AoFXRMi2ZNxJKH2hagJ
fhntFbG0VyepgGftloCx4E0MzigztLhfPZgx7L1WhvLOCFUo3sxC3thxdzSzPzUXqGsA4t16AdLp
l8XJT0OfX+Tp2ZFEbSqENdDqMDBf4CmDUX/neUftSZPseZmVWS5e33oH9NTW/IgeQP8NQKFmhyLM
ECtQI3cP43+qlDZGt3wr5dMa8QcxOO1+iC1udqah7fDo6FEEVsWuN+LAmW2JR2dfDPB3dVTfuAxu
ACIDUzxxxH9zNyVdJ6IBDgoISJSvtdNk+DE9y64YIiVhwEw8Ace29uFv/m4sw3xsetEouupnRZ84
7/+5DtkPgMyhku6vNntsEszmrbWjJhLFVPX/1Nk7/AOEU8+gdrhQJZsZJp/szUuDO4uZ9laKaTLN
Jo4vrpbs5a9lH6tWG3W2TNqN2QMnxu/vFboQ9VNljYvLOkyznxNXyDbwyijKxB1B0rCj9TsGPRNa
68gd/8WMlt5pW0Vhsh2tddOR8p3ykx0OCSRrQA2327nTfuzpS3O0neLlr3dwEqeU1NYhJI4qg+k7
FDmz//+JkV8N4K5LY+01ce0w1pPW2C0FUedQptxxsFc1v5Po4MkPj8R8Ke2cBb1m1ROfj772o+9f
QG6sw4Z8in2Jrft/FX/qREmWGWVMKVZB1ZYH1fs1FLstvpvGI3Hvz+jFs6MSfMDHkxJ73G1+Yc5h
fm9wwtz3AcW1kiFYJkkRHNxQm/8oN3K4S/QHGNWE4+0D4bNNVMHVKsj59WEk5Wa/i75Fj2ez2fSR
NyQH+pGG9XUqmDrVMSbdBh0r69V7Ta4wyh9lEqM/FExjgfYYba+76JUEuhjP5qMdQaSm9VL1ZZuk
2IQo7dG0D74sqCMIXAmlTE4NaoXVMNAHcuJS4o7z2EwGzgRrZHxermiTDbFY91uIRwkHW0szF+Sz
l2SwepzL5dZRguwwQZvJjQt/UkVs+3TtmlVcsDXv+vxUewa631t/l9sBgybs5mEtswNpIV7oi26C
v//FVQ4Px+q2kJT2fj10yaULWzSR8qNw+vae+ceLgW56MyH8RWo8YPjHPFZUk8nl6J88bA8gdYVF
5r4MrAahjIKNyeRvd5smLm9DJF5KkUA5HQWaOTMerRIvnWRQm/8Rqn3rVFSWJTTOGrSVc+5+a8bc
CQ3Rpajdasr71dkfNDB3jFh1bn1HRzRqOqv1ZvIlR64kG7QmQKT7rmnUBJLYz23/qf27Lc+TV1Vn
39fsfsRLdxO4g6Xx4BI3Bp4/Flzacmp7n55Wl37JMILCrs170VljnxnoTXu+bBv+hFNaAZH9BhWH
4RpNDAPTYPEXWMR2fhqBRa40wMqT3fOk6Ihed1SWflzxEpfUi3AuAXk9+YUByI6LfEFFGXYeWG2E
Af6Ke+2bjD1kT8kbqU2uQp4pKyfY9LBGD9oInqYAiYKv9RBlwV/kBLxP39NyN3FlU5yY7/lmpTMz
YxW+syNkT2d7LM5YSUii5dSlO75wwRa8+hWsL91yRlnbNWFG+2pqrypAEaPPUsB+jYvrBbOFn4aT
Chc/W6MBRGRZfwffYElRT9ayCveXAdgc/X/XSX4g3m8qfzSNnvLNkF9RAHCANnxnO0YjJZNEhLQi
UZ6eKfSmCfL+BaGHhG4YSnZuqlL+KeF+6uHkXJY3wJsIuRbPihNaoi3tK6pK//GLNQa5cP8bDDhz
4zLnQH9apkQmM/19bbbu0X8NwEyEcqcZv1DPB8B1WsJMLaMmmeNGGj0N0U96+wWibWn83h9iKARJ
Z7uaYkNY/MtE+tycXboK97YrTFuclJ/tkK5RDNaoAgy8fRWcV1ZrS79TssK2tgbftELUKdj0Q3vg
XHPMxI9P+b+qFuogZ8/AB1/dMsIvWZQ8SH0FphSd3EU74X/knX/5NmJglIW7GMrPwONkvnqVmeyX
evHXTj1T127mhoCtLXP1k17peJMzGIJPpTgwWcTG37/N/2pGBXiYSwnq80xxzafWAb4dLVNZWBgy
oD1CigqABSnBM9eQ8Xg28dtBypTJzaZxzJxQn345sWFgtfjvNvT/Uol6kOvtTnXgyq/XcZFQTu65
2iYBAy+PbczdqiMTFPidCkI5leF+6eFr2rBoDE3+Fc6eWXi8dubFuo34biUjxYL6KozX59ChUXoa
A4ZVfka+/hWFXV25Ta2MxrtZ5wa1NZMBMhwiHb9juJ/PCNtX3BxZIffBh5ZFbraKQ2qMSKz09YCh
fGGYJygmMieZPIEEk9h1XuDWOXQVd+H26zCP4hJHKGtS4BRUL74fd7msO2uhbjKNKSaANRwK1ZIC
g9zd8DyF3s+giZpfUEcKOSRtCr/Fr0EG+Qh6jTqwrQ9Fjo0YIGapSfMnB1hHyCKcjAc9loSOWqoL
8912oGSKjrkm8tvPSWb2jCB4pwEU9SUHwgPoEiTP6BGtdZDpHkg3EG/SsgN513wKA46Mvr6urpwS
zOPHXIRgJMjab9jeswYja5rGklKHEcixMHCIKNKLIjvBKX5cxRwp2mhA3SF9LtUT3JOTkbtLp3NW
AKor5vDUHvSEVjLrPdW7InzvOJMiQhGe/FGDY4J7VJ0smF4cl4hDxIP0JOfB1LgqDEmmcbr6Gy4e
TDKAywUb+GG4MmxRRuLKtAoXOXqzdi/vYYNbQHriPH0TSnD2lwSGh1fuL1OL5jVosU3jZiS46tr5
dfilFguvPjywu89hGKGbXEZE/L3Nhl9TOF5Q5WK9nm0zYsckBueFSgC5foKFYU0o06fbOU9hWNSk
jOphD1ARuIn5O9wz7xSZXUCaFkfiQWj3FnvrUbpWNjuZhrlhFNVnz3vYmWtE6yFlTEBdjQ351Ou9
sJTP8EfGJa4Gr2PZ1fV3MKWqXnAs5exvyjrIruNjlV2iG8kk/gEYabH51+sIbBR0jwKETVHudruJ
2+IDmW53h7k9JLGi9zThTzxuNKoitimVJ8sfm7Cti/7OEXeGnLyL88Vx62qQeLPbNcymJtZ72+Ud
GLOHXg1WfVGORVpkBODLAkkSvHmXOQ/nncXFXZmpQsjmLuDERwlTZTf4Gn3wYq//G/w33Mj10rm5
/Gve25PvZp1vjvyFSTCjomAYXRCmykxzMlNR5Wg7Y8hHOq6XU+JyfZb8UF7M1AooRyZRUoPLtSh7
DsERNXehnCR4W20pbpBfZrlRlupFRom/agcvHyeM7tAfppwQArB6bgRZ3u26x214n9qam08CI51Z
3/Yq7E9p2TrD0ll9+cOkC5A1ZQQb+1k2o0UXbH5GVFsfjzTz4PQ/6oe6Z9226L7LyXWG+oUFLNBV
FS+sq8wyfkiuvTJwgtPD/QimFUlkczRQzj1lGngZtgNW3WUQkSM8c0/wzkYb2kw5hzVxtg52cpNV
arjT3aV8RWDAhW2eSKwO4O9XrcHCXfJyveIQOeKnmA+cgbNFqnX/u5NL3buomW17rwYy4pmYSMG8
UK4c+6vPldjDRGeygS+FOzFIRNDxWqZMxmf8uGNyQWeJXg5CUZsyGhilewYZmzQSshB1FxbG6Bs2
eC0dyADSS8e3A++Qwfi5tEv7Si+cULznPXk2StRtPKq54q6WzzjXcU2FX2IgH8smfVGL/HP5XOcU
PvPaUDK4p6sYDt5OjAR9rnz16bs3lPPmLsgrrFbZp864kHdEVBj6b9BbBIMsNlztu9wdTNulmuQO
KXt+D/qdNoBKwKSIFakMMyTFZ8nqsSlm1/DaXZx4i34B8rRDL2Ua7dIefZ8dQJ3z1tRieyKv7IEx
jdeMvnVJfT2MdujrZjqk3lpIWYktWt6nYac0n+AXv816YakJwduzXJNFgl4f5V1acOlLZVBXmzd2
hXkDCKuDhOdO6AeSWPqMGSwytfQ5wFjSR4lHkfqTCCMLNxvWC1V0GXJYwNEimddh+AJyWCFSbcWd
SduGTDFQ2E5u/HkCLFXmCBbY4AvRVYjv7nFaZX+eVsamrIFze2Yzzh5+hS5OcGlAzs09bBPEw8X0
4ECnPu2sVtD6fntjQubrs8G4u3FrV/CxPAV4owOTGVoqc2TznNIgz2ATIQXnMQUWJD738Rdc2F6T
vqrnZxSxl5JB3FHPb6GDiNlwHTRiWr0ImsVbTXeWarCgG9IiYGgBVyLMl+hESJeZPh4K2O7uY70m
k+tcVjhKmx6RH7uxqVDU4Hle3jGXEPRN9sJ8K4+c+s39dF8xoVc+t5Wu7Ql5JG0xr4YquJbOQBlN
cmno0fXx6PLZVOwDi6J8Tep4WEJ6Bc0m6yfSLMkina3xVI22yxCBTCSijVKg1BsbMEzvGfp/1mgH
gTuX/cHBm0M7cdhQ3CX9kErympHOA7kFbV5/EB8rMtYp7jKjNU63RY1O1WUh5zmRyMYO1HiEG4Y5
odoqayVN67ND8F66/tAexZBiEgk412qaGqWtzXb4QRofUMnJQvzddQ6TMauGDvYVibn4949IfFBr
zZJjWxpsUcVh16Je232SuN8nFCJ6nfrEidT9mShhUmTortF3of65P1+mFxjItgr8M08JxrRHGiUo
S3Jg5OpBZvg/W++q/0AijZ+yo+Hlo0Q2tVanpejVmUaDjx/7LCZToX1VOxvITeiq66tTHJtvvUm0
AzMkaclE9/tGRIZD9MzFZv41/4f4f6XlNHUiZq8CSa/Ei+nAq/n4K6Q7a+hFGkbckPe8Nkq0Lx/A
X5+HP59h5pXzEa+J1jOegy6DHWfTLAthpGRgcH+ojuPTyhYwnUU8Bu5FW2rhUqg7hiP8eSeQZx8+
kNclW1HI39MVgKRIcV81rgdZx4T9vrUmIGhAinqbz2m5GVRuSdAshW6EK17SyatBthS+DOHU98lD
lhOuehyZQ3izvMKhIM2gNh/H1c3F2miZ+ZhB6vuNhtxCoFNGsAE1UdCea0bamuvNXjSn1loA0gvE
h1qZu617GFLWcMcGJtdvrCf/m9iQOYdgXldZl16HgX0nlBPEom/FiPXKkbuK1Ykph+MR5m7fcug+
v+LCD7yGZgqfnYC3CHcSLplkpSVb8BFiiUAZE/vaEF/wfgSsXgeKTlKcyNP9nj9hM3EI9sbHRfyZ
nz8shYpB3atnoxEL7UShxQkWyIKlkMmAprn7ljBZa8Cx4+EEhcJxstrLFRt/T6qiu09J9ysYO5CG
aISCky/hdF3CpJFk4IRp+wHhQtQ7KB2xKrR1XdCDJlkNv8fD2bAkmnHuoj8CgWxx0jX1fBCgTVjK
IUytd6Hey92uSJUcoJuMQzx9ZG3HtX4/Zy763R431RQFYtTOgkVQWDbUjzZXqEIh2g1aeJMG6as6
zXrQkTEBVXX7eqxUiUiNDwQPAN32DzPkSDSEzvcxe4IuRZOOQk8WnIigvF7GxoKHxuVgoH4673Bq
A7rLb1ELlB9KSSTaR4hAL2oO9EID/h3FBWhV3j2IVnfMj8drwZ1zGTk0cX9PmYYPmtzwGBoI63A/
h3pt8ivIdWl7bH5NNyIEM498Eq7fNP9BxnQkMsZIvY1BHo9b/mmTrz6At/zVjZB6UHMjWFklzKSV
YrBNo3tINy/OwXjzZRklNpIvnNOmi2pWuSbZ72whdP7HNVytSAmSoY75+Bjt7867W1DDyTYvlikI
nKSOD+SUJTSd0eiQ6YmvNwvoD2EBS2EcwGGzRI0zJ5QNWj3Q8VxwxTlCPRJhfLqvqPVJRxBn/xv5
z+7HoIvch1/9hsswNjQ8lpM4oGUsAUl7SvVtwrjANyJc94gnYM9+QQgtakOxGj/UFCl1uPJwyQMH
ATORwhrsLZo6qEeFZ1VTeYTLTM4/cQa72RifKgiyo+sZutTR7o4PwYnsGtaXDjHyKFFsuIpe5iTR
ogfd1kGQf6efuqbjmibPL8xFGn7zq5Zf8CLSkBhm+5TD10Eik9pW7bIidRXFBJ7y74WYFBiJmuZP
5cBCd+nGqcIy7wzkBUjuQvQrEgyHVzaEug4tZVN0ynKcSJGVI2tUsrwUuGi7AJGHpzQK6G6qaLO7
QBbyovtr88t8yNypkPO6tybsiYdMk15BjM1LUkun4rWsGZwSncFEKvdVH+aeNgrYo2Ryj+H8W7rM
oMKxDUoVef0u+xOWi71jWAaY+UlxNUvhz3ebP+U3ST7YLi59JCHoHw4Td+2uGq01/W8U0RUt3kYx
vGxz1RYp2zsEBRKYACrN7YlWRF4y7/9KKnBZ6k49VgtbMxuaV2EGgNvP73A8RRTcjRexLdBEr+SQ
8e3+rG3cp6X/7uTG7T0IYL42JJN1Jm3x4H5d88NKhSUknOIQxKjM4GbheKSqekzV5kPccKVY1Vj3
QkJ2wwaRs0PC8ow20IDCSnKVyw9oMxV6ibuAJoGbs8owPNFVXtaTw9nAlwSxXg6xg5MI398YPElU
/cbIL1rQTXFE62CPMBhQ8XzYNJW7TlRQ+lqSYEOgUMA4Tl2fb1OwsnFhZDv3jznHI9VHdKKlnv9v
RN6wDiJoKrslVhqd7CaVS09Gj7pEHPc86MqqFFREqc9GxCpBNex/H7sTwLJvioMYECjUk0osdegW
nDeZOTB+ujv+0xpOXqHztPOEzSyMfGA/C5Pn3iNwW03P9l+fWOTUe93ZHSivPMPlMYL9dqMb+Glk
HR3aNhy8+vhato5nJ1NMqWqktkJozbtBmFHfA0uYT7KGuZmUFfqNdmUhbAKCZFP9SASODDUb1CeE
qL9YqA3osWuBTgmbTiYfUWvrrogzFzXeEnJRLv0djRlq1o2AVTe7HAv5iMIN+Sc9IHq5xcwvlP/8
aqXl1YmCXAYRmKRAj4ZOp0TxxTJs3nhGgHPtImI3kZs//ymG4wcVODs7nPEIQAfzwSDXnn6eGhPc
NDsJUxEmILc+sCXF3QAqFsPMY6w44hQFmoW0uR7bdDCOaL1tExBzOAN9nisw2UpqtqxMD1VuQjMq
cXjXKCD+odSGKZkilzYqq98lnWPpWN+yF9o25fNW42DUg1iz37rx3jUz6dUS4/xmCycyvy7YDM5A
PDGbnHTB1QOzYHTm0C5KeyPcXwEvLnF+B39rfGlwiaO8g+FCyW4eFIKo+tBtNiQVphd6E3Uy3WaZ
FzifprAFHz9rZ+aB1eZcVWvKMGdg/hKMKxgEJrNdsG4xPjTVxemqJIWkDYc/yc/NeCDa/d4xdiGI
s3NyZq4UmklmffyNS/VwqgBbwg+VJkGbLoIzPDXD7NmHcJ71DnKEJUY0B6c+GSgag0iMIeQeYpNb
edkQlvLqfuKBqiwJpq/w9GqHf9pHdJhAh8HBN4NRjBi1RxOofADLSg0o+24G9VW+RqNKIvLI3MWm
bDFQ5mZhqO8D4yAFF1G6FmSb32gqnTl5Axzcot08CKRUSx+wFXjv0w8INi942kZxWAXSxc0DqoKL
JRFI1zdavkxT9TZvuC+AHOcQGCTlRzRPYGam5eNAgggRYvMJP0c9EVBi2BBYO0fkSyx6gnvVvvcI
pwBW/bqZWv9x62isnrJlvBpkoZnFyq6KGEU3jjG634n0IJYickMKfuBZJjKKDnfllW0SrZfCHzZB
qr4kICzKz9fAHhoW8rsjN59ceFa2jsq0U21hJn/pjdAPdU8Bw7+S5KDaM+pKK3yNmXH1AZ+AEJ4Q
sRNdAbp+TjZpSjX1KEdLbDG8jmjOi6dgi0VsQy8dW65YY7Vtq2kI5VoqHTt2+Tbae3syhjvj+BDF
iJu23fuwoT7VtYudIWIEjsDhTBzK2w0nkEw9TnkwzrjKRuQy7S7O1qC7KqhRljNg/fB9TO+m7u1T
Egv7NNrI9ZG9reE4WcMoZURBHxAv9ZelVCwePy8odtjJivBKRLmPlNF3Ip7gPQ3yBJQMKzczeY6M
IKOnUs3e63xI7kt+P+eBbhj4l3aK+z6swq+1G8RoFmf8/eRelXaHijUoO2UODMGSShp1+/u/Fp7p
z6xjBMjoC4eGfI/HFXu0KlNffeSihW5ERKWTOR7RZKFGNqr04GKholHW9P0QclGGakFv0S8Tb6ht
O0roh4dEWnV7kVzCxtm0Y7/HtLRisCTB7uWIpQJTvfKUZXwrICIofLaesKNAhleBQv1eAmslfvVw
kVp+mmGNCYivKW/uoY+6wPdlVJA4lyAhQKrD7doh4DGdp0hu2Wohs77cwyh34nqZCR8tU1SAFocV
AVgR2ChoCAO2fWKj+uTM8JzxG8ptEyVkLH2A8YJAN3lpQX5wYgzKOXsPE5SfTPB6bIkVhZISMvDI
Zrzk2kI5fMreqRj9ZBIeBveSSoYBrdrU2IB8Yy1XtVke7lpcMhQDrvQbJF/xNaMocv2GTxd9r0hp
OSx69mPMlev6iscY96AszwW3+gn9kzwlyWEcyYyc4ALxLxSyKpSkv2UPM+Ddrmmp/YuXpgN7/RqA
4lS/w66fnqlhg48a3J/j4nvqxWQu74eLI0VbJl9PzK8vjCRXSMw3fZEQ14tAfTNDBY+QNvYaiFVe
d7hoBjlxcXtyiqG1ALNaqOxxTTcd7WeTznjDUUYA4c/kDmCQR4crFBrMQdaFUhqsp3FISfNt4WGV
YejQTN2cufeeJ+l/BrmqJFBnCNrlc01gA8r0vLKQlMwthfJkbw4+111NZqmM6596avikCBfI25IO
3uNgQ9ggn0hjdXneRRohDeMM4byADOGhBWaDuiLIdkz6bNmfwue/PgY0dNRgWrZ+qeMVroEeU4mE
L+XNdprb2YWyBDCZBS6eyrTFChbjp01SuqlZv0W9BXx/BHQhVSoqbrTnOodWDM9ZsBvJngZDzfvV
3HaHQHhgvZRFAkiLrsfeMNwiLwcLTdS1JJAbFWnCd/9MDl+roImCp+zdTtdxNu+pFshJM5L3YQd9
gqOfSSWdrfD1McRzkrwjfRRXq3OQ590sPA4NohliypO5Wwmnyoi5v7js1SRBrezvkZMcT7MPjU5j
odJBuZYmoW/Q4Re+L0uXOKc0blU2lewwm9bFsbqzqe5B60BLqH62jxmr9dIA8xxjoc1nyv431YI6
e7pJyRpRXQdpB9ICDx30inmbGfIrD5GtmIBxjrIb3AHh5ChGoJ4a0qjsOvvEO8Z/5+GoX8K1xBoy
qmqsI0VYcyGvtNuiNXWmYlktJeBE207NVDxwrXc7KjOIFvY54bYVtEZgMpJX51MeTsGfmYIG4GAG
k7P5jEPpfdvcXJVuvGpfaHiUTX9i1ViiRv36UrSe1dJuuN6VDMzsCiqK1JIRQyPyanIf9WuXkYTr
t6xVb13lymEX5ybr45RETcJnSNtS0OCKO2J+33qbNufAdKt4cG8m3ouOXxnENlyi088XSSxeEYhG
MHwHAwmd/qwXMWFD29dwPqO7R03fIAeVPVECbycOpY9t5QKbJ3tF9QoA9pHlqL0ZiYEtwpjzuCfN
xHtcYctZOQYDcHuSIHtBFpf7TIVpJH+I71WLXkohWOr7NiMsq1PHcxtD29ZESAUWVV0JfZzIb4r5
L/Q98x4aYG4zWAmT/Br3Gxpa8VDnQRffHw8tmlWALTbGKuw53QSJirVB76AqT/B+sYLj/2sxGjb2
dycR4/QYImhq1Y8oqIXY620iV0XliHXDCeF1jt59Lj2Ivl79CdIu3tfoJ5BS9eD/i6zshmzIMUgr
JuaspS9Q8HPlxWE0PiThuh2V+CsB3J+WHPS70E/VbUF0Mcm0ponp0rRcVk6CkhHjbOQmuvBPlrXR
dWjCtCFphuHMTLmK6upgvNgIe5ctD2apgATqs8X+5NIaxFFu4UIqO243Xq9nr7LVWZpjK3kWHsId
HdJ+k0ABnFz/hZ6wbr5DmIVRzL3YRfHc8HzGnShaPsZUQ3ZU34jfe78XHH+6nnWSf7oMrxJ2Q7XZ
upi7S0iLmg37eS+iwWPtUjhAcZeFzbDUmkx94eHSMF5U3Q3poxIk3jijESKeJaxO/APubNaong95
jENjWF7TM3hrNK3cGyxqR9jSCv7MjKcRzsx/2VsJ9kx+7VkmpMsy9p5tJlCEZ9K4acYQ0phwZJsO
H6RyHRiLX8T4Qx97tDkG8Q9PNK6zURUTsLytILVdiaRGV7fOlcJaomzFxPdbLJZx6o3XndKMlRfG
JQlpJUQeGcH2vHZnErj6K87jyP8OaChU/0UKEpsOk3fIC/vuDTJJYSXurm97KBzAJgJwGV93wVGK
/y7xn1gVl7CnWoNf8ZLR2jn9T1exby50BGN0AoINva2dQjZN5m1Ar3CrEcBb1++v55DKVcAJZ+Kz
XXhBltf07ig5Oxm3pwU8Xbmph8fNMvNIU6pEySPs6Cp0YZMia7XO+cUlbanMTYKFW+EQ+iNZ9MbQ
RuZZT4v+Rf0LnYlp76ChQKNRZ6wgFJmIdodS4O2YuFzUsh1ni7ceROhAl6aqWZ5ryxiIaVOIIv9w
ZJKmw1tcgNHcV5CNkElCoFEUbUGRndOhdlHzXHR2IR9MPMP8w3ECMiScz43wJPuYruoUU7/MfOgw
LPaCz4Gh+C/hwZhxrtKoElg7Wsvl/M+yUzaLXoFj+x8ekoYJsRnoOBdyn04IDPsn7x/Zk92hIDUA
GX1LtPvGcKhNtgcIjJtT+dD8pHqe3/mM5nOa/PMcOHe3A4jiQMTVQzMWEG7v8c6jVlyPHMZR959F
17M1/m//nC0jBN6Wu4tqwcm36Rub1PorORUdbYykiqvBq7yZARTmYrL7VFsYScJXAF4zkpzm5IZo
QSuPrTQDVTs0AryRLS7iQZ/go4elPSi/jr/vJkd2X0pX6r1+930avFeSjgm4lo7FjVUS2o+ff7MH
jKeUQaGKaCS5iItuUumgUtBvCAqfCpU0osW0rO4sbDwk/2jIfVxw38b+40EnkjKqbzvdSRHv9WwK
dp05BWGYa45N+cXE+lvKZtmm9ZJm9X5vg1Xt+2iYDDMESc3oLw05CRJ+y90hIGXX7/WHNMHPeHxr
o1W3rq+kyJZHwXeFm1uOVmzDXQTvsqdI48Q3ediiIZEq7nS4j6GIjUXFLxs5YE3iojy6pW4BTXPX
ISohMqEzga2Lr82Jbv2/NzrHa95speox5C/sOt7cv8moRch3TqjQTdimHOdEZMIjIyGPT7nSfNjp
Xf73ez9q3d0hfchpzfueE3Qf2tWqNjBX2ut9cP26YWkiRQMWpFX+Rl6Pxq/aL/BQxQDQhcfWucLZ
/5p/6O2Hg4SQoGPbzSIn4SBtsyTx+jsa5izqtNkaumnvhyAn7wYVjQufwjVM1jdBSspEG/OzRKn9
UBVr3Uh9Go6kW3yva9+zXy7q6cugCWjNeFbgAkqQZcKX+s5bl3WdSFWqDC4GMfJdCZnH5ZacPJoW
EU6PBaAobN3KB1bCdSecDihRgFH2+E6/A0AgbzEaPCw+XcWJ6arY4/qCg71URer0Vr7yhbtmZN55
Reoi4I1zWgKoGhc0lMhbf0/s205Lt626Cukgnlf6GI4bE1hVD7lODmmRYnmvljo/gRXf7im6q4Fl
Gj8dopWabQUT6lo7dBunNHvi3rE1StL7z3fvtiIJXSLBQL8dzPSE7i4Zw20MCJoKBXZffo6GuOhw
agqzSepcwvPPFZqVyO5BqsUiEESdfydW5Kwczn27eJv17dKuN5kUGbexytYOqYOLHce4fYGyCH7V
X2UBB7NXZl8dS6buPH3Z7YABo3fo+QzEOHAeTFGARZx3w1moBPViMy2n0fWsCm1qmtmHK+W03VhJ
eIy8AkAm8pIch4pMFbmLfaXcQoEDnQ+dRo+FtdPtgbcsemi+q+B6eIXkSIpPnU2qQKdhaCgS0jHc
2cWBjdqnaY0OYP34zUTGlS0oD+a7xkqsZUGO7W9UHqro+lQYGG0MxCujQnX2WGhZ8pJAZ9plaEm7
oL91Qw1IYXHFaVf8ApkeaWBlNKxu+AfCt5ZhfIutDQD4T7/tCRw4RIROumAsGkfRrheyLctb5Rsq
gX9wXpacJQdRZPTC2KKV4KLMiwabUW5AHKP+HsMWAadflyj/psQxgAop0zBmQNcOgbiU8PyJiDiz
KdKlD/u3I6mNy1GrvoBKTIdO2m5EbHj+61vxMQvTbCrBOxuaODIFZFb4jRQPFdHSINuWrp+QfxZu
3sMjxW+llIkwThsHvL1iO6RTBdBrh6ayf1O78eAfQeH/or0CGSinRQBjM2hr7Pkh23PRmoabcMhY
Syl5BsCfKWtyFiAYeDUXOubpe1ybCkNqRwAdHMn7Bb86z1GtuPSJncVMzx4jcVEh99X8trmk2b2s
Fyue5EVHX1qyFtXUztocYigNF0TfjzqeAnhMajg17ckkX6g3uR7v8IMELDCudNVF5DJyIsCJx+qk
AAvSF0RuHfsAsH64YnngpU4BBb4pTTC8A7v8l/2jWHGhs2m+qCHZJE9ZbWxWmNDCjxnWdr/+oFR7
0XNmfijjGSGmXD3PSrSLzspv0M0LubU5FTFD/ML6By/oKGblMmlpNBtyPNfw7g3xgKWme2l2a+r5
CB/HvlQbetkxGig/L0phLBkOAp+Pm2txSxA2K6krL7iaJ99MCITHDSXH37+/lYBgFFjrn3Wdrqad
SEYqMZ5zfxfJhI8ItDsFtfWubzoM6+3bwE9Kc1PD8SVnDmNCjagx5v/xIprIidyhnttiwlmzhbRv
uV+53N9JmQQNnNiHDWaD6U6wpPBb5ZWrxuYRz7rUd3gGjrnL2Oazj68+86Xrm6ltL4g0gMK+5Lmq
Nx3q06Pr479pE9wPkuiGXRmB6l8vPPnq/4WL+r3rIJY7DI8QwELpSoQaSuCkSEbQm661Zx24ey7r
i6t0avLOutBsCAiEcsgadeNTz9/CghUf7irOranFOgDGRBtdbCnlGnF+1xAIW3azIkjxirsEf3d9
biDUkIKT2cFvbKEAOzqii98dbmM/72ZkL36c/xXUmH6vI+mOHM0W9p0Q8c182D8i+9B6TvM1FaTK
StlMsFl6+5pKoYA2bDKjrh8GQJWXtR1WnVCsI0shb9GW3awTg4WYtCeRU9o2cKlQInwJdLXAqi7v
i+j8Jn8Yi6klw2xHy2H7wa9ApFSOjaJuag6v+oruR7g6o5jY30QD/nCXe+zOe/0tlaDKBGMgm8WS
w9j4BanlWFlRHVUEbM9i5y7oj2yyTMTBxZNX4TkScZitB35q7EF1c7C7xMsb0nBsPoGX10mpvVgn
Dt9Ol/6jjcIcdHZiboG1OEHRL7N3nP4LDc2p3/9LBbJnophqe9Qj2ZaShnfqrX2s2lRj2DJ7ViAS
etzUsXCT+VrTFYtPWIHBmWRagA/nzd42DFiBt2tCgCYHq4Qelx1TLEipGxPcokerHl7SozYrFGaj
IunfgOSCqBWUaw4zdc8hiTaBSS9YQxJWtHDJXSlgAAN39+5ZWxql8EHjNuphHgbssnrwKalZKNsX
4NtPTIE1mOA4UEo0Ryb9GaFBbLOc+DxV7r3OtEfeCzLUlTeWa3KEtMuHeHuN3Hc6SFU+xD9yYkTY
bcc8Au4V/8jSD552wSf9ZJo7B9C/NVl7nma6ddHkx+aiQ4Fn6+Rup9qx8ejU6TZGTurawgIShF25
4VvNrMwngjluq326StOb+xy2eVpmXtLBruYFlf/2AJ7wllMXoSN45r6aHxxcVFZN6wY9xvsRjxeT
TXf7Qw29q5q2t6puK8zGx2aM8e5bkrCVdgUA98/RRSX7q/ZPkNUMk+Nd9xrdeVQlMYj1W5eDEXGm
rE1NFXhRApTMlpt2wJ9J3hvwOD1oUcUEfCzvWd5qX0zY/zwEUJ/fhKcMZORb1RJQeRKmH7vADIkc
TJd8yP9AfCS1XjqTl+KADVMiyEMX8L8gPnoUo83aCtOFVbNE1/jCWpceoXJ79bp6EwKgQiOGPLmW
y2ZooK2HOpt0LOf5/9aYH3e3iFEGsPzOT+XUyNDQjM9M3a9OcAVEV9TZOXvNpVEfLv/sF9LaB1LW
UYdzli4a5INqAp4gT5hbNfB2g+P2hbLlECcnG72rKDbGGP/ZAgt4c4R068JxklXz1VowUsOTI4xQ
rICN10YVXc1HAQGNmPYCFNGzfFSZla9Kyl7JIe3oFpNpgFI3J94c4JbXp6/cIHuTXwtlChhpHt2L
rYkGzwOhVwQ0xWRN2JBMjdCvScNw5wlF9UnjFZQXY8beiKLtrSXA4mxyNHerwADRS+TbwWDqHelt
BSrQ1U10q+GsQAT7II6lCsRQqhiDjC0ICZkdqJBoJQnAGUMQZRrH+nLtjUNeeNKn4ONbBSgr3R09
K4WV/HfIXg/UveBa6YXeIdXa5rfAKd15Fn9XryY/psh2syzc78INeZxow7zb6OHYtE7a9udqJZT5
8fVF3E3HVR/3zwLRKmJpp7jOpGZhtjt22V2yKzgf6ksIa2p+PdHvlttrpfA4bzspuRUuJx3qg3rM
VwyiU4XgC+PjjFpKPVN/Sm+MEqfdCebE9MVT+v9wTlKGMwFw5/Qkf7yqNPrBZgqhrKW6L1fjjArj
frqwiNMhM93Yq7vbanG/dTV9STdHHgxyTafmsqVLOMCf9s4smfAEG7GMH5Mn1E9riOxSRztTZyJl
Qc/ONGtr89VPkN1k9rLoOFmoDbNFHAWcXQwWXPjo8q7fhIWDycOH2FXyhQY9VP/IyEWTEhfoS57m
D3xeYDogAtbg1xecp5LVltbloxrYnTu0wCHpCt3+b1JuNYnh7e2nXZwSoZih5/CKW9witTpJt6rD
caDtxtJJ97OGgiQK6FJM5Sk0KF2sfG87kbS1nFPmm7LyYDTdziortFujhUGKj1pQaTlqP+Ugmr0s
zCB45L7es/fhL87/H6NOnNik68W888Fd8gRnC0D8fttdK8SR8EUV0A1Ad+fRBZQWwmj87bPd6Pp3
lQgM6ylKVXfxLBIBpj4XLnHh5btYUJVymSJHbPYZQH3e4ijnev2CxGH37P0Edm023DXgwqkNR740
cwHBo0p/2walrLI3JjtqIH5UTB6VKgbd759RjNtaBT/ER+fhIuc33Bwl4Yg2WbrBKADvHsZju3RG
hkUGBclBki5NVDL1e5m9/CZRKxdRnNS8Sjjjv2NUgUgrz39p8dstyyujYeKHYJz+IL9BjxjA/x8z
km+27e7ofAY9bMRVY52Uh6wS5gvzqtG1kJBmlAWpVLldMMrmRyaV/L4te+d7Q7VfEyJm+gD8tNl5
Vgs4hJv8QQQejFV/o0cIS0u9A4AUjhd+baB77ZdAZM1ju7/LS1cas3v/iI2qEyoRF7K64HQrwIGp
Sv698+e6exUCaHaEMdLP5/N8KgsL/il6j/LtZZ9wSpz+2uOITMFPvlnnoTuZ4edsm402k34HDEA5
5TqX/NE268hI+DHf76dDOnhP8lekdDlYFiLKcBQyzzTO0phjGhqY4KNRLZJioEefnD5mJ36pSWR+
JsxeRuHiwFoZ5WfARBnJf4JcBdCxQlNzaH+JXFZ2z2M8QMwqayFeRwRO5Gs891huPIZr8DDQi8Xj
6UcE+nCCKNMv8IXUkBioccg+NadxiaT0wKQ/sKFEoJPr2GOpkX49akoEtVOr8qQtqg2P2k5JaGEb
YmOw9f8022T/ok/dQ1me0FSX6EdqcX2KL+P7ZBqqhvv5RcaKu6TMqKO4ahqIYwchI8ttAsuFPylH
o14RYShFjjJOqwpetFJhi7vtcHsrQSJbm2J1/C+q8ojcRfVvykTnLog9dBp4tOnuOBuXM+3xydHX
A7Q0qTkWLmSxeZx84RRlO8kZIuOJ9Gn3HpbpRfR0hH41ApgvI0omOPX5lQUfTBs2Kn/a46HwMe+e
tYSSgOmEBqZppnmbuFAVzTaqJUMCwmtng3R0pJEiGFmlN2QDqLz8Obsqlkf6b98LKH6xLJLuRHlr
Um1WwQR0xDh1hZXuT8ZZqeWcCcYQjy5HMhkQEc6zrt5LcZC5q+2uNUCeUVPYI+fKfSQXNofL+R6r
lOFrTb6IhuQdXrDuHgmHD+sdfQvI3yb1IAuoPcgnkFKJsOfE3Ft9swfaksL+vPq6qVhPnv5O4RfB
d01mhYzeVzvANwrIaZT5I8iChbU+JoFjaJDby4MWagbE9/c36Z48WBisCEiQ910+NL3ZnPWiw3qO
yqrsJ15sZ7z5J/VnT1Ooha2lZOzDqZcVhyFtcXZ9dZ09URimqIflaS6oPCPcHWxkR9KyN/xalMKK
XnXrxciROM2zuSuYGBH8EvEG5hRWI7Rr6IgO9FFDlYgLBocz7oGYF9dJ39vkN0bTOnmUR1d7O9EK
7I+ZrmkC+wH2yIIX4AWZ7tfylsrBtMayp+znovhyY6H4jEnI5LCTvinZylbfRHVjn1PU2L/QoMKP
CP+KT1RojyOrqeN6oK2hQbgiY+jl3zcOKV9LMCqI6uitzpPsonUoqYQ86LhPLnMGPEVbAm+PCNpv
bzZVf/T6cI6ju4FOOHoL2hoH0olklCC3v9qaBZvftca6xPKC2NZVkXCnAmstIQqGrypg5+FdyWMg
WkFDy3496ncV6BBv5+erJyDkzKh01GlFpO53A2vl16DVAYYcfD33EY/lOl3pW30SloEjFabvrJKV
gdgx9FgdiZzTqdRKGatRoHxs0YgIKM62Y3lvjmPgjZ3H1Jog/2eWJhYn+SDlHgMpAFr2Y5OLX0N1
242XcI3qm8KfBuz3HtGiVLo3KFziVp4a9YjmlVyEqrBLqe0T4TZye2WLFyYKZMZ63at9VAPrDOu6
8kNgpICAVyIzOVxv0K/ga8L0NuMufMl0LmiZQKbYkBaU6VQpL0xDTjmIyYAbEQf1uN0rf3GxMowQ
IOK3gTw6ZeDQH8H3bkix0DBGo6OHRrlIr3eJeppO+oTDBR62Dg4oDKwwZallQBm/6cZmWWRcfeE2
ChIs/8hkor6vIEdjRGH/SsXpgv/2sXRju/ag4WScoLdhgckodkLyQGkXMvXTMZswlAiMH0sHJSAH
2QdkMaSjOrLB9ZXaFlcKKzxW5iP2kA8oGWVAjHavqQ8O5HcABuccBQHJ5JLer1XZM9Wc8KHhU0uq
l0pmqxk13cvKgLDQ2fG/kVeep3yBTyNScvCVQcREglXr5iBgC5fZ2nJoDSwkGQbaZr43znvs9G7r
DSyZSAtvWlca5cPJelvdr5rFHUFKy8hHDRSJAQ6ejNjinArVYXhCtw3t62IIx9dv++FsT40LpSe2
0PHSvkdjfSJpzG42Ojv5Fucu36rfpuT5S0vASC++LSj4UXbKO05z1GqUkFYj6pqjB/4HEBvuVS2R
yHcnhXwh46Cruq1+fdeA44h57J6jwccquFFmH8iYNczSDB/dQdZvjF+bHr1oigYFM2/Slgl5drsv
/qaKk3GnSs2V3+e1ZqcQO0InTx9SaiJv8SoCQj8r6FgeA4/GaI0wyJptywJw+XI+YRxOXphfxcxA
VF7zP6kEm3VlhAfHfrfvTQ9603nRY1I7RLD/jHh9tevmp1sBZCVRlFBRJS415Xy0dI0eLINv9UKP
OxkjfMX9xJlZXtfnp1egFWAqnFbG5F+5Nj0iEm4iSLSg3yRQC1aa+3sZjG0VVavah+7hRoLnxDQm
7QFeGo2cr2F8RoU9d2zERLd46BS4mf3FfDyPcRA8jduljjYz6hW0bnL7g97ANwr9Kxm2Sm+jIX5M
C/deEw+O0wJx0l2sIDLwU3wGoaI4pptOwM+ST5apjsNUWsX1WpUgkYz19MEXVyjyef+dL57YdEvG
qyBq1vg/aAHpZPIRv327C8HqxaMeYClSj1PTUMTeqobkpkvMxW3TuxByUzvwYEqktjqNURnLGJFG
UrAgyv7WmId9I0cZUyx9CaEPUxWGDhCZOQp0WiVD7XRqMFXBhQHESzu+Z1Yh+JOYzpcvYyUgyOha
E/R53q28ny5RDatEOqNKEFe1usq4IFJISq7cF4D0fb+yB/I4O67Ns1Z+oiZb7fpQasXLHMQnWXWa
l8jd2KrH23MzFBW0/eRAlPgjJ4mj2pLBL2jA8IovGxDGGHyHtskhBUVen7SHF8AXKXG7hD6+ixgI
hMiE9XPCxDUks4E8+6FX4uCJrHD+fwRpIRBmm238JcmPmUPAfs+T5OYjn+kn4CNe8qzgq0weDJdR
pdaJ4NPNCLyAm+zy7WzTnoY79u6V6DheTHRBG9DZGk9vfJURyFw1MoBDMqjSR2m5DCoZNIgZoF6M
yMEDhV0xENEHHlCQuOA2/iax2soQiJWb4tgSX+RJzRdp3hnylnlqsiM1jWv3i1QQhze4iHyd0Hgb
QmgahgirVm7oTRi/FR7MeTgj7XGfT6hLOeO1NUcWGmbkIC+ofaEV0H0Va9qR9ZXcXniQ0HXJgkdY
vwYh75U5IS51EPEeEu+r7nT7YHuPC4WnWrlibUXJ+i//UgHtLwX76RLCzfJZbIKySFFt0MtHV60V
3+6cpMYGqdH55+RSFXqCT9DbPy7dYIySIQQE66R56hqSIxlASfZ1/q2UhHgvIfZqxya7hP0wiNWS
qBTgPIYGjpe0PNn5tbJalqBAsLP1QXLvzclCgajMZTCLDxL3U6/xPZkNjN0HqNoBLXg4mzjjVeyN
m6PzGqXjnKvoXaIdxd1M1ffWd9ZM/Be3/L9qRdt5Vj22LuucywSJ/vPTiO7Ir7ZFq/wyF3rnIJND
d+sENz902CL+wRD1x2JpBosApGBqh1zLEDjlVZ2ExRVpd4o/Ej/N12ydRb92/Q4HDXdVmkIGs0po
3+oZsimgdgwjPvvWZYo5FdTEPUg6kq7w2Q3KwOyzb2d9G2HxwFJsSJyBMX8+1rcXE1NiwBTXCq1X
sOeDlbJTWmymFue4FAELNXFeR0mbB5KY8m3Lc5HPz81zr6AHE5TphRZ4fPo3H/deBpnMvdWQzCi0
RqmsThGpk3CVHLTbiiOmX8E7v7TuhEJ6przOl38WqQ1PTHSDfJADF+UxOG5/qiO144T5XrJgLsAw
V4yZDpmkEHyhoDtA/+ByCdzRS6EOb8p/w5u6SUiOaFLLMn47Fvvm6APHYCKO9gONR4zxu0fJVobY
uanN2XCs8+V5V5F/j/HHBVNc7Ub9lyNfA45TG/hQjnMfv87MUGVJpc/+snqnhHtQJZg7VSKMDHIo
tOiB9yDi+qF7yjJpmcwae5LwJ19Xz+Wd8o3heZ/nkbdNSbDqikPSqIABs6DJZKFbhTz820fqqUaW
dGQ5AXhNsE6beOGGsE8fbnhrovWwXEKz9D5XT51StOeGCb8j3ebcdsmRYgWs873tyJfMZr4VUan8
ex3BkmJ7ceATHAJBsqsxfSVrRcYUH8rSq0l11e0eNJV0kYhZcuDiPWxaZyx8CyLJfvLlPn6QsAEC
PLd01NpCs4cXL69iFfp/wmc1JcG/ARWz7xfjrF1k+7Ies7Z+5VoAZMlkDU5OuEY4AM18+e3z3Anm
W0HaleW3hpp9XcEA+EnQwx54aJLCIHUTIWh9fMLExP+YOJExFBFBGKhmsTWusnvCT95dB6w8GukF
tfqAwdItErZF1gPoTw2DSHtztdExEoPKDAQQjxklg1o13HAgZCwi9W8dhHroboRzsoVm65p8HRvq
vCDgXYax0O2HyV9//c/kbmDZ5I6G5TMjPfg4u/vazKss1AdSrSuy0xF5KTxzkLqmse06A7qbxFvs
F8+gyyZ283BtPM9TlAP+ZYQPYLGrxQZtUNHR8vIhEQrTjUBRTho3A6MGvjuJx2K5sxdTh3QDfswL
WgRnT5YcFJE7zB9ZxLZDfiCiLqGRDN4RNz2149h6Wiq5MgqyHw94JWWNEGuRuGU10VLSuNwTt6/8
0nL66eynOVlxxNYGZJcmUJNY31MBbdgTKjKnyKXOHxATPdGec01vb9Ua5n91/HhMz5SVzT4iseRn
AVk/FvDhiUQrAdBTSzR6lGFbREF5OD0GEZ3Ek6Q8gBLqVJqa6HIDtA2foactTKk8QHrjJT9f7Vjp
AY8LbjzcjdNWM5auLJmF9Gmv8mO8o6I4DtVAovwrRIUPUYcCcXYHxmOsKywfFlBJfpDJpKlcr7F2
ehJSEme1gRC4k7TjI4DsocxAjVAP9Hnc/XsPDU9/EvDxhmsg0f79SHc3P5GjEvAdfBP9OHUr5ZPu
jrv21QLJh+y7OPgoNkbzfJdVP+3lab5iMvjU3rJ63RHvAJpRXpgYbnx53XVVWJcP2o5zN6t3u3zI
CTI/SxYZwP4MSA/AuUkW16BYDgruRZkqzaBJdHUFm8bQu8v0M9cFbthUE+CTGClMgusD4mXhYzUd
/ysYFS74TPonogpm2GZu7HTL+Xqr5WZMUclUF6iwAs7sbshtM5rXOjWIvD8bE1O3aiWO690Z9+ub
9UdCYeFFTs+mh5BzWEonwiGfjYBe4Pt2/cdQ6nvF8RpFfFAQadr11DyZIWW5rjoZh9yFpGAwROxm
Gn8s8t0Vt6a4NWLyZu66Y8PCYwYxmThk6MbM/Blp2R6HY78124i9Mw7velZKrnJKrIgvtC+KQSyv
Z5a0QDxCD+dxKXBPhy0fK369Ud2Bu9Tzbltjx0D14FkIVOhOy2r3VPCwnUkyQAz6O+YTJGCj+vhM
ZygfYZYzR2HSprJ8iAMjmDrfoyXMuv42ZE5po7ujhuJ959QR+uVg5if5qOk/FaRUeq5sOTzznG1f
xSDwRIh4V2IXYDrpNlxcFvGcNruX1slKiT3ta/c8JYyPkd3GG1U7dCUQv/gAPid2v2ZiwDvGDVIu
E9frrLrRWd4Azrf6xmodmPZ5/LHXhet/869S5lCOffVDY1WXbRpCTLhCsMPVuNAbqMNRM3L3Gug+
4XzD5Jl5Dj5H/90+PPVsErjCOqJTfOFjH5RlolduPBouXgDdYQeCu5yQaN0X20Dyl9B7mh8nLMpC
zdBPP1hWqzr9D6H7AfZdbkyirXtbhVFm349Rsnpxr6PxZGDqQgPrC4+aGL8isucEC9xmdYUh0daR
gF5VJSJLCZMssvAs1o2RFdb5f+fYnuAtxUfxO1/AqJNI5ZTNJECDLugad+Jxk0KGvSkZPqFPUApa
ZKzWbJg8LiTCnFeozISMQvHExmaJgSyPhnRLK6355enMVnYQNP1K1BA/2ZpopUEL852dPQK39e7+
eLZLaLWe0eQx63yImFZ5wFWetwW25vKnQaZJOUP/U5/cDsHeu1fYChmbrRQ2NnDvBlMn1hW1YGms
zA8trW/t3pQ+1CHA2n1BmEQVLiMELidYLiREx3RLemXXM885G6zbmv8yNGY0qsdGKw1vQAdzV+dz
UsWg6WLUTmYferzxgybI/BGTm4cijSWS3gnxluCsI+zv/zy5h1GSlr/KQaxvlzL0j9/iYeF3gioB
EZ41bUD2U6i6SI8OU15GpqBLC2LbifEUcy9pUEa3ntFqQYY1OohXADm9QSZ1AV6uQ4btPh9KXGM7
1eWtcrK4a+YJqY32Aa7dbIJTS0FoMa7/D84C7993la36GDCEzDA2C82x8x3kiK9rO6KSOfJwOUSE
azdNCvAcV3oKCmZjUg/x0D50qFv/REzQtzFEV2kXfCupwJJWJ980syv63WvktmrgCXqvwtLs0AJR
qYVBjlR1KQ7sQSpOG7H7kfNr+MOx2eZE+wFgz3sxCWPXNM/+8xWnQ52oxKRYfdPYOIMgxg4o5NQQ
UYCw7O4roXbn3WlWYgsjGQC0GXdByHdrBDqfnsKj1Vt/AKs3E0doFdFbLxj7K8VGIYxsASO2S1Cp
qDo6aeRvFbLUmIJL7aY0QZANmW25Wl1kNGkHOenFyul4us47hMDlBjdkE/evi43+EJjyjFzHwg3Q
QaNTFe5WKhYga5TguJemLRdvM/8xISSycETrsEubmWZ6eOkFb3OswXIS5FmPFKmeLsNGCM4qVoMN
fgBJxSJpsO/eUbVyWx9SOq6aUHIHU5IWFFZ/NUnbf9TfrYSbbjBIVM8i2aw6RRUmDB24g2fN9PrW
fnxJ3loVP8+EO88XDvd2LToKZbjgvVCA9ogfoEZ8HQeC0mojCtxSHYLAK9YE8FzdQL7Gccy5mkYX
nFOGKGVsKkyF2obBjtMu3TCJcn4+Av+8sVV5TCIIlbln3hUFk4NzoRuy8coYwpmCPitZ/bCTSfUa
PZHxJqo32gqgDAi/g8Qw5d4Towb6XiOownbBkT3UCiw/KhU51uvnJu3cZG0F99rNPvG9V8vJGtpi
/g1XOdnx0ObsbtTHm/60LUMIzTNP6L3wZdsQfH/IET52etB6OftLBj4Es5KMxMzP5/7gQWok6mxC
KBvrMxEO8UPVe3FNV3EBueadsvLrJ/oErvrz6zUPgSXh7o8pTYuY3y/5b9UlPEek8y38VIzNhhLp
Jue8c8SE1EyalyRdfzA3hDz/O/jq+MNg4vuyFzEU3KoaF4o/JSvUXEWGOW/hXcJWSOZbebOQ3+D5
n1PxbeiGojwvVGP9hv5YlFpXnTIMmp8vwtj+v7X1VVoDjoN/GOC3+0I7ihEiDtD95DsqRoYCBlus
Mpe+qE4Z3HJqqrs/W+N8sbKQRKM23fTMCVmDPa/D2mBPJHRinvK7YgcNkXLjpDwXW7Ez/3Yo56XK
KcgTWuoRZ/YEvc+AokyGj/nOcpwZKUKcL2S3UCIvGbQSc/n4g3bzApEkdwRT/76dCpmIdomnNvNw
k/+7hSj/xTmbKuehdDbHMk+E4JvyrdGgHFZEy9JSQ+zVlaSiMNCUybcE+OpL1pjeUEYn6KBs1DdG
TSVaxTVZXwCuufGJewLsyMFWrWfaB4EDIZWmPe8nqZglstKnfA9D4xok8k+UZCmPBP6zqTRm4ltJ
qCVwy2crIp9XtjuxiI9oCcCksauBwVCANhLP57QZxFiRtJlISaVgqv9lpY9H8Z90t/7l2X+U/6+a
2d219yGjDNeqnbhM9cZUJu350WQceYsf2s2KOVr1P+c7+dAi6vrJ9FSzhVG+wbcnUZqQYq0YOgp6
OzFNA0+TFuupgx0jBtRiLqMJiWF5oz5QU6V0ukhR2cQBgECHQqvfprlKM2nwm8lhzGwbEWcHrin+
CtEJI8Q+7WKSoqWmsWT+yCg8gxx9SMmqjJGifaUFp1c+HX8T2qbEuEhXx0yiTFnJjXWMXWGJbdVS
Q5IQYir/Vo70LcHhnS2gbZvCn8gCrRV6isxIUm+g30Z9LlbJ9HWKI8vpCXxuHp2J+2lfp1Zyf861
QyDJIUHTvggbaBBGf5VMWyocN/Pc5T4zCaeygVBe4oGe5M33/UFYpOMrQIGWbnRETni4vx4hgm/p
YjAZd3e31upOxFWdtTJKr/0LfwXq18ijeOvHMB5j+1W47sbC1Xxj+LQiMK/BeAq51uHtD4D58sWM
NbwecQicxUXKmN6I6NVqrGXiKX3iuat4IfBE5Ln/uhm99Q47pWePvSsNnDRT2WjXwfSXwtiShIyK
u9HSa7XvFCthaBIcMShOu2swxe5M7ozlSXRfIvfXSKfebhnA0g/rXxlSTKS44Opnjkw3ILZlSRxg
jVa3Bgkcb/UQmxo7hthVRRa2z3yjXdKtaUGRkKEjI2zG/K+/AxXO18BLc8NS4iwc2LVSeB9+7BSh
3+2F7bVFIPn5mWHkyz+PS+p2d8uUngvMAWKet2/+6CIVYsjsYnk/25JILj9ydpjsw3yQEsQ0N3Xx
36fdhtTK6fdh3CDs9mKPiKFJS9zni/HryJlz8zW7EAkSknp1IBvfaEvyP9gwLpLdO2ekDNrPwfXC
nNUmGByg/Wi0gJWbAEGDdJ03xKGPUXbqaLPiNDGmobuQhsG/gGNyHsAWvV+HLn1nr3GkS/9w+SYS
O1kPHCdtxNxQ3UXO+fT8oxPuW4iUsMSGDVRDJymCQpc2oCtVHMw6iXnpNWPmhd4ZZZMt0H30utoq
fhczfP52ZizZOEMzf0X4Xe6y7BJX9R64GmXW6MAfwzCG4IerJsx9IE0yt/MWd7WMbQGrwMJ7uFtQ
IsgZM09GhwaI4td3ev9jE1qB+OFpVILPu1A/SXbF7tSslSVMXGNb2zEgCxxDxf4mXuF6PusBQqie
gyO5PhyCUY/8Q3x8RtiWin8lmW1Rk4yJRhk3juLdb7Fw6sPVPOJLcAlXGxzYyEtyNDyDxEGD/Buf
SvbC7Dn1iLAETEAKnoKeyKBgzKR8S+uhMW5juu6o29D2QCwTodEePWJ+ELqeEyiTCLSBwfd3YDQe
UIdc3J7A5eSJsV1Xpg60F5otze+loYr565MGxfkNL5RF7QixUQqFKLbIwlocwHZJoek5cFqUI8G5
aGHGjCqfwodXif170r5Dd/wb4GBNhsIFaeeweDWDd1XVASkoNBwXxC8l5pzw7SjOxGV7BrK2IbQk
Ejps8VmhNokHU9fk4rOaBKdBgMF/fhfwcMcotT42KAa15WicjOE9ySguBTlqHc12elEm7VqpM5Fu
XWUZ/lz07/PYwDm7PyDOZWdy4CbtFi/YGOvx5RMxmgcsgR1oPnzE6VuK+ybwvFt9369KEZNxBe3/
0sPyd314r1e6RsesjHnGjaBGKPut6JnAP0ScxBf9zzHmc/qGIyDFsejOFizmwbI3ffVtBxBDvkCt
h9NJvaWGFP71VCv5gmfG+BVUjSgFXPO1ZradodSTtdprS5upj0fzVXg5TtfH1win6i+EUDsq6mxt
JXzZc51z2aCfBg8uzZ8kpfu2t1XF68XAPUPK/5vqAXrkKs09+8LgsaiG/iJ+HlSKri+D3+2OxVIa
mgBYidxxCKceS+tDIl+rTuNQByeoXFIw9+FZ4wHTio1dFudFsMtLTw8mbx3VPVvXg6jalDgFr8DD
1s8oeUI1zlX3pouqHhDoBIw7qndJ6vb9q69fGKInzs3Aj35GBQVFN6SLJiPO+L8poTPWL5FHCfKe
XhI3MwQg8WNQ+1s+LMl+QeNY5VyQOnnwbzSZiG+0rKTX2WYsVOGt4fKFFOO0i8SDKi/zeBCIkxUr
AC1Q3/xZsxNGu2uJn72dJCaTW3l3llNpcnrdPB5GRCD946x//WuE/Fs8GV5AUFsKXKtQXYBRL/5W
8hwoHTpyj2yZ1QvdExZ/2L2HNQkts82WfejOZ7VlLEklbjwwIeGCwE4HK8AdeIa1vv55jvOasR9O
SLo/qjen4zfkUFa70EtLHeQdufmrMhWCKl9piYtMXFbxP4t6qN6awj5WSoGuApdSmfP7fhugZRM8
jXrGJVMLBtIsRBbMcr42pX/1QIQArC7ouxrgueyLxVMdZBlXVDrcXG7mCBYnA2uATO7NFwzQ0Knj
7DuGWAc4H7HAg1R4ut9JahITJKeG3jIDqunWSE5ES+kbWqSRCStsqAc7QPClsWBGoNFXr/3zP5To
8ToVQOFv4W8GD+VH+6SRQ5PKlSvLra1i20HMrFPS/HAp3blMzDuVZSL6bigwETD2O5JksQT2X8Fe
LgSI+vbUuCsMjw2DbQ/Cva2j+1JQ512zMou8tm1B5UXDdn2mZyhzy0EtVyEWswbHbKn6W0RvddwT
6c2kO6WLEhlbdU0eo0REqFN8pWvBKFx+JusJ1C60jdvI7+KhtkcRPv/fCAcjB0kYfvMOyRJ4rywt
h0nTy0jnQRzX35ughzGLnSECTjuaTUc8ALb0t9m/ivUXj8O1z2jwQpNfHeoEqbhgIWT3om3lG/hJ
aoAytQIHQJViwIPOrZtH4Kfg5Y7n5ttYA1OfPEKoYYPoC3ZkoXzLyIr+eUgsPAUf1CXZlcypj+rO
8Uh+3ZZZDXlChKOopy2MWBRj8Uy6RxQvU+qyfJVGWUEBILgQVG93fm0RRbxSMuwtjNrAnLt8zB++
ux8a+QpgLXbz9rxQp/rTM6OIvG65v6RkONCPQtJf3kCVQDoFtvQcT4GUnICq1ZKwC4nSC696iQnF
gpPNLo0UuuSY3GPKtk31O9XR77d+jSN+jyIayN6bacvyKyrg//V9lj3wWm2D+nLzARAMY4IN7DH6
+YA6Zih2brn/AwC5NRPI7t4RJ8vO7cdvl96YaMObzooTaPwlsnkV/zUnZA/yQGIbBan+Eqxi0rx+
rv7BHiVUCeFy5GLGIVlsGKu7R/XSIKxhhfTtrbcZmANrwqDZpMhfRh97kPU4PXo8p6GCM/v+GLBu
xxo1hgViHBKYCAoRZ0EJ8Vq9oYN/6Tv2rqDNjQ98iGdO6S8vx8J7kVWC4xGIa23Ganfqhshhrawy
xI0jMdP8fgq12rFyZcNcMhconq94IeJ28k2R42YYNV9rMqCTZ3cWyiqS6buXMmsJ17mQJKimtL49
TfHL2EOdavm/CduwjSfNjAJ4PRHnCdOcsrmlQIAoKixktIOBC6So0XPobIuXZ2M+dHJm23qE+jm/
1JjGkoCV78C3Yx1XmNzzY/heqbYbyHHSUNOjYCQO/GPLpgUARtr2sCr3WKwQ587HLfZX1qzBKgRV
lbDpufQvZQWkaVwpKnbRaGBnZ7kNsNmhguEnfXUKpMNq/Ju7HFP8lfFhihiehredYXyfDZP+Gy1Q
iYr75eFJNO4MdlP2+AZycUOD0GVW8hB49OYKUVnvGU5SlhwoXE/FlcILwBuYgvzI6HXvA5e1j33p
0Lkgs7RzYB+W6YpW5FyZP93tafWDzhFncYoSAeOuq9qY4DkW1aYv0ysJNpXP8ZFucphAmQJLhbXU
0BOIkXVXzFI3NYrCWp/hDepT5WN8ehPv6q4eS1nn2+Mt1XFtEce3wl/cgSE126fSokylKpZlExI0
xXLyAizaJgdOm4a6wUsTgbpWg4gEy3OQhEGs9K2Sg5NFbBrSHpWqfWoKKirhtxQdGjnRXrw6QoQi
myLDQzPRYhrFVDMukKyEpUuOOtsJWSgrL1QExA5zO8v3KCckaPBKqeQlj1VJIXmL7eGFYXiNUM1H
OHSn+O4CiEJfajfmchsHXHgwmDwzJbSWji/tTymhBDX1CK4KqJ10G81/6kSZYqtDsx2kmBvKWRZA
4sKgWSp61yGCfrbFm40sZDRdfVYfmr8Fam9sF+IHqjGW4VhqFGeIrgbiQ+HgYVoPjaduQCYYgmAD
eSKYYdKh4974uUjRyukL5XDILe14jGihQ5qJIHpzWZJWnWEUlDM12P7c33JeNAiF097olEkE0za9
/F2xw2ZhdO6Rav6J4OP0p10Bwo6yp/ZizkFFa+QMLEROgPWupUxuaxiRq1Rc85sJc7NEgVFCjDnu
oGC1MFSaRFNIl739KJlP+PJRSLwuBJpBI3f+aMgvd14+5f2foWTZ5qnTel0FauvU8Gr0xyw3Ino6
XlKD1N78I5fNJS7CCfxXbcohWcLR0jmBQIodZSZgHtB6iB+d/M3AtnENlCdftgID14k8GZyhbVfY
UdM0lvCUei5QSaUGzxJRwyrUEpAKL6/k79kCeQ7g4yfwZ3KEU9erMxZHgiIo6zr+baCKC5pHYnHQ
ezCP7mkhwJ3quZak4UieBYkofi2K+BrQymq7VXEVqli+A0jtsZzlFWINxjc/4iMU1Vx8FI1gdImq
01IiNf8gGbuIrHaJiydz1JDFPByi95yXQ8I+X+FsyXvN1mVSxMtPwfZIrgJrodXE0RFWJLYISVZt
STd0LiZwvw0RDAliJj2mhHt94eqgelBC5kMQJJ3U40UtnOcHoAuE0b9NW7u+py8jso7Fx/ErSG55
PQF4jiqYy+93TPuiPfX+umH+4FmazQ9/OS9lhDcAlzAronBB6ceCHxijiNdY6LoZCuDGkWCyB44O
hNuDEPEj8giUImUlqgjrmHIUZtZ7NThIKXHByNDDR1p60jYzESgB4GdMjFRg96Q9EK/oGhXzhzeH
2wJqTCniqDmQbCfHw4pNPo0+EW0EFZKfyNNVWRe/IRATsevlKmjn/Ei5MOjX/i1DQQsU7DL2MVuR
aKCCgPE0954hlGOUBYvO2/0gO/GrUAjlloc46V6nCPTOdIn/AzGT7BGzU7atYM3vDnaR4wRFW6Dm
17ylWL9BfTTR0Vynnnh4mSaNzka5ow8FYbo28VKktM5xJAQfZL0vpqlJVktPZN0ZBtWLeXfwmaqP
7EUhmtIFH2CKZAovp8SxHDaBptb2NufC4EIgRc4ciqqeZJwy8V/jE7u4IwtPa8wCkozLyRF2NeAe
8i5Hp3ICvHO6fJuLc2DxnOlfMrJ0C2/ZOOQKaROkoYCnhZ8xh26zXhIy5BPzAoOpcrqW5xEPhflD
sOtwxxa56CdCw6cbnK0XKp1vv0I2NAH4RA/hcSjLu/8DsmtDOg8nrcjPwrXaeeRp+Nbf1tjqtZKA
L6qdu2aiyc44T/j+SpVn+9DA11B/QIqXYiYaEkO71UYoTbJyI0T6QiM5ljDMbqvW+67RqTsVkVEg
LGH1wwp3RvbmJ8XIX8zBn4ZRO6VhFinc0+65gnMAbiKMSmZsbzKfqMSj/NoiW5pbMwiekw36VJ+P
Fq/TRSLKVdBUVqBNUR37fLL/pYbx6SaiJaFH6nK6bTv7YkxRaZPzPQMjfXlDXqFIl3ZgmgWrZ47h
Y5SUkt5SYXgNvkIS8ZI9UA4ky2BumtJ0wqy3Z8S6lPjz8Ky+lbHzzVIaidnUxBCgL33WYkqm+uRD
FCL5r1J1mJrMtQe3TLKLbXsd+EQKPfRqZrwroQMc2ZjxjYLEbEQyYU/vsDQebud9SYmdeaR/YTj7
0Zeq5Jed8A+ub99yx23GTD935714NQzO9J9DIZhk+Pbo0fRLvGPaUo769aL10MZj2bQ8KdEamiVb
ZB/aBTaWRKsqyh3AlE8OvZhMeSdohx2fEB40Jr886sT5T9mLd7yRNzu5/5HuynQFsnmNRTzew5Eg
9KtkcaNeHTUFSV+VFOIWKR18uj8rw8AJHQVIsY3RdOvpYiUL1woD/xivU14vvqyNRl7aXC1mYabE
/QfB54y0mLKDuBwiT0swV3ec4QSrFC+L+C3zrMmDy4rPLURtIoqxboZZxqT66okzv9fl9U8rMFLQ
tTXUznL6e5ufU6tziguUPMljivupOOMuKGixif5LbKuvYILqGnqiwUNQ80UOUB4igv/kaLqpcFR8
XXi/hBJCBFxDKhzWn4ChOMi58DeAz9Whzl86ho/jjVhAwrOkB3HFWHm1g7kIGCzCpTczjHd8NJIj
7LGmfAhLconNQe/68txswGHkJ+XeDTVErrptvouw0mYfTPqm+qXJ0W7fOEe9jgVEjRri/KLVwmTh
msGMUqAa42kWHP47VMYkSZgv76T+469XpPfU2XOtCIWQ4oaosXYZdiHDLQW/JHoABFEcfEoH9h5B
e/IOlQ9SHhyf6fp8OZi6vcSxmJwX4e7oJzE3wM+eAg95sUdbyHwSqqwYe3EDCYGQBdBSgZWnS6sB
xrFkCUhL8lnFDRL8dUxVqvWiJ02lJakx6jzJ83J3ngXh/NiDhWOMSLX8Ozf9uXct8G3IRvhzELd5
sxIpni+3MscuZQW2fDCC4NSCpt4+7AdDcQi1iOSdkWJaDhSY00X/pkYFpx40KNXTMv6ANoVDiDa2
Qm2x1TAJx4bp8MnxYXSDfMhZPFVrk5/yGwP/Cp4R/daLTtMtN9iTsNw1zTnU9zzXMgfxUreagpk+
3OJcorQJcgsDzQyDP7Vwp408Sup+7NFtxSZayczHcq4jssnpx21CBj106EQH/ghGB7GPxogFiCA+
YT5PyrR/De4hSvh0vYBjz9AEMf9R3ZowCs5T1KRB3yxUI2Ywp20lms+ESQYLA6JNcr3VRrfcQpgE
PNXjTxUpAt1x77qEpgwdWSlhdKSNONSKnzVIInG3NUWSvmOb5M5Csf8JzYHphE+8PiCUJh+Y4kf7
qlf0VaZiBSRdZRg5XJ6CSiwlNuQszI+RJ/J/sh4rr6YUCGU+YuskF6sMeD7H05LskxlmtUvWjf04
wwbxFMM33qAQMJornHckg+4gcT4pckjdyKhpg5GCC+DM5XXCt26h4u6O0QXxCIyhpLXJ9NhMuMUq
x6uaHYWYpTNYAm6h/sdYbrOWbT0L8dSpizKJnYp522zGrsJUKgAVJhqkc8BaK0uiH4y3JwpoYp2u
q+ioSPJyS8Q4InWIpr0UpN3k/ukKKiSrsDSPZvbjsc4N5sd4MhcQ/ojRcGxKnzY4A0CTQxqjg2rw
LvwIDUUx1Z0wjmqjeMr6dmPsPb8r4nBpSO2q8tDUVB9EWIUjwok/8ow7Lj8u7m1AdVcGOwm6/t1G
CaDMEpYwk281ON8fgI5eHgaz/50yDGLMcPqA531BoiuTK7c3566rHfurt2xUXDR2QKxPoBDT6+qf
qcbCG1tpx0BZOSUr/D1zt15XQfIQWwWD6FeFGOoWN3u+IE8LehDIVArouy6axMgIl2C7wxpJbRbw
t4uFAPVA0G6lsEkNTWO5oJyoOsJfqP+1YklqfZacXtfikv6UCBNjD+5wE3+o9rJv6bvM3SyxRMY0
yBgqC52BlSzN/g6WxKHQWcN3OYfsoz6M2YXAMP1tkZkbp0grNNKWz1cDmrXDg0arp9Br8KE8AW+r
5+3zCys2emVIqvgylMHHFUn6CZbPLi10JqA6ljDh+CHrTo3iiYItLwKDY45FL7RRJOwlk/1Abz6U
I8syxdDDVHdwxWyK54ktemS6oZXiYB3taj0G6iUjOfN7m8uMp38xagK4Q7a7kNGCm1WF69PpAtme
t6Nw01Fvh4D9/8EB2Ob0DQ74juC9HvBqBvPgmEtNQRTAUow7CC5oyEB5JyYkLsQIJZWxvQfog5ct
xSTVM7c9qH2Kc0i8ctT1tCwIYjw2v7KKKA0hEVg0b5XzZqL3vXdYRr1EILX/Ar8N8KX2spv/02YW
sk/uzG7CkHE9yzCo87JWE9gIfl6VaOGqZKqhA1W7t6o2Ig3sY1R/Bo9oM74j1kmDpdf+C27a+Ovy
i7Kau0AP9UiueS5Xl8J0o9qllPijDZXkMK9T9tFhM6JRzZYhl8EZgq+dImMMFR2PZTn0GdHxZxbh
L/W+ldgzs//IQ/C1QLFFVHONUpGwbDOj1J21H6ZI3MItKjr7bKzVDzCOa8BtWR2su0gOxdaXwBjR
EsAxntM0UY+hEkJafMDhH8iPTLkH8yFat+M2UC0r5G0Qi2jEqGzPZ79hH/hY8GJNyFbpYMsWixrK
5GhXQVb7z2ojmzbH9BdIwHXLQdUwHD3Z+iXM6ONgfQsK7l5jCjp7NP5dotX1rHywiZJPddZP0Wvq
OcGK2f19NLAMLIVj6DX8T7prNdWz5G5v0AdiTtF1B+r9zOzKROXSjUXx9RHw6kwoT47wht7VOrY6
v4K+h/vMSVIUde4t9NfR6Hd1dSYPvRvaET7WvjWbaMkGeTv41Dd5auX1KfdDPwfxDyBP9WvsXzy1
GwcDW+7JOlAyevQt2MvNv+ZBjwO7pg4GghnlkjJesz2q3ChHyg2D44Cyx/6l5iOxxqKnKs3vCdLp
KH3QBicFTfb/WWNUPyc8YEspIBpLqj7cQ40rBMVvAA8W4u00oWZGSlL/Oqqt2Ep6b4vczxeMg6n1
vqYCBADZ745c0tzJo2zKipX7P+Gf3NYKVKKbJIWNfywQ16gGvRhyCtLbiE8/z7jrW+aoDxnXOMGv
bQuV6raf+h1HZxRP8GeJxdZvRlTvp4oh6D1vl4DmBgG9/pXfB7rPluvzBU2OPw9vcKqArmrQEt7H
oYvVgJSEtqvifBRCmfVm4CBNTvRSasQ4mNmLxg3LGBc9/HkzPYIZjEJf2qKktPgndzflI3aWYbg1
bG/XmMsA0rzZK/rtQqvbBPLh/TRTAJdisDQU1lXeFfpuUBfX10MaKI50wXKqGnHfO5O82plTnsMH
FmwyOY/XtLIOywL5ZYTu/a4XxJvlnSY+/DyoOqx+rsyaHDF8YCd+sjZFLD2EdfelXAqhIS/tSgDf
lzE2pu8e4AjwuhcjE3ghXRDLBPaKQnP4BUZcz3JReAlU+gc0hieaD6Pe1Dfny2SWGq1ywHa1iqKN
5/zNfWSNWs2Hawobhe76HYMbNZL1rc7NwWMI33AZng4VQIGdK/ehq0RW1xkedZNNBlBwnNIjqpqM
1jnzrC8bnQfhad0+8L8gsGCHk8c/JHLMXcPesbOjEOPfVE+42REJQAGx+8U0ZAjM9hYICqo4i1eK
TE4npza4nK+iTzUcTQmffK095RPbeDLQRvg8EhFHsbtVGrECdtTty00VvRN8XFcZ7vNOUR+t1JYB
2Hlk/Ax0ZdAIF2jaUCqltFhLtovo2G8T6SDjIHNjDiRBUlX2zvequcowB4XNkN3csDn1N9S5yNuD
l5HrAo5q0kQ3SG/73Q+Zp0ZjcBKbrho8xffD78QOwqTaFQAK9bbpg1S3wJTqHCuOlTg+P1ZXtcub
CFmMUeJOR4NGvWpD6oBdsDWJ/345BehzFygismKjTfCrFnfEDxLX9bNYVwvpqr/0sWyq1HoaMdgG
2MVACpLpJN/ssCI3EyeYhmv8HzV59pjJt3vWiF+LJDEpVJCt9ek1qauN0nJ68dXzYEVfB3Uo/2fV
v4KPKsxMxWlYJYw8m0OEZqz6KjrCcgo1zafwr/6W68KrtCoJTCMocimvgs7Op9AnxOS5aVMtVchm
L++WH4mQvg1gohFL4ABuzz09bSn5TMOZMZdgy7n5zSXIPuf4JdgEiXNKB9cnOgRBJBmIgRV7qOO3
UWTph/xwe0vVjyqIxmKwTr62vDjfTRMlKO+4qJl6e1b0Tp2qF/CgN8/Ml9LRsByg3x6rDH/vqeTU
zeoaEtTW3xmQScdmzj/Q/OOiLldCNUE7B7/gJjTJCbup79t/O3u0LHTBaPbGANRt4+VcBNPZHdLF
ouhaMiTryvfAV268KK4FvHVEnwuvt+xb/CsqKBU05l5xRdUujdNeZcZT+FdwvMs/ahVytV4W82Ha
aWfW6MPPNctJ8XUf+jVrr1wzLHCZg7eWIJPwQTh/SV5AALfGUzo2JnZHdpuAnaCkj1R+94e++H+8
xaR4XUaUCP8k01BjfO6RiJSoo/N6AEhMf5o5jDPFQhYykzM2mBLHSBPZCoM7ubuxfN9IIqq0XvR7
2ob4x/CchZ+wgx2WcJF4ISDz2ELPluyC6tJeGt7KzP9DfDLXeER99/GklZZr4e03r67wXhdh6/ew
pD1aayb2/o5+fSOqZpyq+WjCjHXEq+R9CM/dLC9oihrcZ1OCkmmG35zlMBUQ0UW96CiqDJ/Ld+1h
3xeA2tey4EjJgqKfsoqfOMHM0XYeFt2hY8e+fgc7skHwnZsyfWUVz1ZWu75S1J+ZPPWXzx7mlgVE
HFySwNTJEi2a6kCKVwlHYYbBsKHr5xeXPgUfFGYXe0oVEw6dwlP6N+UAToi1QRZl4ZiJeF+34YJY
lgEqqYUSdp2bn0SkZfPMRhwkCsJEPqfhkbOtP04p0ok+FJD5aTHMU5WkRb53eNmWdfldNoZJw5Ku
Iwg1jLTOUznh2r6TrBpOgGzQ9l4yK5qjAaqQuyEweYIwIhU668whNacRwDrXBJ+0sGa4x3Pmt41r
SGo10xvvcIN6LvLmkZwV6Zs4SHeoI6r+/FjP5SsE5HjdpqlzRSskmA+p01NpBP3gEpAvQYJG7zfG
8gzPzkkTXCLIyYFBVvzEiluLsBiWcS4SbA121Y3bWiqk9Z42PMkM4YFJdeEd3fL+tAdHSMVy77Ny
CS2jl8S3xINxi62uNBI9BVVLOQOvURUu08fY06C8WISbLcz1PctFIMHZujOS0vjl+G1SS9jcE/M0
jikUr8qKQkeC+5vJuyBef/01oR5NJKDErn4t5tzT+SKjHcL//zXllzZ9NCjQoqGT6lVFqePDhkIz
1asks1U5o6BjmHqnLcuNyjDHeHtwXQsFMQOvVpgGqesxY9M9d3LVrzsvukaHXApEzMRnWsC4vMNL
Uf8VUzY4ahfrs7ejfO3GQ9W+KzBRgpcQPUGNmUBPytO/aAleXIYR5XiVbppM6yibX757VDX+8bTH
i0Fl5wZreDn1UD9hEV8T7E3XRn87aYeU6DphuAm/ILxMJmgx+oNy6jiG71TJKKpFZrFEG+p8krh1
/dWUlQsU5vqqQ/u6E3dHS/yuYiWRAvWU+Vp9bLddxI6pz+I4rJGXhlWixUcQhvFZIlxtmy4yDI8N
riTLbCNqXkzjz1PS5bhLxDrFsnY9BRIXlt4qPMEwxAtcCxLEoJbDKwGaDfPqFI+g9Xm957BKB5Rd
2iDjBohyIKMSSzhe8MUQKjh1ev+L732/39aeUP1A2UAc25BowwiMzdEs8yJ6NiyH6vAK8YVBaQaM
Bzs76/j0N3xxccpOMqtqVnz9ij+n5FsrjVscS9ZHtHpB6YHsv3IVLq5rYnoiLzQvPDdXG+H8JbdQ
3Z3S2d0IkBf25Vj8FqrILg0jN+gmG4eYS8L1QqLacWTWDgPuHgRnSVe8HpmJxiAyuBD4SQuDOuoG
u0jrHee8eb3ejsfFmPC6zzgzHHEYv2YSW6ya0Xmg0oYpo/fWopsocGanYcHHt1LtKdhOAfSJZ3Ip
HVr2Z3OfRIpeBENsq/ygzsSwqzj2tOzu7YR3fMXRKM+L7ANiPuR04PWKd80cYh+vwcsYKOoUJ4oq
kmdCd0qmEpzZBi3KSotouUKTVGw54hI3Ef9R1TfJTDPFukmjqMW6nc/EwFu9Hismemn1DJDZ/epy
SMvjX+YsghA0+825iJU4aO2nuVyKhNY9WbPiDIGvayThgEMKWSCerCZeJQQtz2Iz0K2qC7jUd503
ufkKNIagoC2Fl1coZQ8202CDrg/3s6JRjesGYsPsZYnBjVere6d/qNXR12m0sR9IqCLJaUO84FOw
pBcDqy5xbvptYsf3cqLu16G/lVx42g02cLU2m5AlbADtG/HuymA4twnPiPX0sZ9guM/nez7CktHr
pC96CZJKrajtXGwXt5c/R6TaxOKBEWJObYtVGLJHvMNiRq334K/l2rJOrfx0mnsOqiOSbeT0JE/H
j28+xnL6J4RZ6TWEU6Sxd0yyLCS/DqDKSMQ6m3u2X8MwbQkbSGDG0Gylsa3LcE8hp24JmDiy+WeZ
J2tuhNNKmFHlvsgNcwujWJLwuFCow/FkEWaBiwk+GdFtON619ikXqGhfIHpaeNMkVzvCfx7uRXe7
enJHGdgoJ6fpjhs/n9hSD+YHvMHFZno2UNE6CYlyrxZUm1CXjOr5VFDcBuO995eqm3ZWW54LLOLh
dXpDaVq3xOHrYPVscLWfJD3AdlPef3+bs8g45/YoE9lxuXaGApht/Z4N+51I1qbcopm05ylxBJyl
9XCYFYqaWGSF4v7J75FanWyCHuH+wOUJ++hx4IRs/f10vYKtSdv8BR42GMPxFvnglQM3VIBFCq2j
J96GytJqR1F9UrkIw992E6cMfLB9GJsI8H8TcCCQEOqTgRy56IXLJR4Nn+FU9tK2NSlxCTzgqC3R
vxIQjPX5MEjc47Y+7z/iGsOjZoC92idLwrFyfm6s1mUX3O3CLMJjDxnHanBGv7FQnKpGxYvdRUSM
LmloHjYS1aj6J18tUY3Lh2d1+7N5HoQfFTTu7DmZznKO69U2QjMGk7fsA/j1t4Xs84PkRqr/Frvj
bZJLGnmeDlnVgm2YdeXYQCDTJ9OAAMolYRnWcn/tFTHIK208TFcpoEM1E6kS5JsW8hJIKF1r/Cuj
8x1hYFBS457wItmJ16KOCg+Wmt/2Ktd+bfCUyF1/5mnTtxLjJonwyrwArttMApR4QEvQAj/4XUzq
f3nVGXNIzxO+3cc/gekrYaP/5Mzs/H1yCwERTgP5k8eho/Q37wpux1gzCWqXQu4CHAcv4a4L9KW1
baOX/wDwieLBUfNI0bFaNdM5wICOqagZAxjirz9uXTRDH77LcF4kW01MbMX/a7t69Oo4Hgod55HE
oKN+2i08y5Ty2T8bMZakGIjSAEq3I6t6THDMH2Owr6b3ltpUIBWxdee00uwpvhpOL0FCHEZZ8D71
V7rFnD0O0YlYz3apCVopNJ4FAnHrZUB0KFvWQfKbuZoe90KD86EkJ2ZHC8EzPBr2IIXLb3Mn6MKE
5e1wsSEwz5q0JLRxwexIgXFB+Rs7o3G8CWBJZ286MqJP8ha65zXYbR0jtXK9iThraGH11nygStJI
rJX2LbTAZfQON8a97vmzl08YaCYGXM2/tA2lliZNT7VdrLoWFt3sfog9+5l6y3qGghBrFedM5Pg1
cRk4k9Ps9ol6j3YKLqnT7+3RK1Q6fuBGuvfGNzphmIP28FspBCiPtDZ8Xn5zD+bvdIViJG9M1k5S
eq+wbNo5/CISkCqHzV8DN0wfqR89/EzFldoC+Ym0/YYX+4CO5G6VClG4Kou6DMy3F4Vaw8MIVwzO
w0I7hcNtFM8ZebACye3QZ7A+1R4+e7adq687bT11WCgZkqW7mfH9OD4LwVTHwp32oKrq39yPUIMV
Sd4UMl0fgw87wV/etjKfoMGU0KTqEeaMUZhLdkGboaIizZD4cEtQJcIhPhuamQh1lkIK/8pG4cPa
U6LBYDgzDem42intjcM1LdzS1UXiHKs9N08YuIhOEHuI2aB7vfhHsBnFK+ry41MLrBUmEZcNM22t
zNnlnZ15g7PELJbpkeqNj3pPfWMDWPxx/9/D/aCuMI6J38Eq2ofETuPy0guoCI3Sh081IUM3P594
mDFD+Dl7JLK38naVoMfoAhrnBeyBTPbWnubE1idgQEZXJBTCXkaQ5PikzlqRFv3QQ/KxaRDdaSJo
QSXWw/SOV+RxkYNE2hqk9a5qrdv150aLnziE1dW8myIli28DUYF0/JokoexksxfNUMDLQI6LcMTo
biiiGGwiwZcjC3PytWHCEQoccnMyXKZDKJjLYHGBUz2Xl/UhIJRdH7ea8+2qR5zs6B//BNIEO317
k54R4n8P6yajABSMhpn17/fzGl7cy6e9UaLK28jJfkxDvQxPEAQY5ALc8xki084/26+JjsL3FNPK
QnDV1K2U3JWDGbYNE5J7Wj8I1Up61N3xwQmNqHDIC0jpZlGiYzfBpRkFvDX2saUbazN22xEW1uSO
6AcgqaBsYC5f3jsKXGBZpYDdbiQBXxEJljCVsJV29fuvTa+MLLyWhMIepbmAg8sCogSMbeg7J3jY
bABTfxW7cUe4dhQJI1bzT3sC58f084/ODCQlfUUFkF2CyyjNOylDW+8j4mu5bwvcEyAFpO5Of79J
e2rkbqfgzvLaKdqwlSxBHFEOm9Zo6BYuYAPoiejMKdl+yJA2z6aljm6HbSOYtUhNVLKo4zrRwgku
HuuXYYP54+rcJJ67Vro4t9PQiwSZGhI9SsLRp5KPebqKXuBuPaL4J1VJMSbUT87H5h8dXBbv4Txy
7KKqV8ud35bKOK/almCMBjci+AJkNGvDLtRIBSqevIfh661HyBR+oEXEOWRW4xwz32V0yrNpSmw2
piCgypIVAS5Z7YBhaGdrMiWuBu8/mhSYVRv7o2KGEPu22l3AAznmeagwqZqDjhSU0+MCGgjS1idp
MjzJY80eT9+bXPAa2/utIe5DYoi/mXMQhPBb7mv9vx/0VqIrDdCXk/Glvm+6FDstwuHq1XsXBIZX
buuuydwKpTSLoJfqr+q0GU+d5LToi7NnMJ9D7EqWF6JnTjMeima3Yz8O6Ihc3fCOXZisFjRq66+1
6HBQlhRy3LC1g2F97+BKXvi7YbbwfqBa71u62axWqOcnO8BOPtinsXGOxVhuOXsErjJjEcQjf1DP
q2UwX8r/Fkj1FixuagmTHEuOKxb7SFpSrhOoTDGDAVoYpkyMTz2X/UT6CNatxjRo6Xju8ZWFMyiF
NHhFtK+K0pEL6oy1Lf3oKKxKev2aWp66IAwpz81w30DYRtKsQOJCp0OhVUGdto0qC9A6bwZVzQPg
gMXaa7CKT5dyJBHCKf7yo/jZ/o26m3i+tK89ld2b9WD/ufCB3Efb2tGZkZyHAYnNgeCPt6SgmNhE
GFccq97QNSJkpVeKUJu/znxEcaP4iSFGRUCeyD90CNtJ57EYGhnlRrg2IwALpp4/h8RsjdRbYTFX
2ThkJNwcEEMl6d7NDI6uDsZrua6DF/28fgcxYMdZUeeN0tNw5/UBzbEAxqiBkSgoN3NPMMUPMJiY
6XBfyDl6qqZ5WPjk8W1CvoQf9pqFrhq41zYePXWZR2e3gchRjZMOw9T1MHwh55XUPIz2/g3igz9P
Koy0vSSOCgrXfz5OKFEiJsfWO5VtzmZaB4kpbkV6DIuTWI4+NOaJPJbjKzQxSu1oeHj9Evvo31eR
mZDNQpZsUCr/wQ04OXfT7PXBHoNNPcF6HlJRtYJPdcJYIugAjjNhVju07oa05uOszv+RPp2mZmn0
JjB6aoATzmjXgxNH+qKVuLzRJNikEc2e36ACHyfc4i2qNVqqs7S3+AoJmcMce+C5Fb9JE3WrXDl0
pmWjUGxuxcTUYzWuR2Qnh9Me6RTIOZ0S+4gjkqd8u48Es3hBSOHs6ry6uzk3KQx03WvLOoNmmqWY
PSpGSwNY9fqKJiq3C34yEFql5NJ4HVB2iQi48wCIrvvggenTM+zv8f+b4Aqg7xi0pcbI7EnZjsI3
pmcRuYjYYpUrU2fjK9jJZG5Jg0hMa5U1f4RMhRlFn17cEo0VbiFQrVkqi/0QVgUN9LXi/Lv29rSG
io8KxxGN0KvokBIAOfXoB2siQbS/358F5P+l3RXOUBToHMkh+guBl9DjYTShX21QaBhU/uUtTnOA
IjmrSpp9ojJ3ayKs4kf9GCBstRKPY65r+Eq18Ah1ghhCBmWeg6MaajL3zqYJc227/iSmfg4oRgbC
vX6L+jwTj0SXbgZHxUrLqaArk+VV2F6Qlq0sKJsuIzoLnlo3pkebzlRBcgKNO1Pna5O4i3dLE3Dn
EyJJfLMN909xxZ9QmeG6uRpRz3wN95UC73AJxQzcpj7ldjjHlXjsXewGOT/Slnk3VgdPf+wrCIM3
lums3g4W5wDdMzSWcZANWtPATUYUFgBSdMkD6z06iQrOZC4roowTtiFTuTorFc2Lkq2EX1Y7kFnb
AIT/wuFvxfZ6Buayt6wGxYpoCsmIAWg7OaPAxQONMiKo1dikCVA7JIj7RCQDm6nphAXhJGu/Tc8B
T17uQyLXwyObiZx9BBmYwb4mWDld3V0BrSRJOq9amlT6p5Y0mguiQV00A1N8Rg9i+sMhrkOJ99tG
Q2xvI6zFEJUaq2OjNkAedvoI55NUvXA8sIzk5fYVMFRrDipPy8YN9S2XyrOnY8LTLYrcNdsOoe3F
I4wOgvZAlfixn8zDR3G4N9Cp56krs60wMBSD+TnDGvVw55q0Dlrnp9bLg53FU21NQklmV7CCllIQ
NHqOSY2+CG9JrKuzRzgonoWFyJFB2F2ROzZD/6miGb4bFbLjmjr900YVArBXrscw95gJ+DH+atRs
tkeRksndDL8bM6+o8XImFXDg5lKfpHnBH1rhcgwZsTt7mmuHG2lhET+qt6BakwxQR8m28yAwC+Cy
GVp1GB0z/m8sW1AO1nzD6qd+Q8N6wNR1TfhVqYLoe5iL1UrGEv0xdTfso1atavT4yzxzxPvBBbdL
PDkh2thjZNHRngKUYsE8S+sN6RnaozQpeAMPg7I2Cbc78xTOoAO66Kh1vqZNLxI2PotLEHzz1waC
iYUV49ARorgU9qL2AtJJY55SJIdMgoc/B0uhhVJ30QKUIyzS/6svnK89Fbsvzh6i6v5zYhKCzGHi
vqtwWDdBEGnbzh7JxJXyX97mZO6airidXwOtq1JwDOnidJlNWkB3BXJW3mLgFZKa/Ul8hyCRUwsN
eBEKwY/u53YFAi+N5J+q0fHd9Z4Yk5Tz0iBNnsoWWTpBraFXNOSWh17lT8CuoScWcFl/Lp4KnXLg
7IFjVBByuDRd1XgZFs7sszY0VuLd31QtEmqZrITBNQfog9LM3O0F8NILJi3MfGOLgm45fPSCAtK7
uhkuQoZodZ2sm9zhaBwV1vaFr3yalUED4JTsEAwQ20vdI10yi4lBix4khFn/Pz1XQjco/4np3L8o
XePjnThDiLiG+5csyNKTtWBr5p7exbgK8Ocx/PUAAy1tFBQHOKVBsvcsHUUJW2cEdmV7cpHgog54
0e04/ZyIuejC+f4lzphaHvKP5+Z7D/j84a2D9oDhPlsHmsY2ijM02XkRzebC9wtibBy+NgUJJ/+i
u4VeTyKNdORa/NgoRyf3aOrDzq+mN2xrqUkKFZKHcPIFFTSVfYYCdKfduWYs/fG+WO9pnpFTrzCB
2SSCYDXudo06kQIT6xOocr7dLlxdM///lwKRverU8bExzhqbBdflavqik61slXN8qNQSzXNpe/+k
yZlVbtJlkigGb7Q43ZVBFJRkdK0yzDY9gzFY3gn+jpgye3ou39kLv7siUxQbcLcF206mqYNZxrNa
dKHPKgulUWThAVQs1PbGk8REy4QJljvramz6dCWCFuPLwIMtvMALrz2klnEy9pqb5IPy0/zV5RmX
OUHw2DSveYF+XAD7pia4tX1Si4+8klwQZJaLsf33h694RwUYKrf/oZOH49mpvYgH9zpLaLp8Piwi
nAz+uLm4s3IhfPbhhOBLUyxXJjOtFnHDOtZGXNoZ4+PpV/3pLcvWVjM6imrjNHHvFBcxMQssAZCN
5F7YcKWq6DWAKc4ZWy3NoZz9ibEP74j90/yWkq2hsQ9WFri+rFA/m4yyVV3cog7CLzg/xkRQLA9c
oJqWwtMar02Vo6aMmo7Ij+LGpVMfbYquxc7APUC2G6SMai7N3I+vyRlALeK/JCVlpR2Ef3mAY/pW
+JAMLauoKePVuUycYRLfMIrUba/mYHk/Ewty2z26z1IcBBIdQn9XaDQMGC4Ccs5mawVtRjPUvxbd
5/fwG3JUgplFQS+RYjNg6EkEm1mtJxc8yc+VOmDg50HJdbL79/Fc7Rt2ko88gvEYQ8o38B627zys
BzKCQNZ1Pnqf6R6FYoAO+76tjA8A9SY6D4n9KQ94iVsIhQzTAzoAgU/J6OB5VYNpHKKDF4HMZ3rd
esavrcdkCPgfoLd3X/mKWzIAlJ06B0+vUJDRv9WYsTLOY8X22G8/1X4QHlygHHXVOcETdG3pooK6
K57FGnQUc75Zyhm32B2mJPCNO+yW5BVjpCOgqA5BN3V5xP+RSF0QXnUPnGt0F3DxY95NahOGREzi
IqJTzqsB8KVdMmb3WyAMeU9jDlLGSffDzLjLUoB/hi0emSQ6DD3piV8UUs8sutNmhS8+5HMupr4R
co60m2yBM/FMTGnVvGvN8xGWTtmp7NN1i9B+eqfbxRN+sxNrr4NAfaZmst3QDwjy/FT9PIbMzWid
ByT+QddIq9RypEn43NgXyYUT6OLynqmwKknxiRauT8B3ZIkZevCNYhRepULOE32ipiMNpIKJNDc4
DjXADNKKlblY75b30VbMIjed80fC/ZpHQGviAZ0vZrxORh2zvU+mcUVjwSeoopJ3aArFnkGjM0qg
3z8MSVNGfEpQG4EssRD/tMWDPzW2wMw1waxLusU7MoPHlMxJm7uGcQ66zhUmA24uMj0lHQaFCDnR
kSx3hzPqcY11el+clR9T/ydbZPumN8LS/VI4vfS5kODidsZaRU5iIuY4GqXDiqfB0v5VYsZDIoiY
uF5LWv61wHV9FStNytLY/+rw5BZVPk6e2FYZqZ0xU9rXXI2VeIbWOjwjZsRpYRSHDDYPAHWj1+1j
Is+ZwwAnFpp7zrZvhJbLdW7IidJwNdkQzFB0bFifqRFTYBATeAbzqafOlneseVHVDLhIg9Dqn1bI
jH48cjTbqScJsF79H3Idc+SYR06KTzKomf3oKNBeSNkHEzf5q59IVwgE+SnCzHVrfAXqf9gyggfm
/QSq+x557x+fGiVFUDX9zkb/4TruL/I+7rJevlOwbtifEDKLrtseW7kCSbiI3hoL8MqWBZS3GNlV
pLymZAt+g+MYg2zqGP28mVpT7ipNDAP2IwY66OCvsswttl8ohtJFmXNtUM2z8Nroq/ExTK7fhHT8
5VJ3inliErrqBbsZQD+Dq7L3/McIymEVcxic2ajP/WvBojVYdAKThYIR+KDfgKIb7eNXLiuoNgwg
Z2ZldzF7qvNBkErO3NkjZ44jgvDsxbTEgPO8cmKIYisPSa0jR8yRexPYt9ctTltLwbNjGLPinQy/
bzwznc9jz55jddgLcBxmJcV3U02q5H3Syg5BhWZR4uz1VgRu9bIG+7ZymmgzwNuku0V1cmmgN9xz
wKkOLOqceiV1k8TvjE3Jy/xeTVLPk3WpI5M9U/ixJfPAD/W+Bs/IxvnrJqU/W5XCz/RRR2x8MyIP
uk3Yf8Ahds+xBLsUXoDW5afzg7+s3FAOkIFs4C8HMqSuu7QGniTLh/MNVABj27F5tv7ACqPQOrD/
UKgv6XksXCNOkYVSb9tRe+xgJZE1DFY0MA+cd9EUSnuHN4AWSlJY7RgHGR0QDu8QrHgZH6CPkQmL
Skns8/ULhIKgs8qpjBknLzQoPmYAURUQuDiH4VFs9HvBGmG9kghUidl7qPSSndYulNv+ojP40aGr
ravHDLCwuNWEkaYo7+NP1YMAiYBwmRZ/zq0aTvSaKDCSSIsTugSL2AH3CFEz++1MsGhYTKpgC+zc
ngwYvEY3ntlJhpJVRi2WEwsjTYtVDTL8lylXIkd+uQZKPtr3vXLhD0QmxoTAENxpOXFtRhnVxXFh
aRGDYoJ1D8az4D5eAadykXz+dIwtwVohBSTZHokffJN9pHT4a6rTv6efy881NwwhcQ0sTN+UD/WQ
DoIhXKD54FU8SIQ5/sVmBqPzpWYpEoH4Q/e4qUgRDzdGdB0DOIu4y7RyVs2iC8gAM4xsVi4xS/QJ
K9D3vSIsjmoxGCEbssbKPYJXte7eV8ljS1HJiukseKRKFge23+/hKjnDMhTa6b778zBsb1r148si
cXKrApHrtRsWHv+wLUwu92/YOAGtIvEjBYBNJw7mKSVrecKhS9OSQ/3s+YplHpVjMFIUC23/fc2X
a418W5ZTqJczdxrRMpypHP2/hz3kxlwG+amsLoJGvIRJqadrmsQFfYVHHdMiEmOJiX3GZtZYQxWR
yadOlLiVUWOYBO74th/7uXlc7IX6kps0POz2TTkBuq+gT976SOyenfNrR7qnXSuD3QEGly/776+M
TMMucNnvXAHYzjzfsqob+K1rbYaWTvUTBRJkTQTMsD4g/qx8J0/2+u3FRVY5ccqHzBPfVWUIYfTb
Z+k+xtw4Q4O9TJcld2K0mkpK9Bsth5b8gJYd1ieneARCwug+OlOrZn6geGRKwOcrSc1oUr5Cvibw
dHEhnpA0PwXKa6Egul8fuzNsbjA4nonCOvPi6VL0stmb6JL0tuVuURjOXdnUA2mpmgCL6vmjRt4X
WRuO8bD/Y7ZAaJWKecScrUNw13W7S3fEnwtqb3B5/AWHvGbxJcB6CXkGeDRxF1Cg6TtCK1VMKD7k
xsKemGsLACHu9VWyLb17XAGwm9AzthFARmrxGp+Dgmw/O4EzOjym2KGO7hVl67Hj5qgFDMk2qPLg
nPnsG0UV/yY8t311EyfFr3kG64LYjzEcRXhgnw+ABpw5t92ddHtLgpdOBOxphxbg4p3nI9BVxeDI
daSPRat9VaGedAXX3zbh/crj/DwHzz/3FLHgPHKmQ/JSEbPTtgs+jU+JW9c+sNQbuoR3PYPSlALJ
7BHfLj0+wtK07ILUTwzLmk2vt4pKI/CCNK1+6W37hjzwQtemi79IpBt96FZaocj62bHnlcG+QH5a
+E3rREqCivMZ+isCPS0JNnO3mwIDsAMvBtTBEAK02Yaw0SMVLwxMn1ZuXM/1d8/llVTU6PJlEkOa
nhUjPiAYIeb39A7+851SFlFsrvHbk2Z0xDwxu/QUzZi3LxhSPauCHU0A7mBIK0IC1FaWuG9U3sr/
8gG3wjyVGdOfZ5rt8+itCfJioNCBf6/qSI8zpTtTFLWWyVbFF5h1HS+wEG/azXu/wSA6IFgiF46c
+A9QkeRg4zEw7ckneORGJEOdwczescW8FG30foeEnVHaH6sWBRO08zesCnRPN407hjpBuY+9UpaA
xapLhoOYpPrvCt4jPo/NDMBkp/lCM3+B4fSf8KsMjRvVyMbx54wsMH3BDq7myyGvzKZje0F021ls
r2kjdhl7GZFOpiUW+g+bKjdGBCnxtnksn2zEmP0gDn42eiKlT3N3hqQzY+A97duyQRU44x4T9SyI
3AWthGK/+MrlO4K2PWvLqe+xjv1mssYVqaMA0kHXjSTXHCNq+CGQPzSip0sRVRVk8pssGp4XQA1u
swSKwBdfNHk/hxRWFvdExH+L03sS7frEliR7CQ3o0Dt4J2XC1pPy1Vm0zWVTGlf0e0Tbavpq0c9i
atY5mi22UqZd6DJ39k/K5UhYwAY/0GAoAEw+vzE09eeCp+wTJsPquF88/41aarDGcdfi5NcG2iTH
ojWZmeZSW6Fu3KnvoNfi/X+kIFzBxkv0wRAJzMWLfiEWDion93Q73moddoGoH5AWWPxVJB0ux0hq
YmZ6G7wNAlvLLtIAvO+qqVieXJC9isFvuwQoWoD0riHojlQoWj3h5If7DgwsfVtTXGjMIoUHkswE
i5nPDqvJEK4qzu5mod0di9FVIFqX6VhMG+Wvn0hVVQGZgFNTyI4egJ5UdYf84jgetJ/bLhLgqUZz
/4sskIHyV+Kb2vhzg+fE/EmskzgbuQDkAh5++y2LKJSfvCqZYUSsIZghn9r0oRw1M9Nt/4Sua+SE
Aji4oG/TEetR9uKHStI59/YlsUubsO8hmEUJvZxk8A8WrQ0wmsnCO/cpXdjDWOFPzF5HkGKySSht
+QFLI9ZONRmtHnj5TQIhChXs5iOpTQHZyZdTvlSBeYrEel9ZiW+J+aBcKWGdkdF2iktmffEmE2FT
WMB+Nq3QTnKHPBl30dFNU7x8d3E7XLcW521R2tBopuoOkMTQPM1/5L0uV/BALPQ6DJnV89YYJNrf
obxUDX/yrsyZNtbLhB6YLa3UQi/xyTCFE/KXHBzNl0dgVViqLcIytlXsXRrO7vOkQootlchHl08u
2uOPzYa59KugQSe/76HnoxkW29zct1RL3TpeEKNIy2pdmfCmBVQ9g8EyYrhZSu7rF+ZLS5QYyaBE
lV9g1bANsV5VyN0i0Hfy2j3eb2iZxVUdArAiAQT2T71XkbF6fVPisnT/ruAwaySiMVR9+IlzhS2J
jnJsQSmCGPonZvVevkXhS7HdBVH905K7WX6n26fFOWlhbsC+R/yWwy/EPxbePQgzs9mad0irMpa2
T4ltWSeDFmE5kqiEQWLR/imxRdZ3cfqa+AoT7wGMdudngAgnFlXtxQTcLJfh6e9hON4eGv4ZZE84
JQC2lRozh52wc1cqlwgq7Cm0sP/Wyji/OscpMo68S0qPR6MoQqEkKIwopsJfrWgrL61wCc33sUaY
68Fy3+kMfiUWII93aIP8efdRm5gTa0nHHse23cnbW500ocdQNncUNbSTy6mgBzhUJvzfdXgUoyR3
61ydS1Wmtv8xtXShfhu97GEx9QeNW+a1WAHJgT061Fdag9OT2N0ODFy7Saj/eWe/Ecq7kcKiop30
VENmVFjAJ0k5D5ku0MKUSj3Xt89cUdZqiM1u4YS6IP/2raULWAXI/i1Ohdv7Fm7dr1TobQ9h/Ki8
zoSzRkgVw32IZX6u16rthy1oLvkFFuFp6RAsTg0iDOHFd69pV6d13Xk5cBoqwXoHqDsrykmjHLDJ
iKIARHQJFOVXhQ14/9beqJK8rSoz+rLUr4UROnDxnRROUJOPIdpMKBMiJ7ef16jX33Vb1l+xqCm6
kNEaIq+b54ECXi9hqSjCiImoWUSCUZDidMExuWCPyggBs530RsDGBk+YinUYbwMyZR/C9+mht9iz
4UUd2nv8ADg/VK46K0BrsFxmTkkdX5/C71bWOMLRhTLRuSRGgLU/6BXoTHiVD10v0zvsUaqWrDwm
a8YqGcG6aG+BDXehAsrndTIjyvGwJwifZvc6W8CZl35rvEQPFq/4Ej2GNH/H2xWwZxMDoskVyPE/
oiIeB2vWQ6Hs9QK357QiWoZNpzgvI/UpTO+6V1t/3AYwqffBWGJxgDNieZ/83DvSPaPy6my6Vhvm
oYC9/NsmelTfE6QRUUk1aeI7SM6KD+OFODQOqQgmAT8q5vtgsYUwy7F287UQkH0Rx18OzFmMAm/j
UJUq+91sj3RV542wbpi9eD2XQZC3WaStNzX7cJZGlC5zLniFRKGzxBiz3HlS18+On1yqSeKnn6yj
UB2wTtSoA4tus92+NMu/Iusshxrq2k3bZW+1txHDNHQ33t6d9Y+pl144Z+JyzBxNOcF97eXTux/t
gZ05RYQydZEg1sDGsSMP4/tnkD9hJ/BFJAzD/NKUn7pqpxzMFPgNxAkHdk69XavAt0KsFtxMDVO+
yAx0EAnh92uhSyyM7wsNzTg9XMBUKqFcXcsmgFNFxZWnIYJlutZ7Xw2g1rivuvQBwz7YXDd8cldc
kL3batL8mT/3Ly/ng4XRnEq5A7cl/RW29N17nx8azN+cZdskYdTP2FzDAGbDKWzfhw3IcpBtEppI
uKG/3EtVUiz3ZD5IZbgkuouDfVF/rN2rE/X/cxAcqbhngXD0nybB862UhMozG7zj80vLYbnui6dA
krZW3xj2lVqb7NCDI7YFLl/Czxms8aAkhUJPQmeu9Nj4PnWHP+6ddfMTuDHwEGqbN/vF8OqE60mA
RXsiF9mReH6DrBahcnF6JMQgQKhRef7DpXjqxs3DUI2i1zdIHQj3vLO3idnBIMKqVwo/704S+oHn
udcMu4NyZJ5V8W+30jenBKLjo6G4VUN8h3DqFTGP/0sQVa2xLNxynD6s0TsaCCUk1F0pu3SmKd9E
3rJzkcDnUf+ZOJztmp0n0jnu87GDpl2GvsxuMngqatanbqe2J9Qm1nIS8heMVN+Hkdvz4lGqoYzY
N1rW1p2yAkSjR5eOaea+9yvM4XzkE9StihNSUmDoc0nkjXkIoYtRVjVVlaw9lY8pbEJMwZcrDcaO
Y61C6TLMbeEdysaFgxKC5ugDCSjds7KELT/DdLYOUXvORFvgujVNxvjjXGHqmhfrBGBAAn/ouL/O
/MIq5gdnDso7GeheM1mb8au5Ss8ewTjssSZICkQxe83N5EyvL6J2E67r/8UQNIY5H5M7E7633MuY
Dt6FuhLk/ZNmIYHrwSTZXB33SU0eEp6Z/iIV7UJA0qqmncYGmHvVzlZ1Aw3lKg91rQohKIANk9IR
jNkxcaNKXYYgTKr1sA4m5FYeljss1sPyJXQVcIGSpQaHxPIcRN3Q0a7RJwpmd8QD4hPGBpacuGcZ
X9py2LdcatuwLXxGz6g6Y5FMS++6u818KHDFD4byjq3qnY331jZqCRh0aEwa+G+K0rcyFFVBKjP9
lYmRSNJOc+UMO9xN9ehY4H9AWAdnl878HQbkiwtgq32IJDghsAkCU/4VpwIxU8K6Nm9kPKmpLgAK
wHEoU01qyg9G9WAzNLXaTzm6KeMi0l5jZ0Fn1+d40DeoskoCStGCeolU/9U4q3wcxKDQV9lcr6XG
J4jYvGGysRelcB5IJbdFPChmazyB1cwvYVbPEE8Z3dLbAzQLsaV7AZQMsMywmdYeV89Fc14LlCXl
McYZ9esRdKoRunF+7hufC40zka76NuOcJGQeqAGSU22UZKKaPXy5mhqyVeamB1hF/j49S3HCXvZ9
XGlSCcqRW+VICG8er/F+ESoWeH3aekF6MaaV5qAgmXahg8DUkWp1hA6gfJh7hQE4UyX8luicHiS3
Opb8v58n36UnRJ2AUDmkj/A0O8kLuxBTweJ8JLUhszidJnedule4xayugLs4dCqSkba3hYWBcgk+
ei6Asmy5Cq4BESYWria/SLcFIygtfTYg+/bQZ6FHsom2O271XowJAiKXAkSEeGilCbvS/7Pwnco7
s2pFiwK4Ecc9HiiOZT9wCgeIJ4y78KZXquFiIQmaCAu1D6G5ZOYqdtRb2ChNvDEcMlXv7epkL7Q5
grxdkXSfBy1fuE2n50zrpZK+B9zU5e8fvDo4wvUBB6tGblwrpu3n9eG+TFBGJYVCZUQqJRQ+RSiK
r8Yp46VEr6aSkalGFRqdbBzRWaHru0VwOfjpmxwYglsgQ/wDVWHNLQ6eT0SY+eQ/LfLaW9LUud3t
F4S5W+x204TlRvfCgw7LBSJmCiY/PSw0VKyIHxzD5ZjQGT6M1QMSUWuKVqAPJypXI+qSdstwevLA
RCALNkw8/ZWvMxS+3P2d2mruvVjS/Nu2RuUCGXD9KAB3Yu9Ibh3kR4FCMilrpi/ofW5oyRYsVo7O
c70d3iBcXUHOxA7vqYPl2aY8+iDG8O5nz3w2cAti49ASSbURQ7d/2qK3VctILsnOkYvADsFqd1lN
vIfdInEJ1bHEF/ehjds74wo8/LoYgCrdcc925D0sHHj0g5eKVDGFvQwGOsXalPjypS5Ymw1mXVWH
Pyi1t3LgRwsxUimEHQrWVyy7eF2yzjwhiKqIB4qwHpmlWuOOeV4IieYTCXGyd8k4eINUXFuTMe3c
kv51nN1ALmAUPxWS77MFYadLy/jlFHxJPJtJk+nAun6MtvN4vPOnAn323PDfvdo+iQqltfRveSgO
UzP0jbsTVGNh8HKxiedNusc7bX4jx4HWAyhN8AlK1yLgDeBiMpwLquQbp3bRt8jkmLIgUu2p38fE
xZFgu0A+1jTLNKRuBvONoDbox69sN/Zj5JkG3Q33idGYHjBaVybea6Hoc7GshO7pG0JbrrNmCTfE
kpRhar8+zIwybtbk8ip9vVQLXyMF7JLcQSkU9ak3w7YvlTv7YnxYJsJyqMjn5cTJA9hPV9JCmy0d
g9E6aqJdvkwXkvfJyxPokd+p+XQlbbkT0PzBId6D7/+rKLf67B6LrHx+KsdnMwbyNXuLMube/Ahs
pllp/vXIpu/qxFW82LS1sKvC0nXK1o8l01Px9tMwq1fh+VElO7yiRzbLlJan4er15NJwwOzeFtsY
Q62me6LYPYGRoY8I3YlYXDJUvM929H6RESau2KzqAtY0q/ErcEZDfSUYQAyrVztnlFVrgtHNd5V7
C4J1yooGGKHUx1+/uP90Yx/Ym60z0a1mswseXg8bnKON751pbyd9oYr6OeIox7ieCDchgbciWZXU
fs+1wh7d0qedTRN2nRP3vbRzfG+djKW7ysh2Pt8jfUHnskRk1Tzma9eSfLVEFd1/soYv0/+0xvRL
B/yEXtLoWf5zAUq0TxY158dJgHLkeaVte5AmraQWaote9yiWEUyePiFA17HqkhuT4n6FMxjNPirZ
U21Xzedf/InclG9jCrOpt6OXZmwbjkQpIpPYA3EBUYUwe1yYf2rfLoq3GIE/uCS+A+TT9km3O8V7
78DouzaQpn/jzvaHYn7tepRyP/ZnBHQrhCeNbGGiSOUGmc8ppGy3HF1rgTAsDCtLYPE7Mva6O8TN
CDg7VhKUjx/EGTrMnU7Z8MxfOHh10+Box9XJf75EO2py8TzdiBeuZGU2bs67EHupyk17mWtOf08q
tVgbn1sTekn1s+atASqZPOQoVJcBA8cX5NrXT0mfI/WrIKF9gy+Djf+0LWgoFpdWTcG58V/es6nG
+yQwLgNSLvB1Df8b1OCE3aXQLRWcJWNUu3fTxa+UnDCyQSdTRTlglUPcfF6ZbWWoGkcMmnJ6QtaM
4lUyex7V9i0kwGWKbbi4J4YvwOl4oG0XEynM4LEOjKVoqPmsjl9hWgLKHGZQRE25AC3ZVt7d2mQz
TsIgShmosuGAmGGjgDhVwxSgkKEIPZ/rbxHSkILFZqzY96sBM2ZgH/j7hiwVPlvTCo6/4pMUshyN
PRetd9wXZ2fg+WvvCR+IPdtFNdNOVzXYSkGDEjBonZNDJzgYZx6paXXlWvkktM0W6blLCigK3Sj4
o4JvlqcoG9SDhASwWnNUPWoPDacNIWNooDZ3qJp3pqzLIyHAdYKuhdc2KOA18Ok8kyAS8ofEVnoQ
Fip19erwO5vPTJtQGTarWdf7OFttR3wkH5FulZWAV5Bx3wJK6HR0H0tv+npCTijDGg6ZTcLraKoC
D7/MYpVXkFC0lugkhHCrVi1kaHldjjLp9YLolwVhSaWE3gm+GqKj+VKesi4vqFzfChNx5ZKM+7dC
c6qaUDZDSgwTn4BM4JbEZbGH0UV531JAyiqakTCO8SqYSkF1rHB/GmaUbDrBA++ZDb1s2ios3aUS
FHLnMDNNb5v3jXLwqF97ne0/+UrAV2fS80EFhsYtujNwaNpjzfMAUuasbRvaGmsKZD3eFNwecTwt
U+k5BHPa0N2IuqFavGXuDD7Rf7lohrhC9MDHh1jglvmcCSuWnOPwEf6GBQ2xwPSNoGjL1w5jwMvU
O460HBJmT6Fk/ckeklVC4/DsWpUEjUNYfjp+BDg9Fg5roGxlBRNFD5kRR4TDkiVJlZlvx/F89HtB
4wd4leFXECZ2LJzj2kvRiPER+SdsyPqUUf2aAB6Ch1ImVtmG7Mhu4FfV79vAXJuZcU/KahDaTo8i
HKG6c9spSmSl6kBrbRrNmiNXdEq5A5YqmOC2rJVaXEM6CM2HRcI1cHWXVYkkuSMCxaXnmiTP1pEW
D63zzAO9yzexfxz8YNjtLLC04hId4RmQFQEx8NlKTuV+eN9ttEaZ2rqZ/s9gmTz6bjbVy+eAxGjN
5erALJsbl8pvzncwns5FsCiJ9Mokn09dsQmXe+jcfDpCdvdQuZ5RmExPe77vFJblcMhI4RlFhxIn
CzxZ5O40jf3WHoMlhwMYixHBBssUFx+3m0LxCrcNtCyDuwy9ZrkPROgrPMo2wbMhN7mxQJU/tOi8
YNXfA9XStDDDlMLwDQoh/w6PWJdO0PxIKodQyq706ngRJB1ywQ5dtZ2sgCWhSzh9hqxYCXQ6ELQT
vMIFr8gCaKneKo3V6ViYZtNNQBgnX0lyriPOTbXOYOiwO4uNheYH8YDp7JIldBnUK2UdAccyCUDt
Pev6HSAQuHlx2yzmtBcMy35awhkSxzy+RQqwBtz7Pb5jbNDrHb8/isa/4KMPZT6IrNWyUoeG+USM
aAg5O3jPM6I9pV6ET84atd5IrAP0bLfD/wqF3wHcmw08HD6irJhwp22dJnGUZlIgtEtpgluYBSSY
1opI0faSDMZ+cWx0iViQ2gf1Guf/pMHgSzky4BMFRD1DokIt8ad6olLVk980o8mo3GLqv0vOMhL3
PaF8+bO3ibvpJufDoFY+V/ARGyqrDozRA+SYuyNFXbN0ce8AjJr9gR2qTK4CPfnFzr24sw/ogJT5
H+fqETZaahqo34QWNsRFM+4nf8TOBxDtVRzV6EqIwt9UQU9UHEyHdreYoJVdMp1sw+pD858QG7bj
TNvONlSCOXvq+a883/iHSr9x1+3jeyj3WpChhMj6JE+m/Ls8oGpw2sfJPMcPTbxR3xI+tBRtFzsz
3GT14eMqJ9fKFrPgQNk1KVa35lg2WPG/fOHP5ibISvFF9016QjEaQsQLmF/vfK8deT3dcpPuaBnz
ED2boKbQ2iFi1l8jLG9TThqmHDvdi4XA6E3z+EJOOOgc0FK5R0ggrcqE7W4fXXeMeiQ08eo4TBN8
+4X4CBz4kMwznunH4SoFwrugq/M4DArYr8k79ymk7xKMDY++PBuBgIeXc17nMS11k8q6mV1TfOqT
IDkgeiL2CbVr9dGCHIpvUIL84baQf4wXrKVV2dxKTWw9HeZQ1AT6Lz8TbyN+NbVWkB/3fFM64NMa
d9YYvMoKJeNJ8CSfs1sk50I/CFW737D7+gmR0aNbLQr81mtdX0Ydi0UJZoLpqrDjhzeabflO4ZJA
v5JxL4y1ySz+Mum6pPm/0U8H8XXsPZehR/rZ9SxYHLFSYv2HY8bf64/pujv0XVky0HLqVMFbmMcq
O4Kg3XJIVws+YQuRbvz194L6hgic4Q7udtY3kQRIaRGTZ882lGvqPNLJ6MnrCm+V1kZqrnMoUCSb
TXQElQ6qgfxovUBnJSTyPI4RYAs8s213SaIb0JosKiSCPbj5hFj0GSzHdysUILrhgqfLuOrf1X+C
jihjE/piFc3IhYZ1puwEXNXkz2jxFq466cM762Cltl3LzXrP90kWwOuwz9DQskNdSiaihRdXNq/F
byqD+ROgqlb8fJ7OP0q5/Jm10sdl9w85AkSUwysph3eVSjAswvbauweSLgwk7GotLJulguZB8nOV
o/YAX5bA55QyBREH+W1mGjEuiTZRlKXi/fBrqjzP8lL0eAqhwfBeuFaSPujJ5pjcZcbmjxE2xygm
UBmlT4f91SJ6sEaGpdx+BpUTKJcOt4v5kvWwTGw/718Oos5jRYxVPgmVTZO2y78P0OSHFGVAUJ5p
4eofvnyIdmNELLsedG7aO/gzfQPCfqFtBKsIBDSIfZ1Uv1tqYwcQfIoIxxf2pAGazGAjRTrKyykj
Yk2s/2BqJ6f8hUhYOfUYu7FKRGO5VadpPQKQSIziKlHK8n296+Soqq0XaMMDEfSgM8Nl7nvU6Oli
Eo86DEqIiIht3GBQJy9vOs62MPXKigy/VMTVL2D+dFjvqwdM/iWfz3Hafd2civHd28soegcRCI7r
oMQeCS6QABqXJFscc9rjmaiwQ8asQcOEkhXaiSEEdV7CdDwOb/cSrHUOBLSwXANxzA9J6KM03qKG
/uWhlzxwUtqex9G7NCX6ThbwUgY0MDHqhLgk7gIr6KA8anWETZpwnISVya3Z7Ud4KrckJGCJlUkL
BfgeWpacHSeCL0ttkpCFEjIa2YSAkHnu1ebDaPu/RY3d3wrU4Qv2Jo/YNtXMB78b6ozBsV4Re0b3
UNvYXdsnz4Zn7e239wilrRWD+XpQstOWs+UWQQBfaYrcoWYwMPTyEeIrcjT/NYWjssQYY0hJAZyU
OaFLSQJnu3CkPgYbxfQL+cpXEfPOtI8JQrsu+OL+P462SG6zfEjD51de3CxH76AtiENUZ3oaAIA4
yJucM7tswEz+BOm/tp5lOyf4HyC6KaGLLpAbuD7emMCwm2cr73OFZhEq721/0T+xOb/Sq+KjgKt+
wAg+VHA80FJOE197JnzpfdtPritiehv3XqodpIWPCvrYf5aogiiEEtSULSybkNkrv6WgZHF4bowf
M+eNmztyX0RKhcJYBMezziqhIhR702GCUW0nXEvl+lHLOgVjaPICoxml0yfJ9Ir5NuWRfNZrbTTA
F3LWe2A+gWpLCWtKJv33AOozsLGkEEDgrD5088OQPxiqIv6J0FuhxVzfq3GDpM+nzu1T7UHNptjs
LcHJtTgbnt6PxNmSrMt8bslwO7unsrSa/Gc8+hHDPZy8DNYAFEg0FuYhhUzLt10GXEEHP823emq1
+dVLsX7swDxl3v7U2zLbancJraNxkcSzuIDcGtHKK2N5aQJp3tY7JOFqFoxGyVh9ohLUgoladTiW
NfwsYJhqolAancw3EhWytKbEpcU324wuYYTPm2lCsRk33svQqyorl2cKUki2qw8Ly2qDDyTH2yps
E1XzX1H6WhgjYrcWY8WzVnqdf+l69mvEPGXHAYFyKTflbbgaBnUYYoaiYL2hyPVAcUfD/PjryXDO
C1i1jRqm2Ho//Sdoe0egr4EwVrJ0LJTVz7KM9ABxRa0Svc5ivAb91xdXfOD5J+mmcc6jCftu/R9t
u0T1YLYsgYShO1HDigow0aXgLP8e83X/0HGxtVBokzY+HYQG/lR5A3aU6qS9uwgB2Ghf3OPwTYfN
bNd5DTDC+tWKBnKbbzYuGD+s8JsyvzI/to7Pn3sMFKStAiV13XKfnT6ZvpoGGG2usSfLYs2P4T8D
Vd0iq4xU9pz4wdjESZfLIx8J3e85r+DK64LW2GWT2oYAN0nh73eEzylbgnGQuBwucWYeT3jeTWaX
GFG+bjG+q2xb7UZhx/WnnTHm1Tk/jGQacRAf5dAxCrTbdXGGsQGQX6vUKH82bALp7ESqEp2JTBVD
NNxiQLRCYms6DcDiVA7UL4gibCNolcs6gvbxaNszHyjnLw83aqVWLyzIlv9Kxc8K4vzufz+mzW8C
gM6EHwtykjq0FETSxPa31viYfHs86ff9GRC5EG7VUmFY1Zn9r67EY9YFKboCEz3ewwTVBq7gJozK
KeiB/ALJcRcyz5+uU5/jUGxpatyGcull71TMGqUvFAFGz0a+71ZVyOncSkvPFws5ijH1YMaeibFw
Y/j/RrNSSA6E26NOPpagt53jvpN8O7fptK/LqZNf6tJgft1s1ZAz/LTHD6H6dhibhbHPMEWP4crZ
r/JSzjbQ09bOwAeMx8+LNLDuwYthTNaWlZBsYoEqw71hASr+KsKFhl3/KoJeRHzkrpE8/WlJumOs
LcInvN6dH8oxEPGf1N+ACD8qcf+WBo7JIlnel4kbIKYHdDZYFxIqb7AOn7/k0/KcIpoqCMcxSISg
f0OFRdXTVxCrfga1bbrpivjn1Fj34QvgvLHhtQuaMYcllDV6VOJ4+f1Yw+2NxR3sOpeEadRD+VDF
iQK5VgAr+MU1xb6BviV/Jjh1H3YOYdwTeS/pWlWYQT40eJ40mBFWQX7dX+Le1rsRbf0AFL0Za9dj
4YFjy2euJraZ+TFHoWzEjc93PK7OgOG+iKprgv/tIXzSbyKLZk66TV2iIVH6RCfvuoqU1QSZJ1F1
Xb0whtr8DNvhTpfmWRgWfSm1B/AeYgQrlxegN0oNK1lfXxC2hzgPmk5yesjDAkHJofHD1LPX+sLa
e7Jq0zt3ClkmWOkZ/128KN4D2o1o6PLSGKk9Lmod4AQPhiVT2uuxnQQ5GzTPa2y7u+I+WlhzpICo
OypxqN9ItielXn5IC5+gxSxGbkSRsGLWCjUokJsXNGDHV0Ghd5E8croF+r1Dm+UHjjSsIei80QXl
s0p3pKCXjWLd5QwmBw6LxtBGQ6eTY/WU4mlaZVta8jnqgok0mhteIbnGpZfJtRtCQ0nEIZK313/R
xHdsMAE2IiILaUljT8rUj2cjG0vfODkLWaCZLRyuvoIiDXaZY1wSHYKAO6DE6uJyYU1mQvy0vEPb
pSRTKTIbReA0Uut8LbDdY0pk9hDzsFCTEXh6RBVpKfh3pCji+eS43NARLnsnQrpAQd/64HL7xLLP
dPb1KNm7hy1rj4O72opsOFJkOG2Fn49jYNwRTT/tCkFlysk2RQdXMFg7r1GUIILf+NQiwtXZV8gT
SyS+xjPvfiZk3txwKNU5ty4aT41glJj+mMpmzjxfl/ndnDMFnybjfsKBNvwF2kncqzz7oxg5qDoa
HzjnjnabL1HL/NMS2oDrtmwYu4tI431dtSVVkamPc6+y0+RcZEuP057BI+NvqgF8zrNkqQeJ702r
7666L5Z2TmjzGTqDyOU+VDXdZEiw01OCSgTIf89e/BIKD+ZZCISrCN7mJLrK64pdhPpTdR3SFx3U
8dzb58BBWVXKzRWimo0VvehkP+zaQw0NvC7x1LOGB2yDGS1HVJ4rdW0n1zmhHPKcPqEza0EcTyMf
7gGy3Ib84tiKvA4NCm4268of0nlMS6o9m2JR6kxXSQiizXoFyiNLpL1njYTM6hPF6bokRzA43Hya
Jj1hd0Xr+2lFhhYDGq9SOhWybn1ReoTGbX0Mf36ksanM+4HS4tfNF6mu1YGRowHHe4NEY1KZJrSD
roes9ym1v6Jnm6t1Pq4vR3fq40BpNHH1oJurKNY0QGq1gi3IrGdRwFFFwapEaVeiZLMPIP5p/QzX
syxFWkmJNSHT7i1I5zEyYzfhOGdS3jmDU2e6jKY4gck5ZbuHQq6FOL/e2LlwXqa+ienJZEsZqD2Z
vsRhqb+9/FvOG0qyAHWxfiEOyErXMUZTDbFHZte6YSdaaQeMSxiJ/3UYGSqIWnJhgczyP1L9DBnh
jNXUawWcYBSJ8KUlQuQROtTT9UUmpMurUWDnVDRpPSIHmoNghah2PF6zzPKqkIfj7PCELxwTX58w
525tsPm34hsl0HCes0WSFRi7fpC17nR/2AOA00x/fnJIg09K3DfaH5QZrUJgOC5IcE0qF2WRPz7c
lmXtmun2Jw1/s7CU6+ghBgndHPFAX779cV9OswXCDwLO1xnD+TcaaKG5jGW+2f3nJB/WQ9Q5NZpF
n/lae8DA04/5V4BBWGfGF5ySdFz9KevJiSnXX9bB7+klRoUxUW6rofzx5XZkoCTf1ho6tZ/xSyp7
i1zNdivJUd/eRS3GtpUzvu1z5p5D6+vYJskNrcEf/q9mcX2r8xh8cgP5FyZ+AbliRV09beBx4OgD
J6H2rc3dpeWizAu72r2gUj3rSHLMXEGFPFqDf7V3WJrQm5Z9LLbwLR8Nm4oxmFK7lbcvgCDY4yPY
7PJ1gJn5o0osE5C2o+2iygY9DYq/eha0cPDqJr3l1Z+ZrDl3JuT/YWiYFQ5zbIO4q1PvIJNciva2
BmMFsx/goxMmtjYIb1S3YQhHOXtgjEAH3StyPRY4etZKtXU1fcY7Wdtp+/D+XVeNa19TGALVX42m
5za8WSryUfUKEq0GXx2yA8azke9kvwNQmvOMv9BcaPguhXKVUp1uxFJwosNCub4uTvFxLmZeYce5
itj+wjVpwnhEtlY3qn9zYUhGUUs7WUKqozM7AMqTXWWzvzk79jeu4EeEOPUAH/DhWGjmMTeuFGuL
dKBfGCL/YrmCgRLG80gyRcbTnSEmz2ND/gGWlYUAWeLWLM6r4QhVv3wqG2Vd4Ff7cbqUNJMek8YP
hEuJlq69cxypi3CLgcWyVT1Ruqbk4PRRKz1uAB7LXo9CfgXEPjAe2wD37EIm7pCOSnqYVp1PLXWi
tQXdj7MDzesVylKg4czmdf6PNYLrqddzRrc0P43xlzqjIriOQ6XnYUPSDR3/mXrizlfB/MLDcmow
MtsC4CYJVDWmM0cJDJ/7f0D1qpolDt6bS5HxAK5kRaph1J8qviNK1hZ5j84xTNq/3GviGNN7KXPM
+GXckLEun7YjHdSK+K9JBAMW1j7lVOp58bQb9Nwe8FjiR0heEXe3fEgXBzUKFDEkjwUbpO8zXETk
udQG36nS2a8r7t/CB1Hg+aOndWC5SIy0YDeFr3Cqbk6sb7ugUyFwCNIGESqxDOJol+vHqx3jYmLC
FBNvDbDXUd7HLIXLDSntKiNsSYNANakpYftllu9wu1A7s5x6wOSf9dBC1xG7cfIvtC6sXMn6XBWh
e8JONzv2yptZLsGnrtSoMPFmz1r7zeqVIz6YbwlAKVezzE1UG1bA3c/BscDgBbnWY4BE5S0SmM3z
fB/AaRao3Gbq2JV0VSMgeTEiGvYCNOgTB85a3+7x/zBqOyRb8jpCYBuo7dcyTm2JKCgDBvJoQDo3
moBKuaZFb3R4mR3jiAWZ4h0zszZZSlN8/Ju8B5AZE0c7qj3R9L4RS1Fl5s7fcPS4IPKbId7/UYbn
cGSVQehrKIaNTa5tr2zbBI8gIE4ju9WEllgPYJOIn4IEEXv1HQ3HbjCgEqq9NaUq41mdt8NhrctP
e02ciCpq0768vXbnUDG2T0mFs1Tnp6VoyLlQTlJwfu5ASNQJlHqv9EErlUHzCGjs4kMo7UMnu5hO
xbx6PAxQUtB9apnj6CQdIf8mAYUoUecHDbO4FVw1h2WmQ9OcoQwogjnRaQxOagZ0NdfmFQsciYvL
Nxm/GmXMsDUOZHl+5SA1lfKE8JbQ4X5H+RxbOTH+zeqkR1Xmy/uDSJfkULcwYqYR450/69unJm9i
udHXQkTV50biFJtefgUjPTWoHNMnfERyIKElEXO0/chyGo+6+xQiG+xvVGFJgD9c7sl8XFFV3Guo
vuzbTRhL0cL3wBhr6sfDaND/Yq90dxEhCRXlRZrlfSaCXXbPaBjxCbqeq7UPPlwHd8IGVZCf20g7
K17TZkjhcBFjy/bP3oSzes0AKG0IQFlJzHaAcJN0QWqLNUrdSxiJrzfJf3wUr12cJVwVFqJYGoFW
pH5gmdOCfOGF6o5BdZulJurMK740AW6ut7oujCsbM/Ucb3dfD0FuyxRCEtEkS7bSfBQCNdfoXE0C
coeAOx3vZrRGDR1n0aIuIP4yHS5tGW1gADbGV72W/OrKPkQsLT+Ry0PjCENqHYL+xghNXSXPl25a
m3cgQ6+nl+5D6PqNK1+zHeyjcZ4uVjjUHqhNi5yiT/EEP9wxY+nj+YKnPPgAJ0QXEPl93pmB0rHB
xX3xiSSzQe/UhpK41ltT5vUtch069+xxXomvVxgD+bbA4+IFCMOOCean2IiKvx2lgLBI1XQING5K
AwG+5EfEtXnPZopguq4yCyknVBck658pavM9Jv9IqyDcJ7JB3FxUpOAmIYRUOXBtKC4vhTiQGF3h
FudotNkcEFjop6xjWKWsvAZv+wiot9iHbTUwCBp6KRrW/jVxMcvPhEcE2f5UKPZX2PCuLciX5pMj
+G5EfkIQ3PcfLblobAZKNxDQ/cIfF7HcwIzsJdL1+HGU1Hz5ax8zoRp9wNEiF6JBHRktGE+j416E
zbQv245iqqdAerKJ3TZDFI4VWQ21IcpGdMwsFLPXVHNpzLH397trXPUPI3Eq/XnjfMwDBFrS7HPY
OOCJoxH0a5cld3IjxlyloonD5g5PQp0KSVFzTCHN40mMzw8rV7EfHB/c0NBOXvxRnUYHO3zeoDS3
OKvbjA15WIgKKPeorEuxBlb7qRgBIDtJbJhv/MVRUhzDUmInVB8CXPevm5ceGcbOsDe7iMpl4SIu
M7K5tGIggNXSowpQhzH9sdhA8iEfU+jMbbKJIpRKQt0X+jykfzFVNw/1102CxL/bXBcgHxzZbDIn
XmEiHH/Ds4DWNKJvQQULgmSpDzFyUh+Ua56ZTUGKk/Mkb1ykjV6QnVXkkJMDUnE5lThMyvpxLPDh
2m1doZj60nWcB9ZNG4S3icx9vkblnNESalR/CQUGOZcD1H084VKBKHMMfOGb9PqaOXCeJzWHBJKB
5R+LO0S+YUnb2fP64qGrXLA8fmvvqYW8ch7yTMv1Bb9btdCmypRaSmUZGiKl14To/2osafKZB9H/
EmUKBA52kMQ+ipxjeof9ukCe5GjDYl1g3zcTjcfoaQuC/c1T3jeyxhIzpXeTaJtsfyX1n2TGHsty
oKqZb4Ku58Sutsi23aFBRXKyMDHdJisZd//b5ItJwtiXPQ2uhuAiFcGLQcQZ2GxTwimlZClirtS2
9uXRETDgJAM1DZFtTSQem09aJwoasoRD2OTjkWM5TWNcjPOCRhHpPSEcd2VRAA420yaSl154QppZ
8728vmL4P0LyFmJgOq37BGJmzdRWfSoeJd9rjM/03O1sgBi1bRJVgNw2yB1jzZo4XmO9n5gakXST
JiBdDNBnED2XTkrAqyaRDYHOeTQ70tpk+OXjHWKf5SvayDoKMTAFo4hi80sdQeSvAapB/q17L1Yu
sizNcEWGCDBtOTHGXL5XZZak/J0Awxjqt7ZIFzAb+Z6oXshq5oaMppIcgqzdBwnYf6ML6D3UHgDa
YeGPKbMi3gFzD6Iu3n9JQgvJR2js43AWKb9uren/2OsCZ/pXT37okrdjXHEmkqeGMvubXVeg9lDy
8vaqxDzcQm54AEzIinfaIrDL8u9CmaXpuyc7ruX6KxMBjmAKAyI5fILtyuFpoklPpVFsGunUlCA7
+LCCB8o9kkXlau6nKoFhUzCSKmYd3hqdjZy0ze0mMoxwU7PNNGyfetvjh9pIlJaQYqqpMjpF5wae
SDWlO6KCZF0fMEpcgiWqoPRLHneWdca7Y+K2lNCF3RV830v6HLhOls38tzYVElNpMbLcF9McG/iy
J+g7b2WYpqg66SvY56hNxd6+dKrhs/Q+EyuwGDpXUF9yEbtSOGJPmU0bRSXwBNeKbbxmPFfv9sD7
dXx2whIzClmqGcmfFJp342LbswHRozAhqCJfkJUEUKaI0HkTO7Qkx0CYY8ADlpUsgtZMU0EHYrZT
Z6U1AVSh926hkHRpKAXcTvVpYUsdKt6JX/5/k8GAD9bf4MrFusq6qQarAZvdhO079ZDAEwR7RKt7
jcsmCiFxB3gOtxjgo7PgUYHPPx5f00ZkAn+E2U8hMNY0XpTWRPkw3eJQ5TNMiHGsQ4IkaTIOTdlI
ANDzhBQ6MD6HXqtjAML/Lr6VNLvDILnCLWvr5ON2uAnDFu4RqohhPj7QD6qPhNxFJbs5D1gyrH1s
h+HkH3XdilEAi/yA3146b+OaFmABfJWNXU6vLhCLGpdgxX7HlcdfXmt4e7eAcelzmgAgyioB2Awm
2wuPqjdJo0LBaMwQxuPfTen4O+QjDm4aeuZS+UTKv4ZE2JOlhN31w3oYDChDOVbZ0HFb0T83A7rw
HCkF/J7zD7F2SDPNc2cNU2OWQrJJTkIDI+vC/mSz0l1ZZGI8E5n9fuKbu/0Yxb0j8Q0VFzd+gP41
6NqeCCmi1Qq6dkWsLrlOpyd2c5iS5djVJm4/H7f1/kDB5Dh5Qm5e6IPFyRBxtLD5xBWk2bIWtl1K
pBOBJk8SRegEECBfiBPi/wJvnD96SrbuiUAX3jIRtxecPB/zHoB/g7WNGCmYGWcrzYYbqdppemmN
4bWDUPGjz92Mi2QlJP/wCwB78dulsXe7r3V7qBuGbtPn8jotsT3i8zYFtHUGU5dlgXCNqy/AYZdf
AYKDb9vlD2xdaOXy7R2L9u26O3klLTqh57WhcNLDVRJ0od+Ne7ay9sUuDulZm9WWbodIew7Bm3Dl
iBojTVvZsZe6wUY3sPsqjH4pUXfbvDlGobDbnX14T6g/lIXU6+W31GePMOU6zvwYBAP4Y8MoqqcY
jYYXv+eUcBGJdUQ7+HR2aedhT77/7PjztcR+6RVTy2gPf2+jymObSB4r5/Y3JtWgBUFpzvalOyLr
WVV697G02Q5E+Eb9ym099W6rB5h5NvNtJ9zgdeavm55Pfc6ol60okjTidVK0ETNfqhejn0E4aOkh
dirxrZD6+Is310hW6P9WH3Yj7grslNtnnsqWusCe3eaOGkGtuR5+F8VD+6QAOkzzjTbLTDO4zHsj
F44Gas3JNiSEow14MlYZ/zNNjBszh20cwbgnEbPd8FSypmL0rQXOb0I5Q6YHAguynBbrtevH0lx6
pCsVkBM1waWTYPIIGeoQrr9Spb6IJZTxpp1s1wCzgkQY1qRD+O+GsRlaxTgfo4TcTHwYV24GrCbX
icEGU9yiV5TrNVAXDZ66IboGN2Q0VYDE6szoI+8RxVXSAWw7AVE1TgdWGs453Ey0xJNJ8AeVHIXi
6CBL8ZuISl7mwnkpEZuvbIMoGWQwqVPO3ZL/AZ4REyGQah/i7ETwhzR8Ds67L18wLIULFE/GdiW4
cJaeP/szUNaEP+4/9KoSNaFc0q8NPsXXr0CP/RzeejhBpuq2XED6og7d/5YL6o2jISX4QqAzyK7Z
lD+uzwFTX4nZ6KofVUVDUTF3RmCZirFNVFEC4ZV+qv4viBFC1ZEAwPpXJZsLETLVAQEgcukY6W9U
/hhT5qr+tP1yr/bU3i1XOKN0V47uggDm/DDzfbJvyEosZuFa7PiaBTVUlED68i0bM+xTPS0+VPcY
jrl8zyZb+l68Z7NsxnxGDH1kBbq41SGGzlzn/hPiwX5vmiZ2PDtmhTIxXgiyXQiytvnduDXwVvI5
ACcu8cM1/ejNI1sc9z9onsXTUVEdLaJkHXdCmE3Jn/ij2b4POBd/P6YEOPZZOkms9eLYUUqFClau
UJg5JiuiWVxA1eaZcnAaiUjxPniWyJI5EP4iQ4othdvAsnCIzMoSWhU5SsfX3dmnIMuOpb8mO3+I
rf5NILGKuG+6xPbgc8vIBETErUdGCPEw2wjmKU0A8DuCzcFLIiIluBqAzOvRLWZf1nQ2SAWstUKS
Si3W6ev7U+tqMP+W1llyyMqi1rUKBSzgdd6g/SfjjgAJEwo5a4SJhE4jGQ/RaQXPNgwqcidPkDvP
UggkkKXYsLhLjLjmY0lLyZ3njUfd2VXfrDHaNxFLuBFRy7AxaHCAMBVkZkU3mBXFyq4oo1vbKw8f
V8EBcur87iLJIjpj3b3KD9KJ7f+50hQRaHKPAlSSr//3eeHpT5oEVqcCo5KzTaMH26FTFsxcCKt1
utTcoBMY6qDcee2L4VrW4xnPLh1PNuh2zRsPR6KebIfaPAxIl6DM+klzfT7BA8UQjn5UIU/Fdjl/
cZaN6m3+tKUptOp1JfIj62y82dSp7APnjVutJ5C0UBxEa4hlKUz+agVK1WeKtarsygcRtAOZnprU
cgKOfoF3qY7Ntv3wssiwqX7cBZINirJaj4Lyl1GTmGvCvhRMAGewK4EDtLiU/sRJIKwKDRtiNUCZ
ujudUsIYmS3mop04ZhjE1PxlgHApaE34Tr3HvWOG1FuT5Fm+vfzPD9YB7EJIL/9ln663OZOhxzG3
9lAUpcesu3VU5Ize8DwGZYOr4b2hoBrctUSVIR/nXTlN+uwqwPgsyYlpKJIF+S/uUOy87w1wYCf8
F5rnwUR7XtbErOXiepBcgUlb2v+dGHBZ85h8b/0ZQ8IFhiDVrm+yCSv/L5X+Nmm0LoT/VpkXQsFD
HkYBxKGEWuDkKP2K5qPTynYjaEAUTe4IvU1cmFUGlJnV9E6+JwgJYU6XFnI+Wgw2uqJVxgfFR+zw
PseTQaAtjGBt/U2h+3FsCOgfBOoEdBJ2vSvnabc6lB708tg2RYO7LsgwAU7eWctDVuIqvdCC1kIZ
wPw1ezYeysrEkYi1+YG06RN06WA8cY0wOUqlO8Q+yWQPmQLjD2Jp5XEf/CEKAxPOnNuHvw/e0Uqr
WSXuZHBmTPuTilzzoYhtbU0F3tzUls8wt0HXH5u39bcLUkWS1+/VWzCEik1R4h52ALbGpLvp1uQY
JhftWfGegZ+q51Mc0/5vkaH8eghxuJY7Ykeg4Y6G4VtFjqd2Za0blSWTxNGYkwGyTx74N2fERtOW
EUz9pI0vvE5GyPDxONiyMzzM5FRmlb77k3sGG1RIhNQvBWE//dX33wOqrhpbq8TUpAi+/ivHYcBn
Q36r9ORZUyCr1aBJtTro/z+ldIBh4L4jrtQ2uYlDPVz+Eb3b09X654cO6IRm1MwezTUu+0FawgTX
0QRJm1VN3DQx9dftOFktNMetPlvDNIJ66wRDplbgEnf7Wc32TAYwIhPbq1ham22NFqyP/GRFzalQ
I9xQIND2pkDt+3pqa4yD/ULU3FzaxNh9E5qiE4/n+WVEGwJqEBZwOb5uWU9XkOcA3U5jc7Ie0gq5
rRk+mb8EEDMYWyiQEPbz1Mff0B+qtaaHI4LluyOv3PfvfG9Xmh3M4+HIhjGBv9k1M50xx14bMsgz
S3+K3sS9e2Y7fwZUdtHK5ewp5BKU6dW+gZSV61rIFmdqexCOuTLVkf4YVwn2aODMzd0+GrRyIwdo
peCDBrfCKu5QZ4A8abLSYjT4IYxKZ/97hF4mPkWyiIGWREiYX1J3btLjtGHtysUiOmZKYwYRlHK5
4Wd13PQL08UsIosAzUWdMjeQ4oUuywbkQjho6D0WarQxVvcSdClXWayuYciPwHkRDxl7HzqUB5D6
/PRqUbqD71RfxBwmiFlFtKdgfyAYauiRe+vnR597HPu6E0PaR1eAzVKEwqZhSJYHUx0xq9TNL8Ac
TfNPWNsPlBdiJf5JIgPQW8PVfjGtxPb8UpJ39nuq4KD4e/i+A4P4pWcDSVD9eGxBnOj8n1XqSt/5
dP/6zDCKb3GbYwagmtvs1O+QaiSLR2oSE+cDVkBkG0YVthpspsz1gnduY/nG4LX1WNP4vLSHYAh/
G3RQB6EycNx1SGc8Jw6jdVmqisoYH+JbErGnydB3cXUEft5Os9RffQpr2KLRsfP4D4oSBMDQWTHq
B763ETPBo8gwmr8CxTNkfqfWLpKioKWN40Oqc0RXaE6CZdkV9B35JOM/zT0lanqMjMx98ME5CZug
b6blY2nuoOl/hwFOMDD8Dh7E+EFP/79OX0VoU8fj0RaKblujDbC5mmOOZPqk1Y3dc9J0MmAcei4b
x+8odge/2IRH9TsNA4OgqQCaJZ7A3wwO3YY3ZbdMSyNHCppfYuEMWyo2ZKtXM5Obz5m1kagXcquG
xsOX4Hcv4TrC/+2efJCm6BQsXiquLd8aiaCrxAW7X/g9KRU2NHlauPU37iFCTRmGaIM1+nfdtCip
VE6B7v3tc064LLPmVY7L1ESGylUbyaKMjve37z5Wv38SVnt2AAiSLn3hYczmxrMtYoYhL2Cyy6xf
RaBhNx3GIbOmFojzil6/mLSRKzrha8KQsSgUS2q4Jx5mYPSsPWS8F9Xz4K+IpJnb96qdfQChL/gv
tHB82WlzF5fSRW6iZP1MkrUH1uM50FlozFDtNxOeChXK3CnPAT7XUABQSxdYi9heLL2Ah42mDLX8
1FNG2Yi+bd7izEt22DgLU/ffnH3G0MMshn6lzlCYzxmAWIbn6Xi7RsCqiU/4QdEDUC5B5xqUE60X
qnxQBakrsdIIwk7gWPamxaZET/90IAjOvoQi/Eth4dIoxdjICtPrynWIp2OGPlHL31FBigaoohmw
KF0JRiHiqyaiT+ViThbxpfcHKM0P3D8pZ2U6C64FMmRgo7GbAuZiSWDETc5A1NwjcBW+n51DUw/v
E8WQx6Nn8pfpYbGz9QFqbzw208YIpUxkTLAs9hjy5y/pOX3j3dDY0leiWnqmHx2Dk11zctVAYZ1a
klV7PaOGXb4h7m4+DlbmT2ie3AYTG7G7ghSFp5T8QMWmSomTmkHEDZVaDTTLcDBRhJJjcaDtxNK7
0r2UdM4iBiAP67P1i3RpVhPFwJM39ho/yGx4YE8Cf966OgIzPn6Bb5CyAHKed0/hxpH67Wa8Ohho
eIjR8kAUhZJgCT0ml75HXZkPJDicC1VLohWUPQd4xAn/1nePXNif2jvM/y7DCZuiH2fE5HOp+BNE
zA3RSvDZSZhBUyKaWX0BjTsjoehyKTln1bsbXWDX0vWBLQldKuVFaqdgko2kA9I4mG5m62f4zX57
5TeUe00NvBNZvPzhozhHKoc3JQuUYU4SbprZ2aT79pB9rU3aGSyUJ02BlQrH1PT1/+WR3u1DH0XG
p9daTwEXgl+E5KxUnXxvlO5L6bX6LRpifnvrAFARxJsc7rDv8IbCMXhodmh1EeRvpnqZ2ZkTpb0d
zFZdNN3q2UjbPiqoSBaUqHXcGhcnDjhaa2LLgpiIfiy18eOiumhOX34KULOQdCbWLH95dtHq3WfG
NtveGZmW3HXG6Q5mxPjKbWyXW1Xn57Ju5nex1jrjVVzaXM7NK4l2KgWsrhhyQ2Z2lbUR7Y7VUZaA
njvMJX/Fs9j+zAWxF+z6wCg6SilOFI6bjGQSgrcNibEF8bsks74mrcdR+U9Z3IKIAJCMBZ1D+//p
sduXhnZhHJwDvKsd+T9g2tIlWCbQcOrcD0SJUezidRb/mvl58MpyPv9ZEeHu8ZvnxjoUnh3zWBe+
iBML59WzRikTK0DIuOjHzSkvABHL++iSX+2iWS5ldz7GXxQYTND1NwNZYAMPdli6sGj4qrmU1UZA
rzupGJF9flczRU3HQCJUpQah+pTUXEMk0TIm+Oh+jLd7+zOJoPwwX9FO8Wsj4bP6IuLVoD0wv/nI
IZilydUb06Je6Cs5yMoBT8Lh9KrMKugnKaXZDt0xIjj7u5LpYIhIq979svnJjyhibdpj0+dRrp3A
2Xbzp8NHE6YOa8NyGB1cGD8MZRWwGtgl8ref9VpyLI9l8IXMjkngB5JOrmRc+OaAFGsUKzj/f+gD
ce2/KqKSDIJ8+8oTpNQZDfMWR0cwcdDYHelA+kTKRsUHywbyJ8MhbwzHmJbvPmU/fTf01LbrwDpY
0xCSiWyQOdbcb+pT5trcCVXlWWeUkAjUA6805aF5qE4qMlNULVjFizc/KicW/I0xmNw3m8IlmEU2
SsuSTluRpC7NV3X/bPBYzLJX0tmBSD53kwBG+5BW1caP4E7BSK49apcDv715jqnDeYbwPdpBamkh
4VWN0wzS0imfZjKwn6uGEaJ5sEVrmP9P6rXEdOXHEo+Rruu0Co0JcjDiJNuBJzbV2rW+orptCQ6B
EOqSOoi35QSbmo3QkP0Y5jIUMA4Gr+IyR+Hbw+kp2fRW8QjKl9p9V8qUY84v1rEMh7N50hx8n+qx
674yhqdABmVa3DH/dQ8JZbbn+5e6VvcpbqNPQqc4dHesyf8THVpFgaIMx+dHj2CySX+Q10MzM08T
X6ayCNXk69RN59jABCsD8155fsl7bTRXlvCqAPQOly8fgwpo2H2/01V+zuNUxOBGB2wrYW6Ziq6d
8X3RQzcVfreUw3xTX+uug74JR9sgW/GUcsDtCZ7HlvG46zaFsLE4gyBAQQkUin2RLdovE6ru/7eo
tt0T97A1YkuAxt7jx+izL3f43NjrQqrMzT65wPJB6eSPNthzY0epd9Ki/DOMofjfN6nKDBe5tT7f
kIPSHKDto0Y4T1zQbMhxRrplLm0yT9ZcHZK+CeB0xGCG2FcfS3IAl7ic02l7wD9LWRrGi1aTsLJu
Nb1cBIWPeAjZUceNXYwOZFNhl6yK0u/YUGmdn8KPiU9ZX6VHzvqHUl7sotQbQHo/N/BoewcjZRNx
Dc1vevA2E0SvICfmm75Fw2B1J2h1acPbw8hg/zUxjL4WtU2zx1SMT/6a7soMQNUw/iQVMlDhdLjF
lkho0tdAv1449RLG12Q4vB6YGPto2BgPptFgKTWVZdXnfVQPrpDYjzrGUlG9oGgSxQu9qOOEPfBu
sin7QtklffRYw5vLYt5GnGcTcPMqT1R5XMNerrs/3v6TRuEb5nSXc1fvHbJmCdYLNrh79sj5GTU/
p617PIaHMa5IeixzzUn981pT9mwOhOHtYGA6ycjuax1mMl7qassjd6eHm7eWmY4rsxe1bi018pRQ
lh1u+EDvVKcYn0Ihq1bGLTZXYmAH36a2XL3Wml9mz4gz02zePyAPLlqauUC2oQ2zGMEYiiwLSoj6
3qTIRyORwReHo+WasXFi/uB/qRS//jSJTJqx/n9gcER1bF8s6V4W/im28mr7Duteq2cIB6UGaXVN
rxdQW0y+QhkOCL9YU5UDuhnIVT+2xYxP9tYYTwUYEF53DJd9kx+i84YRWjPkgujsaIQ9poiKOlXb
+dlQUummTP872HR+SOmohZPeMonXIIvY/mwCJlD+TmaLquK7FpTF4tX7h9n1ASrfTdKhVxJA5cFs
ZfQ2eCX5W+zxSFaYJgcuc5V/J0Z0D8++mMedF54Rcw5U9yMa8Z0NPFVZYpx23LYpPNjt4DOs+lza
gDvWnTfowWu4JY0EOcXF1DRC6/OitIRvReNr3bCrvbu1S5rKZfC8s5M2sjf0Kfn+XOGF0KVVtJsV
jOvtbSvAuuqbz2XKjjXqVU3/3kBjNfs0FBwQvNbelvGmAiSzBqpG0Ku0q3zut8vVMp7mGq4ghfis
CthxSdGqrXAfnJXOZnGbrCAG8PaAWbaUCKKOGhlXDDu3Z8sfEPcZHD5PkqavoIQtU8x7aqO7ALce
MITtBGz1kfvGmkOv1pI8CV4YD6NLmg9eUAAKXuDEm6vho0wa3BBoQq26hBg5xjUlocdaCA7NITOo
dbjZY6GFkjEGIMz144wHf4nNn8P8QRdmwsMpKV+mmRKsHeBsBYPyAGXXZWemmOmOE4V/0StDLM7E
YpaVei4y9AeioskCMpLwdX2P7MCnIEBYPkGw5TOCPt0WWY1KGJg+/slMxoWfq5y3dXSJbTFHyD3j
H1jLdEorlufreoqEG+1x6sk0DTbhBfg4fGdE2wL0rqShSQgz58q2EcyLp4BA9xDhSxH5jnwF+nCN
a6bvukT4k+W6Fveb4RBermLOazhnZadncybArAgjs11V3Nls7ZMdkrzFsxSXQohOD44H7V3XPp1L
y/WKwlsZjr6zpIRks65lz38kzfz8SZ5RVOFcfpew9D8og8OEQ1PZ8RY+U6a6tc/aFPUqo++NVVxt
JpVkscIf6afA68z4LF6XjX3ZtfR7wTLQ8mA77fNF82nQ4HSVoMR2P4UOe7NyyH4vOIXPsSGhTiCj
/51uYFPp31M7oCLHHEwG08mAMr3JV8LMWeMnRsyC3gR1XNksuKFY6Dvnmahsd4s8C4mZzOvRuj5I
/oSntTkC+68WgUv15E4KjuI9aSPHaBp+GeBi+1kw3YKNwNw+klxdvtEqCIlJq3flpVlO4jSVxJty
gg84Ksh+JRaIOTkkGY0MwdIu25NaD7e7seAUODYwc7EtHcCBGP7AQz+y0/+zeDAxaOAodnPTCB2E
zHAqq1CG4pLR+xQ8dtEFrl28wkHAQBzNqmvlP5VC3yvrgnNKkPqCS3gjIIzSKZFGL1SrNlXNe5/s
CUrk6U/1S34GV6q/UfOPEUHBylixktKYYPPxNNbpmoVuzJHLjGslLVKWTiEbqO8GN7/x7DP8yWoQ
zBX+ar5yX7s9r2G0fYzOQ3pZY6XkZwNONWgY3SrBJYD+bQVhYR3dVhvXJZADajYcIOkLooGG6B/e
oSfQmWe9izshBgdiZzfFaMgPpFET2EchJfjftWA/JVTYLIBc3Kql2PFtCgtae5uLsO+NorGBXZFP
s0FUnZMxHoS8QZExYw/rPt8Du1AGUMV+zeyi7uKM/DuQ7qewDpuBVuhhJMvAuZYAj9LY1QVIA0Z/
PtGbqcujQd6r+yx8B5qVVy6ZY4TEAPOodfDGanubohrvAns+HT1XRw+Pcagsd4qDjphr5qFNJfw+
rD3Xrp0JqGv89mWKs5K8HB+jzqSUY04SZYhobPf9xl7pbythd9jdFFj4OXSTuJ2Cc20xXYVBIjcS
zArBHLCkJ6wi9Hw98YPGPcwvAsufKx0fLTqZ2r1d6WrPUMkXSmPKvWCr4DAdnVD5RX3CuEmrXhPC
ukKzaJxNk7TPFQmGcprj9eDZHQlaM7eNUpLkWfPlGlZsn9mt0blI6jDn3vEPwH1v0yDZ8IvjKTq7
6W+FOahXbP5HntS2vMkScv5cQ9aBwMkAdYw7p+A50b4isqCr5WiW4mNN1RYZGYC+id4GgU2WvmMT
EoAu/DsvdDSKcLYOZpJTFUbdVCmBvtySwqioiQNw/W27GHBdAdVVUoyQwP9FqA/5X+/kAD3R9kaW
sUzLQdjkJ1cZIcGCEqy/1fnJ4UQAJt0ohgkXro3ABSZt6yqVTIUqQRztqCetN69c0Wkf3CAvjRMk
MA0OdpXhA9eICZjzVNGGww6eDOHIKuNQHCBZBIDq1LJXWCoHGayD9vrcTGRf5ptO3gItD9kyPxiQ
81fhs5d0ztnoWer7YUBz3yrqwMuZtiP3urtYcmewrGtZYCUxSonAasq4TxolfVTRbpQRJLsbskn9
KyXX2tjpVbvwPX/g+6fljLMl55anHu7NFIZFqGlYkV38czGCoGDaPBejgoCPgBXWxvRONmUS55PK
eKq50NekQQJuLJ7uxAkdQv5TfY9xYlVxoPKI5BhQfpETjUN9EuinkFfOGMWV1l/yerOxQPLnjAwk
tcYE+m53EP6gClq5f7rk+jrmWM4M6yNqNUIjmv4ePDeKQGH1odZuyCMOuM1S06H4P3FhB1GTQG38
VilGuttz6z/o4xgMtiRk9I0JptsUl6UcwGdpzQueskT9/FLVMC2yO/xE3g1NbdhTzg4MtdhAOI8C
Q68+I1cqgZad94b47+ZDcoZBP61/+3aLqHiOtIZisaYjM61xpwUqJDIHgZiyrVZWf72dQsRZy3Cj
zeobXbAKpAhVKf6mTe6PABxasuf5O+qCYF9bAknxyOL8A1uCGrff6qnWjteFwoykKNc2WqGUePbQ
77Lk48P3ckOSdKT5rfA3qZfxeMPmnNbQ4CyloZIGaa78Th0K45Pp0k8cQ9IJMkk3KU0pHaFlcJvs
ktvtKfrLXbxDSQ/oIDyNkkxRy60AM56Y+x/SE+3ht6U7qomBAuxMug8P7Td0uW5FFo37ZTLlDtIK
TfMvit2J9VjRcoF97vrEvo7UpUJ+kXtPlRcWyCiskqmG8ZRKJ6SbDU8IGj904j3kwLtFiyM/FVnI
jqX3BerqK7SmTZF2C8EmmpoLZ9p8YVe1MsTQmz5YBQqff9EtzOni3fqydfny8pM7MeDTSO5mpV5F
7OY2DMaDkqZJMgJs9PliiWKbMi1E1n5V8GMozfESgxGlMj/NNGJlTf/bRzUBh9IPvTpaKrLNRlly
3+/LpQgOAe+Kk4MQhmg4znB4zNj0CurXLKBSjNZxt4LMMJQiSpoc1esIyEF247nhtitr2SiuO0lx
LhUghPE8w/AAUH4CopBbJGizEQveQgmCQOfZykctghAKyLCfS7CZc/oZYWU8/xbgTLlTZk6fTUlz
hcc5MD+DuHkQJJKdYCc4w82aExlr4QSsVgtqUVXAQjUBvz9pwN79E5+At64tT7NiSdpl8XvFpo3B
svlQhXJIzrtyQ0V9sIcdbpoWGmPkJ9qY2gi5UYvPZMEJfTUnNWyuQwHb2IL/y5b0qWz/o23tX2Iz
kwg6P0FC2Ay9mCPErAq6bL0LexY3NJjC1HG3nV8vSC3/rr2liI9wpGGHM6gZ45uDzYukaafGHG90
ctFFTlQXZ8GWuYTCIqI83sp/lD8NrpP3roAhT6HfRjNRRmUxDnVIHsv8h/EDqCUuf0Fx5NHUlSLX
DhN/80OTfRLutnmSKtSVL4NRu6CXJB6OXpyVrJD7SEfMYTBfcvTqsBfDeK0bYZi64pZfvV82/MHu
IPKV5Bp3dmhF0rFDezYovCFQzHGpGlAvAE6ad6U27GsFaflAHnKRd/URB2fyJXhHylitpeSHUZge
lq2ZeDq+CmxeqCpqbSS2ahgwkgoQXmbiSVTXHiBMZgqB8mUgNeE4GSWAbWM2u+ZwZPjn/7ckV2NN
B5X7y9oIILnDOzs1OrkI6uFyV2s8UpqDDn2WG7YhpR871B1DxVXMtwLFGIV5TIoNOiKtwoaAnCy2
s9zfoO14yvhSC/xhhCd26Dk+PPF7mIgswm3Qem7R1wYlCUrp5tDdukueG41TRvWQcUNIU42bA15m
jdeL3Wu/zRTEN0+77G4Lde22UnHSn0u+9SZbyVtI57bPZhIMe1M6je77IhoCTAnUCYgUjOznfZaE
Q9brbqpn0oxRA4joC9g0CXgqrL+JdBZap5AA2bjrtjcOYf7w4L+kul+rh4ohEiTo6mq+1RlqB2q1
Yal/GGx1+5Dv+GGAGzX02USF0JzVAlFWB2q+08Mkg+KEFPcjXDCdz1KGzamv5sSxuLmrV0T/9c1N
VHX7SxMFo9BvaOcVOXtSCL/6BLM0GIRyyu8PCgCyniBmUGKx7zNsUi3szrhr2Lc176nchod2f9nd
psNVr/U18TaOselXFkPvaMtY6I230WEftFQPo4Sk15CixCWkocyYuACKu2PFr2ZQmCMZ9TjEPXZa
kx8Bp4YXDGpy2jJi2t+rzBpbESoCsv50Pj5S7A0PsdLaHIkPVS8RGSA/mKKnJTUU6rvdTLvuroZ6
kJzYDy8fdPgBlSC68ctWMrTwEVaqcWLf12FkatwLHKxrj170OFrCB9oYTH5UVehK1/HtvvtQenBQ
OTWn328PJp5hpaSsdRBItvNSH1OunTQFyicG6nMjVQkRuHTu3irX+1WnL0MsiusyhLXJsjbuUk6f
rfC1uGjwMkHQ4lJxeDCKTbEn9uG9xDAWe92hlWSEkWAUMzsFCsKPsAVF8e1jXyOaGS3RlmL1dfEo
/5b+A5evYJN1sAMa13+3nkajv/Yo2zNkeoLnR6auRwAPlZAp8UUSmgGqhwx+iDW//e7X6oIxlWTg
oqMnne+pfig/l6YroehFarZD3Vc0E3AJ1NL/PQgwREejzqo6d5VDeiP+tzBDnokin9F0zcmviaIj
jHKbtqLbGGea0GpHl+QZAvSO5J6CzHppcyN66l1rguyBb1ycJhhKSNNbVOf8Rk8sBxbf+y5zsCco
XM3LLKkTY4lWJue3w26L2tKqx9auMrDtHWwiTz4DUPbCJLFT/olU60UxL81IPj93/fegh7ezRosW
Z1ku5TaTjraXi3zvaD8Cb18EteSYfkwJyweZ7IaCyG6G4UKIDZMNqo8r0fOTs2982NAJLPQplYwO
vwQa4Br0sBkTmUiJJZA2Xg25BCUnD2D3fEdqoLRSzhKv3zofjy3Bz4OOvj2P6uIjTt7xLk+OBbze
KC6GHwH8ZgF431KVPEMXvzUIp9xDclg6UN9mtc+zosPWiIyd2BJIE1DkgylHJz2AVhhngEKMoHNL
Mxuxgbv88kofhNOPK+MnksdEjULOuQEumCQOc+cgocShIJgA8DxTLj+6eW47lUvBH/915fxEdFa5
2XPw6ovBcKhr5xLn5hbk5LJIzNgXyQH8N4h05vELXT5NRq+zZhtrIw+9LC8reAuZneAazhkgg5ME
FJ5ppO3MKtINBcxSlpB2iE1Qc5OzG7PazGXSSDeHCzU+Srl0gxNdMNIk7LacVG6bucFPyM+uiuME
ilZnUsU4lXSlMSTcHvVuTY2rEno1hPDIyu21+K2n04e38W9Nip4+BO7wuyw8kIa9Jw0HWg1Aoik1
/J8mBBKdF+6E9WTzXRbDbjAHD6HaJQuDqcreN3u1fHqM/I5fCnUmK934hfGYhhDsAWVLr/Vg6as9
Sw3J3oazI6VV8BBRu8XSwkGogRbOtROzo0p8PCSTjWosltibZhhXUxv46BSXz59e1W//hv7j3ial
IUqBT1u2RfQGOD1l1wRJJYwH0O9qVs61a4c5EbhNcZ0fRJO0qhNcV6hRTHbhVYCp1tbB8WjyZ+8P
iH9+E358gt2jRE964QObz/Lp2IqektY7tMXojn5CGhE9vdtBiI8jrykWMiqDzk81luUEtegFPUtR
tJy2aAISzqlaCN6DSzXC8fPsNZkhVNST6eR8RVdbna099K81rGBxtV6T3DVbPWZ/QqjoCGyRS/Et
Qh9ZcNtJsDOW1qH5DYj/da4v2qySwTnXknelUOb+CXNwjGU5ivL2mg7mGL0FeArwpXpu/kAsSO+Z
qV9Jma86X8cTY2ErOm7VM+wX0sJQW+KCWBsyXgSEQ7i/AvlU3YLHy+PDtZKVPKd145uM0YTIpBm6
Ivnd6ze+fuRUkZZOQ6DAzUNc9TWgAksZME7FYFzHlCr5uKetRDy54yxkx1bQ+haQFcZHbLv6uKaA
erX/vjCyb62UiFANu0k+hbjyD8s1P9jAoIm3CdRg5Q7G6RuYfjY5DuPDfL1Aq7Oy47GbpSbmY59l
td7bzlmB+lJojghYMzw+5PtWv9x1AHx26+QUMn9fnjCIsQn95lFOOC0uwcrWmsfycA3zNok+QJaC
SFf4ADcGRGhix2j2GUq8R4FwxKR0cnm2Nq6AJv9u4yQ45C0JLCgkqbyukKclAxTMojXqWHJq20mp
C2j92DVMZpyQuTKWvPnRvWfnfFA4X8XzLKDks1A/S3Bdcrxq6Uf9cTQoSTYvdVclw18/DTi0Rcx8
OXwvPKMA11KFaSiNy7gcVOZupPhlhZve4uhOD2rHrzloc/uElY2sufxATf4qyBiIRTRm+7nMRnSA
z/+dPiZcxSriGQW5SNZTbyRSraNlVNSERoMtRhTrHqcJ55Wia8ZCG4BsfAnaRATtCeixMbUc95OX
zmMhFX2kbshZUxHWSsxzoyMpEMPkn70AF2g81U6hQm+VEhEEhdmBTF6QNqjKJZYFbH5k/4XkZ/H7
1f3sPtclr+xVd2qjrCB78Td/m+pPcOpigVCKEUPvl7+2C0LPz9XY266G1UBCFHN1+xDE0tb5jInA
mCXT1J7rZ8+wsJR9M7o41rSrZMqcXCby/RmuUpp8B5PqTK8QKO+jVpnvmdsVToob0j7yW7HlPjS0
NAQuuv4g5HClOVUg1NxCAQVxXSLv7qQi0rN1Fslv+OhNWdcNNEeZHR6W9PyjNdRKmpr4HAv2B/up
lQAgX0Fbk2lLQdjWWnc/MmWS36AVTF6gnKQw3JCi+qM57B/RvOBqd2ZhW3nPgkuR481LYy+okOD1
uVNyA9Vs3HBvmsBmEoYJp3P5UF33ebMGziaAc6nnEcSrPCnZ2o5LCr2UHJmzhw9N+FNdADvqAfM5
AR1ydjF/b7sLOwosliO69/IMBUaNNF99t27xOKEx8CLFgfVTqqb7kIJgBiJFgfn3UYLtCsPP5uwu
kcgKBRvlbTmCDHhiihHfmCmOL/KQUJ1cNDVEZ607ptzRg5qnyJgreS1w2kAwENuEHmSDRWgfFGM+
DNHVjqv4XYNUBgG2JZkxV8JFBeuiJQgbiRHcR+TUhM5ETTEnlJnlHr3qOpgDDczGRd6OTuOmfujT
RISHvbbkU5qviL3vj0qfs6v71kbWTHqpXcnFoBYXfmExTojIpFhWDM3g2pi45JI30LPAg/Hcm+eQ
mzWdL/1uXt7y/D95Aju8hxSlLcfpHDwYfVSDBXdp++dpblUSP8oapVgid/mMy8xiLJtERhTVv0Hf
KbabPwydJssJS2AqufOQr7F6QYrx41uEwdaM8U4CwQ03mhxh3Cf86aV1GsVBTbaT6qqjBUWdBCOt
xSDfQDlLHRE6ZMBeHHFrpd+Jb2IZL4qwTh8WHesA9e5NucbTLB7tJWMQvvtzMtNb4ngnid7mCrEL
3S3OZdePbYYoipkGXSatGe8LDTOC9bigbmFQaL8tN4GGb87bcX4ldP2/t2qRbcXCn9KNVNGJhCk5
8VpGs4AIAvzJoIdL1mD9hEQipL6qRh8rrYI6WSwQMl4hz8YqRXE0aB3z2tcfYZ/Fy78S0hII9+2Q
0Lxz5g3UZA2Z2vF8835sNZT7WmLZjJJSLRevGk0MXwICs4bdOwB/uLZ3ZGKduYcSXMKExuzzPxZl
BS3Mm5hn8nIvDOv/Metg/45bTqISMu5UsmMIYCYnfp7bwXo0qAeIIY0A5ZcycfmsfCv8xDA8ohgU
CAR4azSOLLJTJGwgE9UCZle/XJA+Km+AxMhEy5P/Hhr/SyrXMA1C24729ksTTkM/7GlYdsVultJd
oUAE8ZLbyY2RwgWisCUknAKaLNaT0p1/wfNmoqYnqBbPWHp2SjoKm9rw5nXWCkUXdWLEM841MyYB
wg13qVh33pUfQzWzZbHatiY81CNqy/BcArR+gmKGEShfQusMhzJQjtnQ9o/HtA9qOk2CLnAdQXde
ZCTTFt0MosoMgSlsorNtIikk7MjFqU4CxK+2RUvC++fdFrudrFZ/apE9qFOgfMb2Kv4JZKb4xBRN
0Z6TgEhy0g4iUX07JF7SNrVFBzDFsbfZ3kvQoXbHxgZw0M/q68dqELkzvpaFoalK04lvoqNF0Ngs
G4QyrAv1gzsUQEGCM/Vod+QrV89dzv6rvdpV2HGaAz2EuBO8aj/UW/+AWhnshHGp2dLE8mfX9/Xu
7o6z/Yj1Bg8f1cA4PPCG4wDiYGndXASaCuDP1081m2eQ6PKD1AHVZWFeMe7qGmmy626SlNcrWYnb
3YOk50xt3EcYIc09bNXJz7mNOyFZfSWHCaztEA9UhfMulh6cLKZM7RouhpUZ88s2cHg/nwwhEUUo
jzYDVzm5HiWbwwrXvN9FOdqmz5A2s0tEX8QBiRhg6GG8I2bP/y4mUFSQWUSTI4w4ESqw1/7RfAQY
V0TYIPz67+bDqWqqRFOKWMuCAHwOBv9wZrLgqN4BzCXotlpicRvLSz/EeGscojdNKSL2zkl0+vfR
kMhFpGJ7eWpIadhhsvU0GIyaCsP5naB1inttRkX2z+ZQeN/VgQDQnTwrUZPLpc2kmdGxnm7SsXwL
JfoGOEHTbzr2mY49vIrIX46hlZY9uQ0etc5PxTkzI+6ki4YtASBeEDivl5Z/yh0zT+7rVvzBTI+j
ZsxHbVhcC9ztwWgJt3HSW7M+0ZZfm1pBD0/pYUA8Cwf6tNBuAoJRUC1G7tzkQz40u6PMVoxlsgfF
rY7VBT7RtAupFh5K4mC9tj1XPOfZiseWqoD80DN0yxwOq7q0xf9pro7HuwsJGBE4Xjdb6dnuVW3P
uh8jpigzgL49oA/64kB9szQZROhwoWWiiHI6lUVPy8KnTykS1oSF8foySdGekKJ/1e7eYEPIMId0
NOZqZyXBhhVpoedugvy1HOfTN3Vc+vivXk30OcPBpoKHLFGw8f2d+eCcjmMgWfPOrJ9uyhd5HMBs
DPSVgsYwr7X2bD8RjIt97uEUswmnn5omwdBUB9hhYmBOnYBJRX2+YYyqK8VlfDFMxyua0tfs4WzB
5FClyrUtFkd2tw3dSs6OvpC5gj03yhqWVBzq2D5Q/V7R6sgmrZeohmkWxzyuc3y4WSRsm001zMeb
QLaDJKYn1dC30L8Pgkjw2pshCW8i5FoLMMRDm6EhbDcHw+LdaXzaItBO6WHjDPWuOrdguxut9mvL
3/OJVfmCmerOvuHw2ru9xGzm8RyfACwf4tDrmzUVa35dhV+nWYYAtgVB/e4XH33ySdv+9iaa4lLZ
ZVr6cWqV9REPBo0yKGVOI1NC4XSxlYKqiERHzkyEFX0wJteHMJd+eZMm0YqaawcGdYQ/61aHFDTi
oGIK2J1l8g4x2hmP+JrLisUU/Yd2d+k/ZI+N+EXwGNUjdVaVyaSgVKCESUIjf4mjWl49enqW1MVp
GUEG9W/Hm8IcNtCqMZ4ctjdZUSNQsSLJadEYmHOOcmGTC87Cqt7mhnWgPk3u5XYihLcgFr96oN6n
HvWg+QxCl2n59UzIYbT/WIuwLJzVjnMtokv2Eb4xT07Fdp8GSrwU1OoCZQkGg1bcnsHiTUGufMS4
RJdMWnQH5ppfz4FiGmA4TYHXGqXea4/d7otakoVc4oIq/JkhtLfMmSkGUzpBzPIoV7cYMITweBgQ
++77NPqs9qgfqXJrv4GkcZAeME8SZ5XRxxh4YZBr5fTGkIcgMcM3ZohPBW/8UKJqeWa9HIsOZedN
Fd7JyxleoH7HWT12YkP2nOZuz4T7C9y76gaJ+tXUyFs8psPVq4fmBRultt5wrNjRC7Ym6ERacDP+
P76IAEOtiskV5ZldpIwmKEO5nr8kuK0QxBtWfomA+IiSrUGf/vO8A2jB5+aewqw/1jD7Gaq6gA7Q
jiV/pUBuwTb3tC1TcOMm2+kaBViIGZZJy/jIgZVh3dZRS8trciWf9KSHaLEa+TBexsiQ+H84KI5o
yZaKkL2gJAQeax6TbfDMIlfRqJ64/2u7K7khFUEzEPAC3hOAOJWtY8eIrKc7RVONFA1acnRWRLOS
cYQhh6JgGESVskrMtv9I6fcm2LS00q/Mmo7+JWLK+mVT5A2is2MzoqBsPalsSZ8PTzhRGLHdwpbv
BJCN6GW6QJ0uA+Vtpv9v+x4Zxw1sp567KOdlacKzUKCwupFqIsz4CPHoHecw3239COBEwuKvXQ8d
NQ64lLSP7AC7jHt04t0MiGDRG5p5o86UGQoIABl+BymBRslcnIkCy8Fx+39CLG215VUlwQ4CG6ha
lBjQdHTAI2XOEtPb4ds3fPfpEN4+pLLpOPqkNGq1ZdYiGL74ek58mFc0c+MNF+XRlcKkkIQtPjuj
H7M8vggylL5jk7TDzTnKSbUtFI9abJLzhNOQAxlqnsogQW5jlvf8tysdWe88+TfJy8Ah2d07Njdl
tDPS0SfLo6yDLl2PbIcQ1QBvz5N4n2yrTnl5OerJtwBbbXOe2v+wWdf7eYM3rdT3p3cB8Uv1u+GA
trX3SOFbZ+6k8Cote8oJDyqBF0nU25YoJGTeKHytGoh9en57P0sXTbtDAAa519zDJWXVjUYNnLCG
m04QuJx0msm9FAUGHsbseq9NJMq7Y5htX6vJWHbEf44Pc73bDmW/8dPWAR7iHqD/ZyKIqxWIwxaE
V9Cs1PbRtr+GGc8ta2x3vy+8Jjj4vkqwa/1JMI+azvkefE6AmDgPzcA+qkEa6/7IAOer0dz/q0aK
gtkbl7uA/1iMdI1ugAji3BhSo8XI+qXA27O0rf1is0WWM74KgAzGMLxNIoDri+sCS+5KDPBPd3U/
l0pyfxgMwduDJCksdut99onkD0Tyi9JHNQalAFP7uAGLPTwkrRrU/u+nxy67s/HFC/qZ0vFO3gJn
JJ4Z4oIVaf9800pYL511OzK/o3jDMHBgOmDVXGzlcuci6jhO2FTgn1XZvGXSaoqG4eopuYW5sZ5v
HO23x6XmDTqtDHd8jNHYMZH+ur7LS1BnfSUwE1zhs1Va9GQk4tIzfI6ASGkisP2+SHMhkaatguqz
kiLLoZfgLrt2p2EuzVrmuJnhohWjfJqTmYVlm5TKnqeSlEPYKPPkL/m/L626Zg+jXH5966SnWtRb
7RMP2un/ZQos8zg6JG0VNsu2vm8fNBpN8DrJy4pgzH5uOJAVNcDKMRaztP39jdJmzDfum5MsohE5
sYhYTGOZNIB/qMcBjJP9rBlHY+imdBrcUjADNPVjk4242edkrI0PWIg55L1DXlv3iV2fyQLFDcSM
1lspe07kmYEMi3yFvIJC6RiJ5K4JemTCpV2RZzRrLqAKw0cmi8H1v+h4mklQtc5cyPhq3u/QBzQm
FAQXflIr6jHxiudH78khYlpp0aQHF4xz0Q4txM9cJLRUHuYv8Ym+Bmc+2ybd52aQBHxav6QLmUK6
EhaBqF0EBhQDHEL/X99M0kpPy/eKZOyqgTqUrQP5ETqnzdloM4TRM0nKN/T0mMxGAKvB7sz2bjID
CviAzllJgl9g89ZFoZAyB73RgoRXSeHbDTaxcT4UUL5xnWVr3VjXLr4DS5bX8BoiUbZgfaiajMFK
ER4+9Pqt9yzD7Zgr/ebCr3psMsuWh5Qua3emCXRzvrvT+CxJfg+QJY5y7FFPwW/c404oLqG42B6M
RmVRgKpMUU1UgY4NauYFO+1M/A88DtpCWZstS9fE0cJdWdOb+cdHS+uu+CrFO4pnlM3N6UT3z45n
FsF+N7kllOP4NdNcM+HCqamxieHLK4FXPNsKQb0V2dy2gI2VdkRo5OJ2711/BDUIPCyToKMil9GM
sIHWeFZfL1SVZEtdnrfNS5DUsORIpz+7MhKshLJ8nqasoYmObtai+Wws2FKlgIJD0eQjzGvPBca+
Zy2SNYtgdFl1HaETsAXxYsHcdcRlMVM9GPV5bNP7K9DZNoqe3GCJZb/OVtHZKZ7KBmJI4zDpabfi
AbfXG7cXAhZYY4ctR8sJzEnr6zDi2CuPTzRwVp8WLJjxC0gdKMmZxLigVVqcS2CsSHeykah/Hao9
tJo4HcHnlcMt1aJDAhUfh6cZxdhFDqI+kX2Oh67bjci2YhpzkcCrtbFDIcAvMJ6AC4mzs5LKoet3
Rp6TIwcZgnK9NzDctBFg0P4e3lC5Y8bTG7SGskvLvRSuf9LeV/Od+lJTZ5wKIxeg2hfJtF/KRNJf
6vgM3h+N1oSyktJs29yWkU2N09JTh5HkP/ga7DmjP/r7USIXyjURq9jz/BG6z0Hvm289c94yE7dg
+nJHBfKBDa8eSNF0BxBKZ6SoG5tkXq8oZ9orzkNIAR83DISv2eUzfKbbWk0vO9/4HeyPcNuriE6N
tk9lI67W6rOVVvODBl5BIrbk1pO392n7JyVYE32RiXVnLpiwlrIZeoyo6LLipE/Xdn/sf4GJoYzd
f7GxpwRwm2PQP6m0CfXnR17kWQMYaf1bjLnWMtibq2mPK2FqbU7gJdgXNeFaWN4brSRV//MphZQ/
NnKS/0NYbvPhXffUFPeP6WMdjeumu70IRemnSXTKD8po3eD797Zdboyx0dVdMcPMZue2fAqnQMR0
dBrfsoCzHDI+lhZrr+D0RK0hveHiW33Gpx3CLxrEQBn/NdcTAtdwGoefQ0jU7+MuLuYnSZMihqla
Q5qUK7ESrsjuIGmuuoU32cF1E16BqF5ICeTc2d0i8AdndhpsjeQ4Z5/Vd84Tld3VIdw6MFcE3+Sb
1D7BHKLY1j0jJIq2WDxcpZQavqhS3k80WNK9INoJbcOHyZal59/XYVTItt2EEJi+rgf/RJWv5JDd
Jv3tA2Np4CG5db0N+0etKvdzZ/6mKe3/CqRVBrygNiNfzzjV4ZRNbeDYACJMOp2rMlHnH09D6pfc
5nh0U1jo5YQXLypl3E0jy7Rh+b78IzB+G1QWZpyiXTPjVDpziTuFghB6coMKjz/dMiI58TTW3vTl
tvk+dEDN0g3KqpvLmosaVhBUClooWm3E5xq8Jr7eRSz3i3VJ7tvTfQRjzTBUstC7MznRlyiZOsOB
Vc9A5BFNL7AQbj74YrsgGRvbDhCZglLoCrkO434lqKEmtf8psYsJX0kCnDObyEunHbzgW2Ibj1fW
ZlKQn+s0g53dzHyZMNP4ZqHPsRsUk4TT/KFOuWl0mDrAbcTdjY1bhf6hljnSXna7mzJ+K5QdKkSf
u344As1puSYLwNKuF+lQfTOuSxgg0GGExcSST+ugafpL2FcHKYodNkpjB2Rb0ykWHrv4JJEUrS9v
oNzVWz4UBbdapP31HlhVhHFXFYYy9tZmRqg2hzRXDZnAiQ91rMS6AaGI07a2+0WHlohqv7Jk2wq/
BBjhG3Wz+NzgCzv2BJEwk1qNRx7JZpH5bEZ4pSsiMUhufiBSnbd1hQKnAMDjKDs90Ww9BK9lDxSJ
uzYSM/xpC6b+abq5xQEN1roW6IAKhVCND8fUblBsc12kQIlx4HHe4X1Wu1xeA7SsEJOt99IO56yA
E+oaRF6aPQQmuVadP7Q/V2bUNSHt2V9Z4Rh6awg1euqpHTXSkU2tFKQKz1z9XzOP5a1Ahiv1uIB2
LYzbIaT6KfjOrN+NFVpx2F2+LLIQXGx89x0TlUXLrl/GQH+CICZnaOfEHfbN4xL6ZccsZ12giuRB
ycsqn8DIJBpVkN2dmMUAJeY3vhacLExDxHoOLBTYYI/c3gmbT7DVn7wJxHJ29RwkBWSZ5ldFlzfs
rjAJvrQxV5P6wZxk0vxjatfvH1fnH5R7RO1gOM//YOG3/mVCzAc+iu4l+uWLtmwjKAU5Svmc/H7r
S0oYWGXq5RJxf3u2DqVZqIG8O7j6KO1H030dnlSECURjjnnh746lsCq8cG9n307ZUUn2J/vw9ZsH
/A1rEcQ1AFyIObFBd5JHrmYucSG9zUckqLifuRwBtkR1pCdibT/9bmUVCbUi6iZXYMdK4IniaZWe
62u9ragE1R3U6s82GmBHjKUS8wRN6Mxv+2BnX5YBe1Uz3L/edU6Jn6KNIj6tcgagM4a91y0ww5Lj
AQMDzcB4uvNL+Coyk/qR09gHOxncnk3NnMlz0CCo74oMSezVf3PkBjs20xkmnoUWzJMPmL0zVsCP
4g3R29NXPvAY8qoNMfq4v8LxugfbC6vmufFMHmwZK/w0Vfk8jaYFzJ/3G/jVyuyZaIb1jEoRmVhH
zS+Gv2VCH+ba9Yl9qp0WqgSGke6nM51o/Jnsg6JeU14W3vlOJ2W+IjzISO77znoY6W4AIQDGBzRw
M5mYiqZgrfZj+QZIGSmMGn8fAZHEmiGvuDW7NP+0MaM0IxanC9m5UFF+TAXbREleiPjZvk5i0qS6
lcZoKfERkBdt3gk0ra5kRDguj+OX5c77hbJmDoLOX09PKUhzI6AM6p0tijTjjBor5LEc9wZkZAuc
KE+BPpsa+MxSKwZgbLzcIAbBsDPkJcc8CATUCYuS1cFgJcYCDo2HHEhG3iVDapRPNr7g8nDhg3JC
FQ2GQjlGstSbwhegxybu0QjKCuGo5LSzgUc5er5R20eAOR60o9EBewcfZhQdIe9RzUtIiZ8Gdl4C
UfxPwDntjw8GzxNFt2V1eYQmx4FLCijoDe7PjvacFfkhCPgLFc0F/nT9LOpImsC9lnwGApUP5M11
BQXFzAnj5kZRSTkuXIfhMwj0w8N+XrnneTkniWndnyjUFrteG6EpvW+EhINQyozvY8Ht+cgNbZBU
8d6bFVVjNCjUNBS/AzqLukmG7YB+TEUdJlHRarQhULfPR6E6SM4PjpRCU9hMJuz/WB/e1l8q+jW3
WHZwMzLH4zoDTQAuvBs5L+YK59R9/KnZp+Jhsra0bh0p7SUdjgU46MG/rHO8No+C6kRitQO05CZV
wLVfjqwp88s6MC13WJ9gsZiQe7UOa4CFI6CWAWvPu/NXyECSNPyaZYs61AT8MnF1XOKp3u4NifFe
W1joQgM8WNyxKe7ZgDFDm8U8NvB9MFFtQNPeerkxyEn7N2CjGB4FTIgvwrxRW8aO5/Oq7sHatmYg
y1WX8lgAEIGQKhwgNhqVdbG79D1EPWgOnN+qEz1PuCoYIwZyv1zNK5Q+xVyRi3b5kd/PJQefPYrS
7Mq3FTKQd8FOEM5wvbdM9DjYWzPd6cWokpV2LCREOd5S1Wo0efyleItnRDmPBCh+wb8QvR4iLL+D
cAsTfQ8/644R7cLXXb/B91aDwegGbS930ZANJM7lxCkjF7Zm0uA43i7CItaMdVU8ciU4RV9N1ps5
URyZXircGRfcUerxmyC7YZZCugoa4J52OMEYq8n3LEIa4ETlGy8JcbtORUHxSyEWDZurLPffKpma
UgU4Q4JFN4+6y1t+EoxyvLkK2QFg5Wj/T/E30eLAF1Cw+JIrQ3wm/111FcU+gf5nKM/A7ohE3zLi
19pVpeAIgkLyvbC8+fST82cd1C+fkdWmk6WMcYce0+ECwoi9AbYbQmqgEkfxyAj8fm2QY7fgq6ox
vyoGxR0dR3B2WRugy5xIh2pztMs+H6SMoXbSpDPerPQvZb1mxN+Ch5TKZPWtIRsj5m9ZTmrI1rYg
1Z+UgGEa/lOiy24T1ZBoKZUwzthUgJeJ5RqbPd2CB3w2Js1DK02lt5VarsNuM5yPcrL+gy6O81o3
tJto3ZEeGDD5qxukdEXxTJUUMDkt1QOJvgDYRrt49W7/KwiEuoPxe+Yy6LMbe6gAAZLRg229vlKQ
5xE4u9SB456e22UrlL4v9IuhMZH2MoBLnHVojX+bztyhz34BZsM9QQ9Q6Tm2IEodvGe5HF4wIklg
7fre9bwXd0XluGSSKNU3dovFVKYMfKETc20wsAcL/dHQgHtDugmjqMQGOakOiXCLyU2xg7cagfxo
5q2WmMfYLD0hIoJHICNuoPTAHetfPytvSQjchv+swvpHGUIyuYIUB5N9uAiQr7yr9LrkKfHhkq1q
qSrCfLCrNhtiztCYviYrnW4Pjeqct/nQKzM7an2w54omx88MU5RyOMOQ0L4xw8+C78T1TJ7sop3V
UpJEVxMueZ2BatG37swZIOsgOCboWKxYH30RwgX5haEqbFLeWHyQR1Nhy5jarq4Kyeu721OqC9n3
NfcYDAu6cfCxy/FuRdCw0Oe80L0qLAANfi0aG+HZunDI9FDxegX60EgJpzIyRWKotZ/6UTDRGnqz
vY2iz3wRTqkr2tz5z4jCPnZmeTXNN3QL7Og42EwC3SOWs/yf8DBeWW2ldpqQQRO/iYfsADOmoqIm
mYyxotsHYsTB6SsYgdTUbUrsLfR2zN1BM6bsO8qyXPfRfZadIUSFSktK6w6CWUxwppS6dPKYykMQ
yLO6ISttI61v3jwoFi+aJGyFghWpr+eiCgPpmzY/1SYJUsBUC0stmGEmX+cv5KjyAHQCIiyEueYM
5S1RtWe8WHpNnL5gcQPTccSTlaFNGeDNyCjmuwyfKG2Ie5CQ1X1/tn+pPi7OZO+HnsczM9j8dBXf
B/2wCzMOE93kx3P6JdThf31uSt6v2EVozmlOpYtpHQaZLHggipyGZUaxkhB6tgvszGdPLN0jB6Kt
I8v9WPH2n2HHyhtnLiMJXCG6KmZih4XEhc+px5UulaMSUUmSv4YNduVystvkPoJQA8Jis4vWBC5G
jirqg15n3+CvQ2XtcA/ortAhyQWKpL6Y2VSWQlQWRc3NR6p0rBAkQmymKO8lAuhxGhLKlCksC8w6
x5xzQVRHWIBLd2L7u1Ju9f+/6yVZ/Cd9pH2P77IUodEbZe5gKyva8x8AxIEeuIPZ5B0g5RcEIWRu
zfr/I922ZBiIiXuV7ndCFEoN84maqTvtqdF6y/ZYkDYke3tvMU2rZ84IUYbglweURV0kzelzDkM1
a2LyXo8hOEWiI4yOM4wCkf3hmHm9aBZdbjw0Cg+any148HcBbHtIGL6HBxeu35kDWcfJGwJsPfA+
B1x1N/LcY2UhtcOvsxcXyfwfLKOw0wYS8aUeX2+pGkvJpPxCsb4sWEgNoF/ZQ7oB3Pp1pvqC6Con
bIY1hGp5nlBj9DuO63Zkv0q3tXJXGjpghhHPhWlRe27FawJqOkr2E8VgxK6aZxVr8VJ8eN2rJaW1
0pVy7ryJxWyTSkRKuG35uHDtjWFWJGbMTku+VU/vxNXOOGJSRwDZ8BBm1TIqXr+laoefg8pXuQJf
dXjDGOPiKY8tGCvMUwbgwp875p8npbA43QEixEFd90pLidseClC86Xckt4ADNQWRrgBiahSQ/R+Y
rZiSp+LreDvmNQ0MUS3cAaXuOJXgPpWhANo49e3MC/QsPoaawjb5J329jgw+7DaQ2zajzRTRgacP
dIyjVoXvtua+POOaLtmrC+chSuXIA/wUfGGlzYM/Kf+Jr95xDEpfOIHaEWDvwY+HYfvHE9ju+ESh
LYzVhpGEjMHRuEgz1JC9qJDjt1nSERjcfjwGagwsKPbtGM9fwVrAKmxOawivPW+jSkOzy+8G6+mV
z5/ddx+Qw/0AiKqKFz8NwQLPT/LkTbOVp9ivrvlpX+uknMXe5F1B/4dftV0DBxcEVxZZEWr5RTYp
tUcPCmt+1p45bJwL5y/XFOSNMiUI3dpbfPEb2lgRUeHMScbQTZejcYzNTYHtcXb2cBq/tcAfOzgo
tZxpfFQ5c92mK1NCKGVyI3nzhb0DfEIIaeli3J1winIWVaa86Gu/hH12Qahj1/rhbrvSPU6y/ZZU
sUGHuswREZpF3zqxMclyiK9TKQY+oo34/atnHqHnNEBgnd5/Nm0Gtl5NozbV50YqbBKGfkaf8WJW
+4EMZeH6qbFIv07Uo0ygOKrBM7S6eMXq6y1SRC53OBuYkaT5xlc57DNCZ7fwoGYuHYJgY7pHNKTP
m17xNRu42vB3HUH27MJkyAtoGO7+b/aE9qbVhXYH9cop5Haj4bsENIHGKOLsiMdspyME2pfQEap4
+JErXWdK/ue7nKr+iFBXTwiNyEl/Cu6SCHIF1x3TwLtUy3b4vF8Epmm18vlKxyBgP2rKL77BG54d
ON1+bv/RiFPGHauF30JuWNY39QjzAjP7e2/E57vo4i+5//qdSjxMmjBYtgXorExktw3qchSTmlSV
kpLQIcRxHKhIthOq3OCphABCwf08l1ZoJ3xjB0x3WcsTVnja60OCkXxP2ufMeKJq/bWDfRzUDXz0
7Y/4RpkyIoK1oNo7gUcBDtwAohve5nPMKtJxoNgvLg0wtooly95MNazIoO1ALx4zkn3JuMwvRsUZ
LGOVWCyFBosxdIxGDP7iViWqjph8vtMfgSPkDxAYfnadYvURWbitTAUszDuFKJgbtPN1bAcmpTAJ
1FCr86oRiTTlxdNrrZ5ImpLyR2nXNHTcrtidl+8aB/av9StbTVVaDiWBwJXoV7v6MyUaE4LFhusW
LJ79vc1DtbmhERLl/gVxSa/rlrP5hL38iLBtJOc/90tVf6Pplekv28c03xKT+74T2KNipuSLvau1
ITXbStab9rV9zQbGyRnoYptczZKMECpk/fMGC2shlbInEzQLhE3c0orebTrhBKoG9KcGnZaAtw2C
iUvMa9qRwOlsVhJXcexNGQVgZroYTvb8a58OcD4s7A4RFpp3hH2v5dof2vehbaNAdkecA3OAIpVk
RaqbvCweH64hffLcR/iUFuWesdHPj03Pjih4j/w2vCEsM8cQT/3FFWntIErIHUGEsvKNW2AJ6jp5
UnRciLnuZtLy6W2nawNGssd6SwaCJbucGrRZ7w3Vr5a2rxnXlb0WnwVo9LP6ItaECxvp2azQh2RN
B3OtCZnJorA4wdSPZNJCg8i8Gbn0r88qCDjd6Dbl8jkXJImhjtaGDB6EnFc2sdo5f9UWsxQP6q4L
A9Pnkq2GFMeLOoWMpfsDk1YEVeLNErPxhi3sn8jYs/bq4CHcPkqhrgG1zqtGWs982nj6+6SCGWjB
EtqUDnWsaSO9gzxJEhmFjaReheGxuSpQfEq5MEEu6aSGBb4LSDAa9RM+5qVEDFNjYQR2hUeo84DB
nLGXnt0gIFn5MZTBUdRA2MC3tiCYfuAfrF5CjIycD2e97v5KPgIaxt3yYAFITPoe1ubMC7/VPSMA
KWd+AO79oiYZz9A3uav9VXResnuVDmdXvJzvdDXkvGAUU3+gWD5pKAfD5clNsWWFMK8dWATsyID4
PUFO8unb1TIp29W7yyDK0Us93qs9y91uANKl06GCZmx6Cs5lz/uQfU7tbXVdTkh0F0PyQgyiKhDi
Unb3k/FyUqfNv+3XkNPN/BB/WML6jQJPzp5YQxOqnsGzXxvMGdyLFL4nBfsf/aWYHVOckozPkg24
frlhewM2stAZPUBVZtj6C4cTwEGlJcNXOUWfzvxwzU3mWDEUuYWSVOaCw4ruGdoWAJPTUjuL62fc
iLUu6ShJAgHGON0I4ThJOyDMh77BUN+l02GCGGR3/Yan/nZHCAydnpVASlZpQyl+xVIvJPnlogfP
sDRQeOFqqLoWPaex5TZ1CtYtZstjnSaEvHcyIdrgzpttyrvHxigrHj8IFgvxW2WOSB5F8SS5CoTE
uGPJWUmsvp9LnebwhKv1PLC9IZJEbX5UFuNxdJNEG2GsFBlF+Dl586d5E6nWkQv5M+PRP/7N/hBY
3hpDKq75LsbdlwlUkQj20M7pzha8I4DAZ9VMIm3naxowP+a8KTjFGz1RpwK9oL4EohKsN1a/ouvG
/cp9F2NhLHDY3j/QJ/+t+3VNswqUalkMcHBCH/+j+zTMhCDUkk6/dNfOmyopIcLZbY9X9QuvnAg4
yzObtobZrvj+Mx32PRidP2oqNrnMcAIV8h9wJgDLNHmBufZjmBIqfBjd58TKLM5agYdy5iFk7Hwq
YsgTU2LipRtQGDIK5heuZq+GOoNlIGpr0BO8WolUNUNA21/Y29dumzHnbjxLwrS5NjUbiv8rGaBN
tfESjOrDXfviPz0c10CsDNraCOaAFcO00R0Tri1V0tZWqmF4Zjvzeg+RMg9sQ71GSc/UtG3LQAFT
nSviAkE1POMgkofgKXZS1qsiCYLti4jN5aVG200U9ZOSCX/OhDyD2WC3P144PBtZluxyS/N9SWyU
8i1yjSQ6GeyLnJFF0tq7ijol1W+GcOADvtSnXMxLyqpprSBMx8Aaey5Xp9x4ZQn8pfGlysATSRkb
cNF7KvqIk98wM1YayfqIB3Vz/2fxS5XC1+sVr5EePramCywdEgEkxelng/ap+3/NDeBqeQLwnzjE
uts/RXM3sVzBNX5di41J/u1QASQCfnRL3oXjYOJcOgJhhvuY7RvqoBU2xleWWtqbeeimzO2q9M36
xf0giLpNvjUiOslBkQSmbbWGi68E8PgmmD0lNA6J+lgajhQ1OD4kKMojH0XexobnbdEu2uDao/4M
RWOoMq9JIranXBQzB4iVjpfrtLzk2E7RkVh5pT1BlYU58dyv5ZngNl2P/2TPrxJAEN3OlvNwoZZc
ZampaQKW0Q78PjW5qmLoyYbFJdJKbcLKBXT65lxGVudrNJGY8kFImqaALNcjKd6M8V3ea0DgErDg
w9vgnMb9YuC/VYBRprgOsuY0L0JerzichIB0QMD/m9ny0b/KRfXFiPaGlH8SpEcPiw8y9a9KcvQo
3B1JJ7anFSHgqbfJaikmK1aQJ99yDh5Z0v6ufEjb6BNQ/QH6FY0cQcJqBqalSqcOFRdhXLyc3QqK
YCrQeZ5QE+hj6wOzVJXnIEYp7jHtUE/VZY/rQiUl6YT77m/uPdgnwdJjGkpKXnWOle9hVth/qGe7
9TkoqfibOBMaNsI5xFZDmjZ0lGwCNiw9tq6EJE7vK6kmSErDMp5jZ0M+t+nHkuYGWoojLi7t6hEB
yeGnzlHffWmkkCkP4aSmmyPh5seGsRW9lYpFbMl07BMHUHj1MG+6FZQZbK8Lsfunm0lymR5zewjr
zBlQjU8hdF5xs1XUggZanXOb683D0WfjeOoggiE0f1Ks2sX+sHz/Zcxzr5GT8yOTLYpFBqIzHMzM
oZzKbyba9BWX8A7xOo5MFG1I64va/t4sUooeayN5dHku3iMiPAXiqp2Y4fb1qO3t1AZ0vwcvNwFx
B4YaGTPvCrtkojg+pnO7eypXikVNxbbNFl6F+ZOmDBpYH43IIuvbdBgC2L/62MxaGao1oUGdmHOb
CSpJCZ5sfmVsEvm6SpRWD1SgY8+4XkfV1cfXCaSTcIN3nZT5iupK0c9/sEnDWEBdX8A9HXdHOkW7
Aw7yIFcoRTSaAFY4G2VyIrX1lwGK4gckDTgtOXGw2X64DW4IfenUCusUH9bzZaQFz7L3hqunyXwD
RMsr/Nud9+k110Gxfbcu5g71ePUPfG6Qlez9SmNBg5Dj50iMV4iST07MG0PsHlwva1VRwziS7Nv6
caAWEVDfzA5xjHPUWxTtgnYHwX3VQzbzyuckQOh8LspzE64nZznqvZq/08+5jCv1ndsKe05NP5+e
1CYCGz8Ulvj3icjGqIO3i5DEAtNOhMtyjPPh2gs/EP/MlV7+/BjMUGKHARS5e5YZJabfgyrpxqqb
ubokIO4NilKG3sbWW1oAxrWiMEqcm0S3Rtgn+r3nNOaMCcwNtoOdxfFb6GVom5mmdDu9v8LMh2UQ
X492ovOSGRUNwPXALlQcL/+vmsUlIuWc3Tz99cA6faU/BGu897ihusMJHi519dlntX8OcWIfNP20
UVMwphODlIKrrqae1I/9DoKc79xzhMjhHEpCte1si1xp/6GWqFs4sCLagwZQBa62KyhauJsaicwu
00W229uhTS8bRUgw6PYAO2FDfO2pqO7bihP0iR/6DsnULgznipx2IDbNID+jHSB2l17KdNYNlxHg
BTf8s9MZOS3bFjIuTrTy72dp/Gydsserg8eghncVpILWkBd5yspv79/H1tdY8jre/vzdYs+0qtjS
gopL9KJB4BesyUBAr38ZCkHrb1ZMYW9cPbpoIrICn2BgCaObtyhmsjyQ9PYE1UZLmCoKG4gR7or1
kO8mdobJnPGrrSk0JPE/CFCr66zpCfYjACRioj+Nab/1Ebqd6IxBfr/K1t3d4JLvgNBZg5yfjqUv
M73X8zRE+Olx9NxyCoDkA29uC91ApV56iJ1N07ljx0JZkO/4q7s65NmrZKhVvJGIiCXFotyWF7Mc
RUPTFFfIWcVjeWNnB214R5NWFtX8QX+BuSq428CUVqiJkEIHUUeQ/LD5iMaRA5xGesmnqysY+O0H
RomG8LTbWYGWLQsMgFYhct3XD5fF4oXxflEy2K47H6LRQa77OW8NFx07fImqFWRWmtW0zZgjkzsY
INoBBpbVmP+10diLbhZnbPxTaWJlpIVK4kOTiIpYJmTpg41oE1e09rwDy9F1Q+5huBJCzGwzdWpf
SXal7MRqPpOUuXGh5DCV+vsViImTyPIxTjIIlE4DdVthJ+MIKRndTkIpk6N0WmMFEFE/xlAJwhdk
q5P0/sIA/s5tKS8zIt+AkehpblMf1ofCBnxFz/gZ8E049DZ7Py69HvEFX2tK06aya15z/6gSbFos
aB12728yD/24sncAP/NVDZmm5iKzC12iTxq5uS68yXZ8oHWoO+jnI1+vwlr7PjVBukra107rcH/B
HrgiDemSMLgV6CFjvnZ6hZNjeSwVgEdWaA+b/XmoaRMGeDfklF9fvSg428BlJHx/x4ErTnD4XEW0
SJZ9NKXe9gSfYl4Y0oWRu7zcqvjho7EF85HRpbAWhN8Bj1OnFJuvt4iuo6zKP6PWuC2wCs3wnN63
F5G8QlFLNWJ06u4hn+xBPEh+wBkf/vWkeEPNqhRyT6r2Tw07rHROH8XBhc3vN7E5AHncFaoLzU4w
qXRmhUq2Xy7y4VPdeyZ9sI1whnXjfwQPq5hGGBP/IldzOCfePKoJJQnGWy+PCwehrZHMYDKUTV6+
wT6Hw41az/QI1RCRVxWebYFj2azu+MbpqcoMPNXDSoLUyr06E9MK6Z4cpl8GKylensvQhHZ++CW0
0Ri3U7Yeyyh4v4n1ExaQGe+u0lBCU+pd6IfeIZgXUcTU3XgKJYBfn48B994BFL88w3x8QQPUQs7W
TFPhdSZN47XuBZ2Sc16XS2lJmlIJnTvntsqLMXLaWZj2pDUdVN2Rbkky86I2LMrUWw4/LmA+ViDR
o/Qvz/EqbFaYhbXtdsXlYLxb3ehkITqz3GDOAFbYVDAE9XQV0kSz+2Kym1ICd6qab5gSGklQX1js
eHi4CXnoLglWakUTocK2eCTWsaabMnuKB3ALUPNYzupX1HcEnvZgLH+SHJi21bop/CBxiuXQHkAc
N6mqWT9ePO6QxfDFc1EgsZFoaksfErEfpACqdefA/ycJ6XaRJXNHAJt2H0mP176bw4wpgfJQDitQ
UkN0xhIBP193+z56tjyKoJ58yTjyz6YAhFE9GqYMjqP1puOsFjGlh8+D22ZImK4Vrzy9fwqwX10b
0rNnoI+DhmULELihmaSqh3Gppg4naUi8XkLJHOk5xHRS+tN+F67bvnYXzugmcpaMTeDVID+PKI+N
RRhdzOqHUlgK+gysEth1ZRsWM2D3HL9MPdXrzwmDblPhJkaBZAzPVNuQS+afwvpPhDr8DU38dtVg
Nd3x98TPqViEYO7shUrFFCOdGMqqnpAjj3XRuUUEOcZLd4Kb13BmBiWktOEjo1tc+915rfN/S0dc
ojAZ5AzdyLi6nVkYZjHkirt0C8XamIJbroRbHtUkOwtjwvj6+vcaaDXflge6kIUY+RmvxDQH2TQQ
NWcN660Hpa5NScLViFVR6ESyK0mHAhc6ffCk3mwFHpZr8Lh+2rf3Dju4LBzDwJfhmsu77UF4DRC8
yBZS0LofnQJlzhbZP06/V3h5PYie+cjFP+EyVCBI2x6V7/G7PCbkWVFnz4+OmG6f3Dkk77eonowv
cDPEl+yqpTiiIZqQcD0gbnGH04UaHRL/EL21Mf03ZS80tIFK/IHtORN8xwzcMe7yJIRPSsZLPiXr
kBYEqafzu1JirHys292Qg9e/uXpJefhKeXk/GxEry8xJUWFTjUaJmHiKIg8BxebEdLv3H68w1oqN
Hcsd/NjdRkGqQx3/meBYVfh/DjjjAL0ybIYoZT5peqZJByKqwIAAos/zrN5CbEx/Y+dKeHqB8Dzj
AHv4rcYDoL+EYaVCrtMwpbNepknywzFFBavZ/G56QYVwF7qw1bfKCatMc12oIC7Rt0OEHCw9JR+D
7L0jMfRnu+BFlXSUC38THu9v92PWIEgzHqg9i2qhzAc3LRmso95emROlcUi2xRUil4nu2QiRVgUI
s8B8eqbRCGuh9mi7kewYmNcJrk7EPbxx0QLeC0230zhHgQDY2H1Sz/eiEquSyM/vBL8oUZ51SgSR
hcOe7rWKgJIEyx6wunn/zML6SPTxR/HIqPPviVFXePc2pom7gojhW+wcrF8SUf7wv1lLuWDyCggs
m2UD2FzG4pvHplPPo7s2DqtZpvqAFw3a1FxXKjuAfGGg/5O4gy+7dtpft2ESHcU8HtJ7uhNs+DYQ
oTEVkY+W5q0I9mAmGPLkOv1jrUH3KfxR10JAsUqzdpHy7B4xMGglei/KUJDCvWLpJ/HsjETRWxto
ZQ3aYqVQ+AwS2ktfzJ1wBip8bbemR8fRQ9TSa9qzzg4u7Z8wdLIqQlZ9OmiZV//NL4INlOUNpw7H
BkhBVL9RCiOKmL6fYVY09dDrYqZEd0+63qJeal6uU6VDxyG56OmiJksT4Va27OYCWdP6G6OF2/kF
HmSFWI05UUi7NQBvMeVsUyR8Wq2w94V+QoFNxCCFwZd197k9k0wcZxod7QNx/7p2Q1fH9ygEJcWx
4ydonycelBUbsw0pdBWdsjWGwkIZCdE5KqWkASIg0DqhuTzQCqNejRawfx8VYPDsLXcAY12svVIT
C7l93q4zsTAU+Hdz4txhFpM+j9AsJUMcCPTuhTVRvzal/2ldSrnfN3lfk6LKiO2DPzOeUNKhEE7S
vODXNlRZOMmZmjMseeACDPHrz40YnpmHR8+RTQ6Ol4yGrD4URYvqNE7/oY7CdhW1nQKVPWkgIX+n
y4fDp0VmHfWguLKR1ta2sGrn79LlQPSYYsDtHR3QB0fYlzIpWasQQxfaP8DzWJSF5ER4C92sroT9
HBGxR4wZfN2EA4m1/T25YhxUsJpbj8BYaHJjyplZF2yelbDexmYUqGorMvdGG9C1544IPB5QLM1v
EcMWE4QVQ4D29/2hSxCXTRXg1LVokTz82FccA0jvImZl4TQiMX6Qo6nMdMkCpn6YQw6sXhUI90om
1P0/ob2ZJjGPJjbYLXu6fRM6WBM4gMi6ffljvImIGVhpUXuE6w6FH2XbGJEG7NWSjMffmUawMPXo
RraItLqJlYcSpEPZANk6BoIbn/WkC6QLiaIDlWe9drGKyWO9WmWt7Nsa8HybQ2hfA0/aFUqxIJr1
KfWDxZnDYGxVry7z5PS5A1LGHzpFKFrXslu2dZL/xkcJYXJ2JdP3tE5xGXKUf+nS3a/LYG7k0grS
k+ofedxatFoEwrTIo5u5BAOW0Xdr5rZ+vXLnWvldvGP4wRYDQEpAHkSJBXSaIPspy6vbTc7C/Odn
QJImMxxInZlOx/brnWmNqfvhXJIAsO0PNDAUp6iI0JAM0TFLakQbWE50D8c3/L6CnJNiRsEFQMJy
iE5OskH0sApzBF2JsoXjrYxte2dBNR5JWT+EJ64CmmMl2cxQ8qSiRNx1SwNTiGD7ShsXHMm+X1I3
HNVw+Z/zThOY85mCXswntHGrbx2LmiPgkjw8yUOoPCyB9Rk7Wmv627MUO6G1ANb/eA0cyfTp/soN
WzZrYXTBaw7HLFBEMDNBbqKfJd7BGlkusLQ1BKoRvIAriQdnwWXytTJgw/vkbqoFvA2gxqIJOjpQ
WFgcLSkzgECIMm9AfER7z7gmZ2XKpvfRPZwsaAXGpXw095cvwCBr+eKmH9aufklEMpxKyKq+Hv3i
wZEbtF4SEKd8QsQM3MCBJbWh4DNf1n4/oMsxYIQ5A3SkdxN5ntl/y1IMAx8LUneqZRAhKk8uskCu
m69pMpxjWbYZwC8Aah0T9iTIPmh6ljwOd5DGZ05VMznOXlvOkZOsmjdpdBvhN43s+rdF/hle65Mh
VrubtXhiDH+0dliunEdYYq5A4h2BI1gnWQeIpa77J+JiZ4LEqq6f3l0V5n/SfMJBOYtwxVEgGHZJ
S8GJQWZsVSPnkwlM12uyFvoCE4NABeyUZhb+mychyjvwmagWWkiyBiO1JZAZig97zcE0W6qV7qeT
qbstHnFuwfeB/w8ghynwWWyY+2RMq1/qYllaHbDWO/RRY2mLhHXNU9qdvpcvJ8Z2ZkqWiF+wmXT9
RZ815IEy5UXbWjyXq+p3qlAYe0/so30F9XBXfw+qW3wUerw1WnmHc5eJNHEepkKXLt9qe90U2W8Z
wOHZ2wrF1Peqor43mN/C3excngPgYJvimqobKwFCFaaG/n+wWycQcy3ZJ1wjaIimG39WsSoxpprt
0CUMS6LWJwSgzmhqgcU0PySe2Rjh0V4Fg2PVJl4LDAs5WR3HVc6HmL51mJaJB7ydoW+Lw2KL/DWz
f3mxwtsWbxQIpM4qgErFVnxfD5CpyBWFBkc7fuW28gDZds1s5yKQ+InsJKwXP0EoT+bPOzIGSkSI
1NDp47diAhicy/7ePX5plTOmEOyeOvC0lLtI1qdX7UsFoSQDSBeaVCJljMsYUrOzlnBZCySI21en
vBzCrxruHbqMz3qfUKA8zJtheUkC37donxHToygOWwSk0v3UDJjTdzse/DYZsyyzNFJ+syTSG+5e
fntNvrs4QbBk0K/Kb17bP8qsQSgsVl1IX4wJk488tSo1lMxGxjBZh+doSdNqQJ3jfFtwALVCg+ZH
0SAkbdP63dBO1lMYgbLlazjaniBtoxES9y96MSEqupyxXkFPA74mvcbpepxqJfpu8HoBTEApPVgM
tMHhzOKeYqoAR45sblsernK1grE7L0G9bUUUfQLd5qNAjErLQt4j8Ss1r02MwJFTURjba0nb68Xc
UZ6v83x/EJmXJADORuZ3PhZpoBiq6GcoEY/QMa+cwyQHfuABN/8JgfVqCnhRHmsExmzz6Zelk2Hz
rzbqT0KAvZ4q8EbM/odMATIWZjUeCh9SeVaV3o852wNh2HxofItbYpF1vYd0yM0yiLwrda4uCdME
/4xj7eYCgUkWxtAiP0QlO7VtAMblknYpyYvvFDdtBX/wW25Ru2ibrz8xcVXtmD1okCmM8An1DLJR
D+VBoYEdUw52N/76ylLboG7ZjVRay9Eb0xd83/efmLWeH+VU5v/W/7HwP3y8+l/aFGZj8olVS1MA
ySFooHKNqkixzbJtSiSwhBBHppnA2hrGRZcF7HspGmSJPxSdWtKXlzYHzkPBcTb76LqBDHtXwy5e
w+Uv+0VQR4ApJN7BFy+wg0RG/xWcNAl4bOl/jLlybQ0dmgoDQvRdDPAJbOfmP0c9un9N67g9H60n
DIbO47y9NL7cAUcfLvATGYfRHdM8pm+SNwbSZzlG18g6+6aXi4SOc9b3SWiXkEK5aNJKSTLR5EyU
A4w5q3y/RUnNViQtpAiPLwTEmKWtB736LuzAmw2Gon7cVXIhlY7s7Noprq8V03PhTUbU3MSbdBJn
64OJjCcOWjghfz7Kl6uKLwRDXpjR4nduGgpviEMdezDM9QOuBIqiZUYADVf6kIIRz2UdFX8D1/QH
hDlIgzUP1lR6VisnNFB3s74Ub3jvP2ymlMaFKZTPDBQXNeci0ViZyH7mJvJaDLiDpTaDwoKSkrqE
NJQkvk0j8X6RdkQgvdvsi4hsNHFskjnP1432e+kBN5a6dfT4PB9qMwq1okVWWRxwfYyenQvUaq4D
T42k5cOis9Ea9xzaJeOTZEmsCWWkmoE5YfbJMZXu6cJSOFMUh6gxj/7gcWlRfahdLUzCzYVuyoxf
ELPBEWG8OwQJuEq9CMcICHwqIacnm6pLyCnwI/buK5GSIiV9BqwL6bRZ8SWBA2ZIKqQ9x4j5Dkd3
mW5IM3FXWA7y/5yHrffDDp6KXHU/+SsOlzoVLnZEp8DUxnpI+tTxQY5DgJfLw7H6MiNFdxJ2eds8
sSgExO71q68tgPlPjUIv3x6AMwxEslUPAEA9RdQi+CjmlV8oZuGePckgMXBFT3RVcJEVmF/hTjmz
wthh6p4zBuAt7hcdCTyr0vyHf/gLwcNd3tdqTkRKWYYAh1rElbaWPcdXvXK0/wa6XXJpcEyOGF9f
LjawymKbxgirvDMP+WLEclo4WZmsbO5NYSby9TG3NQMYAqnpFBBrAo9fkLtsiuP/4TD6xfFzHD2y
47jGMLp7Mua+r5rnOfaLu093y2Ymwz/3piObMx2o1Y60K3fL3+UiV9tWpjMLW+hUcuOv8K4F8n1X
oIlMXZxVeZrz4BYdmiQ6Ry5bSBKS+J1VIETZZtUzBrnQbmbRJoq1AyiZZOX4CSnN066534dKV/gp
4RexUMmgc2IRIOnA3Egq+f/QwWLtHBfIW1DgREklFgp4QgSOD/BthIobsG/ZsC/73gSSzYip5heD
4IHaAfcqfq3SMtHfRfOr7EQEQvvjOag7oHJAXe69B9Du75EPaaTWS1Zs3BKS6x8ue2Rvrutg5Yo/
3G1Ls30kkU6VqrTiNKT6t289o965O4wShRHxRplGWnOorBtkpteBAhYK+8f4kdnMCA3o5eg5jOT6
pe/WMYprcERQ1c8eY7EznafOvS2KKd//4NfRmBVtkpNbaqEwTLUr0BQkC5Vaqyp3FNNnFtB4f1ed
alDgSHWvYD0c+uX5g2slX8YQMfX36sLWaa0I1SfKc0z9ahDO4HsEdibEW3RdUeAOGrEll+0vTHXC
qWciP4ih5HFxfncIw9kSezNIdBiNVn9UcPbI956wxpOa2B40BS7cOwxce+F5Ad1pSOXJa2HGqK3d
+ARdbiWijaQ0p/NCgx3LIOAjR54/Eej1TyYunRSVS8WL7bzrmX/W+D1coqAhKo2IK9CwCrCz7GPI
AufF5Yg4nDs8FvEX2ZtuCM81H1lLXwh28xIRdMHMCMeAUnvYQSy3YT45Qr2WooXuU4XxtCEVJPc9
SZ1bGIn1iaznTflJK8zvOqpu937INCKDH7g+9//5vFoccdUPYPwHTgslsm62cE5a6eRlr9MjRqPr
dWJkhtLnEC5MTg6GX6IpuE7ItbC8okBDuwya1ZjPZgC79+NrZEtL1eMi7hEVrw+h0AZmUTE43OrG
A+6f9foPVbMvSaTsf3icanVWHnrpvqAuJ32mc8IHi26WJMP4Rlz/WayjqMfG/bg9k1X1XSyE6VOP
5gM9y2ZWwys1WIbC6BL46rMxuyjpVPv1acFidE0ByXphUHVAyePA0ZUYJd2g8PWZnubcQbI9ucI5
m0JEEg9l7v6sPZ0CyN4U7YW4erRsqWJCy+OwuZmUVmwCXtc7JJJE/7fWacDwWpeTWqRmdkOe0Woz
zQgpEziMndgWlZDFxnVL/DGQAAZvKBq4D/1sVLKYreE/8Wcf4HDAxoC/Y+VYSEeZqZallsA6njjO
PSwM5z/Lv0EVL2VtjXfHM+jOqB7hjDpeZE0oGSTe5XCCnGXQGto0XPV8Tqq6zH5n5yimPW2OzORa
xzDFcdv7XH4OIlQBOViovSjhn7ozSBBgdTWrk5rhug+9w2jKYe6qkrPmsUxX+SNDAthdPJtda8aP
P5FAe1/DUfnqKD/Pv93GAmw3dF1lOXJfbng4QWLVycMeFWnJGDED3pypC1GulBipJToGGg4WJzHI
DdN+6f24279vjWKJADoYapuPqAoO5NxzD1z+7OG/9e1dL0Py+gLqkwmpVt3DRxtvLmYtcK9mD7Jk
nuMoi6nz7JQspxKPlma/hAMbDoBXGn2ZO5jwiJonzNg/dVpotyWzmqVT/MOhWyMDIB6sJi6h/hGf
QQ8m6C0NQpsrE5jSniKUcUOm7x7C6GFC0nk1vmP7oiB2CumTc3vzFBFOgl9mY7d1j0neWZSktjCX
Id2wgkVpvrKHWDfmNr+v9y884pnPd67QCeEoRbbgZKKBCSxBUXoCqD3qByhRgY6y/0paS8/8bTeu
2bazWWUYEvsRjSxBB0nXDS6NaHWf+msWFKimAg2HzK8BUDZ7nBneFVb/zJdNWYWueGlTo6kcK4g6
vpF5wUu0VpfQ3VIH2929QaG6XokHjWO7sm6zz41XWdf4qWw9lpxLry54q+yShQxny/m9khqsjS62
Rgz6HPfoPF9NPrToAyidNZJfawchPQLdkfREzUdUsBQTak9YhxHTsc6DAFFttgZGeQbuqQJ5OXaG
T6LOyEd38rLD95WUDKtWszn7/EPHik5rLz8lIL5kkUevrf505H/W0YT45CENZSU0awybwyhb6kxv
p49MOZ2uof3o4ZNqUhZrrIhqMNhTQpO1DtMafvTrNsloHf44NQ2DemieYGCk4YAvR9ewLmvAlkji
lYlzKJwRQ2NXLcTzxX92RR5bag5eK7iNqh1stx7qTO8z8+uiunZ7SKaZL03LOiyEGGe10Dvf1pHK
JDesDi15xm3pP/UrYXkIfKDMQu+WhvPd1QtVqWM/6O64jA6dMRtHy0QGGs4O/hjNYBOZgfewA03w
HmDdhYmlaLv4juYoPzlpBts3BUr1APlYs4paaPLGRA4gXDWyLSmkCNZvZyoSYdRYW27iAl42D4+d
pJCvQEyO6cM2yfgVnELCcKfhzm4LjIvc2DCrwrCDccyIekHABCs95ws/7jS4p0T8SZcopbr+xWlM
N2+4oXBVvLf68X73G71KAceiScsG4Cu4Bt/soA1J/80Y34yB3dKJaguu/DcKiezSv8GyOkrWfe4v
tAPI/z6owsAKiZxxPJTc54ZHKK0U9XL0BoH9SVOMyJOC96s9fgB5z2r7RfT5jyVSE/gYu/VjWRIw
f2u/aMF1bD8CQmxa9FH38Uwm1t18pMp9JLu6SOhbhviKY/hpd+cFDupuyqBey4YxQz/V0TOTDMGQ
qfc+bZwbvszdDfPs0vr9XB0XrdncHDCFzuJab2Zy2QZAyZJpcUXdIQSuspnNKuVaN0MQGLCcw31O
q1Kt06KZpKCMaYja2yxbCTX8AMv0Um1rmGnL4IfyrKlF8T5G1bPCthbFySrq63O7rhH4dDis+BXu
9FsO8kxoS6qBxn3XQIcUkXutnx6gaoTrrwMm9AaPTrUoFOHQZCYSBDjcjnvxq7qOys8XWzwthAr6
5Jhw3sEQ4rfy6DXRSAfIGpi8ZOD3pYHRNs5ZqwwbrPG91KqpOnHDpa1hGDu7ZunQNrlg4i3351lL
tz+DHRy4UAELS7RCac26Cuwt6c8rju6vzybgMgrb2b7pypSd0TOqD9oBDURxX90ELCOtFrJLgXMH
oFhz5UZ+SerF05evfRki9SkHl+fw0xj+K8oEb1I6IBSvG5+7BrWlstEn9XaGM7cu4Ecbx9rAEzNX
4XDzdqcCC9eQPYgJY2JeVd/3F6A/ZRQczGqLJiw2JbOIeKVIovN1iIULiaY/0GCDz58dZ8pBmiPm
pVtif0KxzU5r8gQZ5PupiMGin0mZgkeRmT2bCyVtc831RbkUWjVn+1SMeCO80w1JujMXCTGy/6ge
mShw/oFLNWAl69jCX54SpDXd1snonb9hP2vzv255H+iO0AzvnmA7uBo+LzpffTK4P6XFo6Nqc/yk
XFpk8tR4Xes8BDOt+Ef6efmxHC5SbfHs90WUQy82UlSzGQayp8MWuCsok70p7t/Dc3PwRt7AoT4b
aXD808dMygZ9KxCblXsYVULylkymVdAWrugThUTZIiinSBWHO2k/E83+XhDhflzeHzJ3Y7jViIEh
NrIiZMIxc9aLKFim07PZuZpvCAhcd/TlXMbZ7zvhjFOeeR8m5yIB01NVb7BL6/zDSqA4cvEk404J
fvz3vVg07kqnKXpzkCMWRZjHdCfvVoiOe+mXbN7KEgbNZsFgnt5yuCizGThKLvLizCYwtofUqYXB
e+jKD5KYuTO1wyGL8ms7Ux7N/wxaqGiv8ltREBsN2udwV97k0H2Wy1pDmVUDrSUnftlQs1gFmE3U
3SFAWJczKpHwRaxpe/u/n5BmsLXGEZBN5xZ3XAh/o6HVf/vhSkH3ETaa+58z+X/ZJ34IeYIVsNzR
J6Pp1B2729VuBY7Qx6CU0tJBV73X3+zISEzldYRjqeDdBm/N8Yw3SW94MJTMoKonpMiqw0JTrluA
dsBUwiXZXbrICCy94FT+ESMURN2ttzuoUR0BJqAlZXMgBqivo78blcqH5lR5bju9a/clNDQE9iLc
Eaib9NjoUSXaCfbC8Qg5KQxs4G+oNfKhCuVpN0Rm0DcD6ShURVnsAsf8nWR01VHWjpOzibP27+dW
B07c6rFYszbznpzrChkbWoCL79/Fu98tmDCWR8nhHq8H03jDnMP5rVlRTAIMjFV6rmKpD+ZJzeFY
luUpcJ6Fs+41zzkN3qxJFID5vGPoqnjYZfthSHBGeldaSHUoKe8qQFEbF1Wx46ppGLhjXUjTR8qI
cVdQKvot91TtiFD14UmebIsAe67Jzz7tpooaCsaXb9g8xBJ8MeYkk0ZEb61EQZa04LQs0oOFXAUj
w4U2XNWgrYFDhHVC/j2Tyl7TgDsA5OckLhtd30ufJLF9+Yv7fR3U25dgwf3p+2+Ghb3RJIaBMlOJ
IWRecM8+SUQ5ONziTRUvzmGsIxZ7L318NasCbG8ob9vdbRHekv/H2LU49zWV/zZs2DSItR1wwkUg
mE32U6WkVoWNeJppI4INxsHmALt34B2gEqLPV5NqaWoAMtXjCvaQfdeZo4RRQKCc9Q5gcwY6rX+d
9heJJT+SjjXSPIoX3LqT6scL1g37oxQIUM3wJdqbe7fTinij9OVPhQtmv6RpJNps3OZDaRd3bBkY
9z40XhWbY3n2o2ubJF/zeIcub32LG7am1DSdphh+nzUGyahRr8Wb1jwKdZo3FVZYxNzPvIzgT7Pe
O9C/P5If5RE596exDHn+2YrQB01wcQ0wgj7Xg0B8tBR+fOs3Ml+tppOqTPpeG8bOjccCW5nyBSNc
Np2fNEx3iafvp1Ij4rHOmIDd975yAVFfayhOuDZqUEXKYSEViexbuDVW7XmoIjN+ygKOlTY9YiFJ
nA4A9f3xwYRnMVr5uOEuCrf0oRDjWMHaDs6iOXoo/B9UwbI9XGRy4JvuytBRDRoHkzglv0S+vteF
9Fuk2Qf8/HE3giy6A/0dncAGDKAp83bS+uIkR0kbC3Tcadwptrhpcdz6Ypt/x5AOjieYVBO6clR0
x9k7vxNhUmafhrjPM6EoLxxb91h09SfDaDyma11Xdlk4XJ/VyBNVusUlweV12ja53LH6PAVHu0OL
OE6Qr6XczvvlCZOSgYxj70SpkAjF/k8uWYRqS3weeakoQgyXcnSbaSCG68XXtxCNsGuvvKeTdls2
f1GXhWOsc9KDyJHrkXBAQ7Dc3uO+kZq51EgNLIGECrcDfTiJT4oXgsOSu4OKpJhdRrZWwXUk7coN
L0gO9d843O4VfrknvMifPjagJKVTTGfn6VN5W4sANcuPTurPLCzCtpMSVy4JVS7bnLpxpW7J8pQ6
+D2G3/8G7IleLAVAWo81f8sFgPNav/99lFkuLqC6R2BqkzubL5vLyul8Fo5XSaqgvfMs+HjMhie1
dS0EBBgJogoX2XwKvJAtXUYyxQhiMdCPAZhDt3TLpz4aKiLvhl7HJjp/A46/zJYBMPWqoRWJgyVn
g8SoHN5CWx2gAMMOci+ryrD6Y43JZAX+Y8eXrWMsmyf+VnAAvrHabXMy/8+pQ08XEZlebwpieM/+
5aIh8ZEpsYg0FjSXT8NA3VOPbsykQ55cJcMUdKCDS773teYDh0LznQYPt8DsuoOZc+LdeC9ZW8w7
JlMOhM9T2Ru2p1fO+6qBFiB4wUi0pstEb8y76+0V7SgP69d4JCEnzOExq05xyzg5GEI0q/1TjK33
mT7+YBGcy/0/s0OYM9+0lcz0dT/iP3x8Ss/KqyP7MzACKZAsBMWo588fmxRixkLXYfRV8wfybcyw
4AQ4C1aIRHQbAbLw0J/5SbsNM3a5/ZFIQMQGND863Vjk3+tZMZP9sbzz0r/dCuRO2vh6nNHQTrpp
BHF2E6yVbmKIWXohBat4TUkOSnJBFn/TiYd20NmeNifl9F8+A8emP0bAHBcWaAMEoW75gi59eN3x
kdoD5M/7S3T0KG8sVsx6HBmXoO36Umke0PJu4DlvirTUgKsp+gpSoHqcI5kv3D6h29aQbe6vdnof
2l2UCxzdzBrbv8ddEPbUKzi5zJftj6+JMFWmKF9omCoXCWmJlkxOmWBS8hAl3Rq3pBukFVZkSi6q
QixahSu7FfZr8pO2QtbwqoNYmm1pKq+gFFjQ9MTdQfQqKRP63/9sbrmW+mT2Q6mfbtKBAghw54a1
SRSG5hNS05U33j/ZeHLtovv0N0lc3HvfrIac/pc0+4C6UqkJXEPMcdfxtmV67uSjnvEhDCM89Hcs
f2wPiewt70hOkt4VZ9Yd/ZeontBMg+TPXNIZpGMbWj4n/Pk5AaL3XPOORPFiSQ7MIF42/cks8f3d
XmbvYWd4kKsJ4V30mVlt8WmgcwTT86uE935FP5v5P13IEda+T00ahqkWFqnAQqC7IgDB7EitHNBI
XPwMMCZMajR2R+FZ016y+8jzC5qGfk6tcqJkx3oA1cZyMCIfC66jqCg9Dx2a00UaA5JRsMLfuCEq
g2HtB1t0gBKmHjloDMHzYAf1KnvgdDMcOPQW+wVmNbJX90AOvjxLkW0kNHKFScLhmIAa834EGWaY
5aHMoSiwlLpiQe+cNl8k8+1fR+I3cSYQ55P4eF6Ip7512DYYcpK2vT47TT/PIsL/YR8zZTspLcXX
XXYXOV3O4DoVqtV4xHdUtNQcxxqLKrZZGedqhlJl9PxqddaoSexUK8Mnpm/jTWBZupYM54IRhTtt
k6cNPOT3Z1Pfm3KmUmcbO6yvWSQTtWKkXpqCHKyaH19I8gXh1RiSnzrmEjIAB4fb1SIgknCEKC3e
AhHGhTsT6DEYlMc7PWiWKTxXLxi/oEoUz6BPQg/WmWabHAjwKtx0yjoiQvYbUD1N4I0uTePd+hZz
Oagp06jpQ+eIqjQYjYpqBbgzOOyaGCAcYlpo9LiS3seW5PPvO246rIzyOWlu3n9UE9UNp1jcFYp9
NGj9zG6BpeOo4TNRhQFQX+ejHZP7mTy87cyhEEfKSvqCrTky60Qazi8ofB5xRsG/NAR6lh55GCR0
QwWYgOaLs3G4uIJETf/P8agrADOA6uDtA6L4jfSRHwiyfvDd18WB5hIzjTV2QWRF0J87IDDx6/oP
jHfq53/nJ+Hs5p6s7U8uMcIVYINQmwrKHFia3u1X2s8zmzZAPkB3fLlZDDhFFkBkYPGR96qo4GAU
dtzpa6EQ3VCh4qfFkbwcYmcK8kd6ndNJ5OFBW9xeDF5H0R0Tz98GaXeW6SCIVLBw0GWBNDomwLjy
dhwUPy45v01pILPbm5CZBnAyNoxZkryWn9SqFDHzPLfFiE524Fw+OmyDeK9XpAtB8CqsnGXtjhVK
FVIuc/LyLQargCP3kv/3x1f7TxBKcH3NOqB/lpWbshkE46VSkcleVYMgha3jknTYiM9gaQPwDwAt
6d2YlqE60zhH+0vxcM9W7X8yhtZGxDAk7ZOa0sZ1uGwjApWURUri7rngm56Q067obTF/2xxIPjoC
UFpa2JCjWN4eF6K8jYCzcf61RFRnaeZyssnEes1RGSfp0zrkz7Vl/yIYmZGKT67hi9xde9T223KL
oA3CXsWa/9CVZOsxyQpna7OC/m98ChgD1jFUu96XgUjMhCyrA6h7qnzcyVfs1IR50jIq0JCr5zsg
fW6V+0+dy9Tuvf0Y7VisqSnTXAq75Fsir+ceAgDxjMmR22N3gxO+vAPnB7GVrUwgIfv/wUeD6cDC
k5ORGdYQgLRMciuJCOgCHj/jKsVdMpviJMKaRGphG7OR/RTC/OK8UNFQx/lYg6/i1RssS/2fZbrh
eowEzoqcMBCN3OBzYf1CIegrreBwvncBSiY4wpNhZqt11wapyUJ/7H0wyX18rpbnMULuSQY86Rbk
eybYh0bBtISFYezzQWlS3ehJHMIfrp/BZOOtTE2bNPFoLZ3cTv4/rx8IYiQfjWUaxVBzxv52wPLb
q8is4VzPJ+V/1MvRHKuYpJaQDSks5qk61GyU0Vz9hkUiXwG5KukHCId8e/OyJv9OCAXZo6UAjaNx
8awSbM7WUxLctLQW0UVQMwI5w59LOp3Yr1I6CR/ApnnTJU3TIZhsSenzMcBycQ58FiKpo+eTtwx/
hQOIcDubvWsp8GxR9zG8EW9VhmdsoAbb1Ox3VO86gBJgC94bzg7S74oSWh3cMaYCVZy8Pq1wEQFG
uGkDVnJcLxkhdOYB8g1Cqj0uiYoUO7LMpkI5Rd5IiQ53WSnFOXjKymvlipm0abHMyzOSJNcXjaHY
dxHeuZ02VgU0u6cf4a7M01KHp7C8AmnY4DgviT1OO0qifZ/fImkguACVRs//B0ZJ/NUVLXVLeOdu
nRNUyYjHqZdJoIDooOU+I4frMNtnY/7HEUqzQwmuHUru2RBXHGRsp1P4v5q5nIwoFMeDV7R0apS6
Hm3H9BElvD4pJtYiqe14PR97W87J+VX08JtGLZBeAmGCnd99y4SOWKSIllETnasTLO1xTqgAISRz
xob2OqpIR27Ow+c8+l0q17NMKB8lZiCl3RUtZ0gB2Zl3G9UF0/w/hzX5sP9jECBvlS2Qcn5rhB2M
51uQ9txFQ900Xl2ix5AD9Htbs7wsgRASZHuJ7E03dnW1qRMQwgMGJZ0/uttgg+RnBHizmeFbh7wM
MK30iKxZfEOYRFiRZ4mj2IiOTpA01CxOcPtl1yrRHtodJQJuhGL1yiwOvtd6uz+eTaGAvnOFCiYO
/0uY9UNbrXo7HDIy0wtcpUSZ89yWmGre6K42VmV0O203SW6uwgsv4fAHqxEVU9YULKwZR2+goowa
zL+1C+05CD8tc5AY/aUhpqdG0+G1HNITVfxw6TsBIPT/tZ7G4ZINqRwPL21bWH/9SkPcTdNuOjS2
W0MrpjXdTuN1tM1oBVodWXrHFT34r189qIas2teBB7jvUJ6HQejyijJjuKn7MRL3GEuVciKrWlrp
Xl3I7jnYvkM8a1tqoCVwdls7YR0YFgvg61WKQEvgH8x/9bmXN8gzHC3qo7o8h0+ZTF5IZA3AKgH2
lt1OuLE29xFIrMvcufwg48b7B+JHxWaTgQJSephru15nlkRFBZbXjwxvxKLw1W0LCPqcZV87SgY9
/aDG/ZTDAG64FWnnAtcehGDwPlHjlm9qPF2G3Q7JAgTbWMeqEh7Fl8D8Zpp5zYC2QYkN6ZTOHhK7
mBmSUApK7yJEulYcp7HqkP04mb1WjLS15fKAxujV2i1AsESjeU9M6OdborxOWgMk4Z1AwVkZH+jD
PyOsrLDudOcv28pf8VffMZVkk/WLl3PLgYTOBdRNooHg6M6ryWbwvYxN+sh7sS4sCqKD6fUZjz63
hNhMaZpTaaqKy/mmTd4lkjnX+ZzHeKoPuitIquszAuXOrpue/oVClsSws2lTkoWf6kpSmmq8uW9b
M0dpwMxENyeMZr9m9007FpGNN6+8MuvV7GyC+Fv1Veot0gKXknqjwoEXdcgDCq328b0FB/tzZ1eA
xEdyRuh3YGEAdd66GfTVK2BcFng/3h+lIC4pNpGbjoE1Ro0IGTBQ5gtGu3j/iVfLs0LJnnzXPF5P
M9Sj5BxeWp+PdmrpRk3H7RIIXtRAgORRBi+CBHYnFJpBWb9IZc8mTxol/nrw/opr1n1PcJ4ZKN6m
8nJsVKjo54csZakXw/Uyomb7ZEZoyTMKMzmOAJelIa7wWwFTtEAvtmIekeAXR/iFuG+h6Q3+SUxh
lFnmggCg7oOWwJVzYK20PnNF8sVYbjINuGfLF3RIUIDiD4t4BIcduQJdwo46ReMLYSw/HCft0UC7
ATGPVKiA1f/sM670la/jW/zcVaU572pXkEkKTBFTe8RdzGAf7xr39Dr1uWUtLfS3q22VYZQpDB0k
twzC39os9bx0jEe6AJu7koRFhXvW0n96wCsHOC/GSBIFZXAsij+klGkOwhW5n4PnIaPrjm4DYXwB
BptZg9d/ztXROKo62bsh3onvFBPNAnBsBlL8dMc3RJGRz23NukA0yJCMOXsu6XMtJz8ko6cLh7gk
XbP5IGmEyluaUxrw1xcoQ0weaDETCabX8GQurJSolKah4NzdNayXTIlpI4EMFN1+N6VPE5QjS6La
CeVJgzux+OyeP3gtxfSYBL+W98k5NjHtYlRQmzrTqQnnJOoWg+nzpC9C6g4dIItm9KZim5GjKWNU
FIjchkMleqFx4bivFz//3wJeN5FFxI9zFBvC/+HUGBShmq6C190wZJY88b8y/xfl3zc2k4XjCM/g
OMFSAtPYTTeI6NaSC6A7nlbP2jisSx2s9sdg/D5KAKjckm43kseT3Plu8T13TDPnJcEojpe7VMZQ
6jPZcRgtvN8VrU8eFcU8CHqvVei4iaYwf3dw+P4/07Zl+KSqCGSIaL9TmPZG/kLtnjP35POrSV12
GtLFsaUew47Wp8MEzRFs/vjS0rcQEKlYu86mqS4/SxTAmLZC/l6q3d2fgO296djS083uHz7dpPff
Vd2A8nJdJSgW9V6/XZzJKAQo9qNJesrKzrVVu/zrcMl4Xrigme//SU5QbfKBn+kEYmQEnWmPGAQN
vAdN+rYXQJcETIV+S0MqCLEHUTAamXIcFCSnQzHNE+8FNcQJDpvVlEtY0pqrnDT3xmgfLDXNiZs0
Qp1qsaoWfZ5lo7xuARv60YdyMmuCJAAxKnM4MtGIpW5qvq2zUIYmk3wVuXiwtQkJrdNb3zwTv2Ns
V+yhTWjfbPz0T0T+655r0i4lRyMnlUqtHaEv6a2YZ0C5oPYSqtgd5gJitWOb+xXRa4tyTIch3qtJ
FSgqYZ3EKnm6Gkif3vmPfDyE1SZKV9Lmc8s1pUBqZt6XhZc62bAivcUKtyLVZg+4OKHLMDUnk6Ps
pG5ljx8te+xgP17lmpOyXk8mY5QE/zqvTdfsbHPB7uXg8YOJnoTgHMf/MFP6pMZBbkEXpuop5B0E
ZWzj+TMhnwoQO9DaSOV9czSCNydBD6nGoY7BlynLu+mR1kwGfKaO02jw8+nw55bpdp2UgOQkPkC8
R4x7FXHwGbMTrvqwQDJOSWJZWzv9+OKcRpolg2qJdG8xb1IeS20PHy0HOfDbx9SdzIJ1MkDBGkCR
F7eJJCAf8o6eFLOYLKfC9yPYjGmYWV9HV7K/RfGLQDVKSATGT0fN9JtpvWAVtWG6ERYrJyS+DFE8
6nC2ZzFDFrjygrVIVcbJxgQvsmQO/gtpZdl0zWT21QqRR3kqp4OB2MN9N0eaUoU1eEfGFyqx/xyW
Oy9dQeRwo6EbrKO6ctV0UPN1sTqu2c1Rt7z5Vr+g1HkKRC8GzYl7eYOfzX0wVDCESVngzWuFL+/d
qt0gJMzEqLATXDVEvsZWHGMT1WCxEFacY4n1MMrw1xDJbBl89nJJS02tCTa455t1mJhiCMST1VWE
rU3ygVUt5EhSmWZqjwxv/Yc81mdH3Vypq8jsRmbs4UtHKAK7s4vndt5xWbkDpxvi4hqnCgYMwHjL
SO4vcQymzBZ9vKtfnPSLYlj1LTGNSXSGy9DhSSMsEgVcXw8LjhXiVM0XhD3Fnd26bdqBmkAridOV
U0Ni9gtGRWADykCUxlDbV8ArNMq77hwxt4AWrUI3ZBIS+39lWpO1IQsRdPByTfhaPASWMBTOfArt
AQXj0ezW4Q81OwlN+giM1ebscK2IMMELW5vDVRmpTIVmArx5Srs9rwhyNMo2POwBwVZCD1jJRJ4L
7iiLn5bxjH1WGifL42FF2lMn1UWl5Ynoy254aJwisAneej1RHMnFzOiJJCZITq8FNp0/aYzR53tw
UMbZZBiHjLkRCe2qGoORWgT+/Rmx4MIobcbTpi+ps+RnFR7jO5mrI8CyKieeCU6OhJKLlDbWv198
5ZsD1jTxftsqgZ56DRu/LPS1d1VbpZ8bPr418nYJCjgaBHh4h+ezou/qi7y1f0NmqEW+TTV5Ql8G
sCtdD5WsY7lsMJka3S9ciV4v1K6uiesZDDWG4w2ACcvDmhlIKqqMxevon8CJvfLHdeOT+fivnRX9
XDn83c+IXCBflNGErYPZvK6EgISeu/7RO6CAWpWwSLXL6AVSturLCx2qiV2SA1wrzO+w9E/TgSif
q1Nj6ewZ0tkuab9xyiT1MTcOzu8qN5pPcJKgOdsUxWHBOztl6p+4wCcphlHWX3UtufTGebgNh1bK
H6E1ffTpMnVQDGOLZtpn2e35YMUNtiN8osAFY/y7uGoPE56GyD9pMpTlQxUKckSQ9TmBUssgdH6W
EeZ0Q5VRKqV2RaQQ3aZySkywih2ZVsisk33fX/u8GFCvuECKUxtdWHbXpUPIFBVDASoYs/jvPE/9
pFV2J7grEZtYd7Z8gx9/paxAhlvjNhXw4K/jC+Ct5nE7Oe0q0rBA0dABrxmLz8BpXA9EkPFyH/6M
+EhnHugPbhuXw5nZiaNL3NlVEANvAWhE4NoLu8L1XKYwK95jHtS0yGG1UPlch01DcUiw4de9WfrU
dCtvAz0HECQOzBG7C/YQF76jxvPaiXGZPatLda4o+uoDuUI8PImA8B5mXWqGj3FwUq3j0aaVKDMO
cj0TxMuvBYR0qElfl7k8z+lofBfMQnILRoQQBD7x+riC1Ca4kkCkUfqKW/Toxg4w4RO7oQqFch1K
3CkHOwhTIoUvIdY0O9nOGi7ckzazDi7ZZ33E4blc6tweBnveHv++JVNY23pfaRqPXQ5lWWGQ3nT+
DZGjrHV86iF2+2JyruHNjHXI4Wz5sCseCAPNpXJGNOpqy3CMSgIX1U9tZ2OV6LMoLl3zly5Zi4Hb
kKuekG9C/7oLQZffjtnoGkgIv6jZCFnuebSAfDlzOhtx41vbGLC9NxdGUBRt3ICKlO/pkdvGOLjC
C0BDiif+UDXOMmPpfITTHTL6DH9FZUla6xe2p9EbN/wwc+WjpRisrAHvRxBLWWUc9/2u3T7SUQtM
cE/l2MATQ7jj6t+IV7yGd4F7eezPjzS42P5kAGiShtMjIEL+Lb9z623cea/+UDa0Jt0l4NyzE106
TsdVh0bzexwJiUYO3cL27t+4/4heRpJ4Yb6j6Sa6Csh+FBl7ZUp+DM26YddaTODy9RWN8KuybEUZ
aCHfYATd/Kh4Zsrt61laBJDXWWGkXRPeWE6RZLHt4HWw3TTxt70ww5LJtCUqHZB8D+PpwSdQaBhO
tsmomzwlwHue1ut85DinfxMjCnXYhthvYSmK+IvHlTjGwB4AY8xkm5h/I8ucAsIvGpAUHMNY4ph3
HEsXvqOCWb5YLGDmNbqjPP+1rxZhGEVTL4Gegz13f4ZyhicP9hVInU1155TbsBkGa98hUvZQadDZ
rIwDMs+yP1pMrPpQ3KIJJSNamLbKNCqXHxgUZ1wOwaBARAXo8VsP+oYd51KgSDieMo1rF/3tWkiV
XP111DWZyTYzeZ8QCXzEnXc8+KSDa89aCCb0uKfnLLPYh8DB0/rJlzkx64u86+Q5i5QkVJhBmeZP
pxj0mKt228MTo7aaMNP01P5SfOMELXmG7yVCk9keQMitO7zuKMh4oGlKAA2uMASHkhEczpaCGEZY
NT1jIkpC81vauA0gtLEUETLjHOnI5y791ITR02sL2KIO2nLJRTEeJy+XlnuOfv2IHJWLQS5HamSr
+5Jghcy/tdBhZ/aNunSWKGFxOSHPphrLEfxJko9jDGGeuwHz6li/dKEmAg7Ac1IyiWnkYJqIuVaU
gIbBf2a/Ia3iEXQLdEZJkhB2YYiiGFl2nAlToMJ/uFDEOEttNCe7WQpPLqTmwEQC0TqlIobwwtsg
5ySmgR3rV6jJSASKNK0oNsRUyR22yShqUjIMB5XZUtF/wFRfyUlYdoSMZ5pYcKSpOssQtgq6FKmE
ByY5Msc5NqZe3TLUA3D9/vFHEdPV2oWxaePpTbVOJxmHtshFC6iA3KlVooyKfn/UPE7p4Bbc6k3g
P5zfyPFgKR/3WIthDFtEa5PLgv0n/Ysbxz++t8GipRO19IZHArE/O8z8/R+joW9vZpcte9GKRGgP
U+a4gvpreTjH5wG9VjxE6DQ71gESfSdNSZu27tF51JH+049dbXvD67kJ4LFMR87xpA0KZBO10WXT
gJ472Hlya5GJvUvK/datsI/aR5mrbh6QCCt1QE4tmJRJggiojQ8j7tL169ErR1VMq1JIwhBThX/6
MyEFGIXC3oVDPW0W7vA3A3ZBKviX6TsjtoAlDtGckH4T8v1P7YQqyMT75KZHkNmRmxujrGi1k7UT
OFotSnbwGrNPL+uWZc4EsSArKk6kwz5lXkrEpWOJhrdxkQdcOzwHlYvfAfaplRNhywVl50f6j3Ic
J4irZsEQp314NHHAASMieaKx8hiaJmoap7vXT6pYJlJlLUZWvPvok1xWYveBHUVj3OXjpTuNHF2i
KhzA7wQnhfnVJCG8jNHc4cBeL+cu7neQL2Ah5zM+/sp053OpBOYsfFNKmiENjzgPcDJWuj4NZSQe
0bZhu+JCthjBWmoqy/6mtQBIv21/Ci4XmMom+UgN3EQp9u4RqC2XLDLilNIJvOTpjg+/IgUCvBWB
1cITh7+/p9qWmYdPY7aDS3+IilwQ3P7DiHdLWNQNQwc20coLc8V5wmuWbtFpNb8hmiNqJ8ck15eZ
76PMVgAgB4N1Dmvpe8tjc204EQgXDySiY4Eh/hK0aNEKqusiyDOXZJLrfsTngck9SbZwHm3THaQQ
PoQTDsK1Fj6dKj8PfOe/in5b6cUXOdzdea+EJfST6lnY0tz70nEv/jgAFAfg1b9qOQrX0wWOulBM
HtgOipix1RGJIZsUXUZVsqxb2nf5KCZiz4579vhxJ0t6PvhHBm5C4fi6aqbPImNkYNOocPLuoeFH
ebSWfpjcBY68uDQdiCVqj1wqhyAd4KDMx8UcQ5MUu6EqLawCSy+qoAfkrm4hBpBGMpcw/Nqtg6OL
aWvvG7bUE9pdO3GJTuAOMUmmKoYqLLDWclrFJUteSasBzIiZQ98UglfqxAh9aI7E5dJg0B1t+jPb
2qnJaql2rZWq/t2OwKmeo8djEE0b2+pJ3b8JiJLUgvS+I94zEIxl05RkcdJZhE5x+0VNKqb+5JVo
ZOzTrPWRESWabUOz7srVI+NMRvtWELqWfT20hkkOgKSsInHE1WXf5Y1kGypXVd/fs3mhtmI9smMV
jFk6YCrFiidGyl6vpm+rkf+HBafwnHJlxenQMMPPLX9E6+FeA6iH7oGFgnqCbrQHG+Yo0HZQwgLr
DxkOAaii3PWQltnk3qDwnxOYBqAcVxSdsAn8dL0wJL7Lkf0UuB6yuutOd0xf8C0nBD9uaRAR6wDV
jQsofyA0EIqxQVTZBxDvH6Qd5PcfhIn6jpZxXdidoEIksa2scnXapPm2spg8cKR52U/eR45VQpzO
mSu/gkY7d9PQ77d8xUOFXFf8JM1fdML98sdNgNz86AtN0ooZyxgvWsNKcktH6QHBwGkRppllZcjw
5FecFzOqhztQKWeRO28Rr023dCDAwhniZ7lTd4xADk3YepPERD6T2AebP5HZmIAxk873GYFS1rCV
4R+E02uwZk9zheY7eKBLbVTE3GOUs9purxt3akuZaxrEo/bo9V2xn38mOzXwzGhZBbO+DBCsFtvj
UoCt6v3NYmNX2qa6U2F8XIruBqN1vju/duGgt/Jl3YcCeuJ+/6Uj1u3pKfY00b+laDiTplvRJysB
k/JDfjkmP+vTSsJFbV47vF/y3mLTQ0E6+Zvz97K77HHmtP6FLHkdWpEqXqJy+FATmIrGhS+4rBBh
2teoUJv1Z5UYZ/UIVb3O02lDXounukgtNJUIvbEWsLZhZqd8C1o8go+0xTk2jOCEyzDuj8vYdmRY
H4U1CPUNFlBvVcq2JLG3N/egaNPMqTuJTIN2Tmd2zq3BAgZi/LJeFevDy0E+bWMl7q1VM7TTVh5p
n9/yYGc0SaUGZLH4tKNQR2XVf3yy+2s9aZ77HpLUJ+DyKc7fEvxGpAmEuS5wLw6NVCnlvAmlqlFT
veo/xUBzfPvugFUDqM82jKeSCD9M16MEfydf6a7xVFx3Rpwelc66XY12D0X3836AcTibvUgMSy6X
I4M6iU06UcTDwPVFSwXyxmdpdyjvvNNhJfY4OcRmmfObJoTUgR5Y+d6JhUyzcSHF5lPmMPadZHEs
laGHfDPW6As5O58AbepKcyFfZTyGC3MudLflu9+4gI4UEq/31aSPgwkmQmyJc+oeZyTXNc4AIgKv
kmbYSSIPv3iZJs6IBwQadMKU66p1KL6DSKXpLNWnReHR2exkl1qwdQYosNDkSG1IxzLW/itAXIGb
rJyiChOnKwrPs4EGfeV1b4VORzuNvrZEKha5q1Go+S4kt1igqKooSQBD8U+NCSA7P27WYG3KcOPQ
204AuCxovrvYRW39peD5BpOtn+wx8pyw2VsnqMu6Y1kpaTVv/qP7Q3HAZdOAxBYJBUufEMJAIH6i
jNF2m5tYSRBHWg1UGo1SekYV/B2RQ2BpgMPqnVcuVeqdut7VJnqsvqsfqPRQMM+c/4eohDu0kCIM
cuY2vIVNXZkDwK7yuSPyQf91IeLJLpF6RZ/r7cPM8eg6YxwnbFOSbY3MTWlUL+AwmRySJQjANsPB
OitCallKwHurGgfsSDO9hbpl8T0aXFFi6Pg+PGvUpFqB7D3LZG3gwlsfjBhjid+NEYvPGH5gAJZV
hKQX+QQDBYbJLkxXbF3Y/NuLZBwcToccmJ3wVkmUN2Rjo64kPeg3fGrMK36FyRHYrakIXnscBLAc
SHlM8IVL4fNglJf3Xab8hkY69JKBOKUw0EmRqjr9P/Tx6hjSnLAjdj6WVu5QHJEW8MuNSrRSC2CZ
i/JKS2SlUegbAIRZ1E3Znh/w9p3aUqdQbQOiW9bxtZmHb55kl5tdFgNiR95RKhmEuf7KkNEXpOFw
0E2g0qvTtfp49LpxvJ6/Cz9tvo59xRss1h3wKAv6HCUWvWZQr0I2uzYOy14F9hAzXoeqmMvESJDd
uIna5IxE9oIkggOylJxZ6hnxe0Iy+FHS8iEjlWqAMP0Gk9vxhihjvzdh1VeYBL2kyTknm9/tCf6w
pj8rIvjdOyEqvn+xErB0eG/V0Gp24Td/HKgnx60+1mlD/DLzeqf+9JfnsrpCBLJSbHGFlShLoIdA
2ne4xLPW+HBT9cr69W5/5OVEOQapgNqk5CRjaxxjRTnS3z3zFR8B2LGOIsk2FA5EVHPoOPA/m8mW
WdSWiewXL/STjLczNio2fAhXt9W9qVaIRd0ri9hFusAEZ2WVf/bHFvGwloDdJCJsj/eTnXO5bWPV
RrfTLXuB2mkBC5GpVDC+JOR8KqCBICDUOANdx+XFztCvk3Ai6rzsxZGEENjBpJ6zm+uQw0VbCYJs
ukML+tI81eD2BB7oEEAIQTo1uPhcEqUA1xoHth/1QJdX5chZfOXgGUWAQ+AnBWzLg5Zcd8VLTEHu
WICG8vwXukK57zsx/vngAZQUqCmLXxY6deoLTuwMzdUihGlKkxy/pgu0z7vc9XFWYipDcNs/JXHj
xE/J973EeV0vZpLx9OncFjBYxmQINwRFIQFEu6OM1FEQSRefqgjG2WvmzVSvf4/wChIOIwTEsnOz
PUNePewLBWGCzoK0TEIDy0B1cjmtmB44FgoOYwOAAGzllUpSOkt6wzQIUS/3dDhSusettZ0jNQ20
AuHNah+cCv/KWhenAf6LEd0RFKLw7DS51OYxYtmeopbB8u8BVJlCNqNgj7XwtyU5DtEsfiO9aoha
BlFoF0NTb0WBW7qpKKs5oebwJTaj57b5Q0XclV2NLxdh9hiTF0U3y4p0NBjHWUYPbhlYI9FcxAVh
RkKlbKzmJkvX+0e+0t3thrrD8aZgNyosSPSBdTiiTQmHZ5sHu+72En9gEPnwKIg0B7tqw7jTzdzy
9gp/sp4Q0ojtS9S+B3dDMxAbZiFUQ7RAYMiyDy8cMDMLTSyI4AooSRQiRSEAEToWfoXJT8ReylkN
9wvSn1W2NMyIRGVgQwNP1cz1u6rVbdOCd1xADXz/ivnmP6zRbleu9pHaCg4GMzeOyc9Sl4C3oJDO
7vuAQV/wItBIZ56YOV1ouHtW/ljPrzYxNSeMXO0L1kQd01UBlfeLzCpcsfMr3omZ2xdU7SIl+8w3
KynyhlWn9hxjnlnRIeyYJKzHFkgrGpCR/ct4hHAmNUtgRle8XL0w4de2JMiDfA4PDtHntTgdUP7t
hpatzIAIdgjmv0x8ek4JgGMgzlvpw50YTdSZkJNsT80NjK3SWuvPrs5jhO4U8Vbcp/zCp7hWKPaE
tnIRMVllwghdULSrsozejxBVyqv2GL3dQ3one8OlrlP0wCvpSjRgY3Z6yTGA0dkTG+PJQArZYBzH
T5n8sd/qTu03V/RmOK1H+tq5duu3douE3KCSCnaWNMHEhuPqLQgiHBC+bRbQ58E1Vu6oTYZu7Uoi
Sq2CqsghlBVrX8lOu6ixW7dW+3H7bTdYCSVlWKoSPElrJuKRlPeW3WlGtdw2AjU732jMWftFtPQ2
DBNOhU2QY7kBcFgM2+QxV6dQQaVklMZ0KhrCHqkpxuvQjhaRWt1/QLKq70hdDWipicmBNO5V5Xqm
gExZgkzOYShAlxwP3nOuNnAd0d7ZrhJtJ1kGJl7WloloChs25HTQzb2JJY1CTghX24OAUzH6oSOz
JJyoFThTZ4/HjN6alDeAJw7XwsV4Qk6/vNRNpPZfV8aUEDMkXCtWh/GuSN2RIWpfPcD4PhoaA97W
FEPHhSXyhv9XO5zaR1eJgPrQjzJs4t+XcgS4wnZGRSBnBjw2jFvwG7YAxh6dxznJ1cqRFcAMxFCM
4kapdXVRqja5C+5WAUIjcAKFKd1xVe3Rkth0FeCMnTMGws9Zd3FcGd3EzW7E8ZJ2FyfgK1lSdMwF
aAkROZJkkHflHI0GA8PVNFKB6bNPPaeP5osTG7kCJsL5WeVDKCFtlb49wFmG+j8NDY/Ik6ZTneOO
+jAUKdgfwRuwensEOJWSVskOPUrZyuO74cD//6LpAsWM0/UhIT4qqwwuIHYPJ1cHQL7Ka9qzFGvA
VRXgOlWI/Q+Lq9yzFvPCZ3BrBZbBHJh1O+x9jYwEzIRD62dMN8xBeoPtzOs8mVDp7NOU0SCCHeo1
GoF0fHPu13oYUh+szjDBDdo1wCuNj9iR7OPw3r1y1Sj4WQ3WeQYgsJxLdfMVHIsHlo8Oh7kp4tno
/UQCoYFfHFB1YHUrlazioeOir7j7x/s/0NuDJSZu3jXqzjhRM+5HwFzA9nSqEQzlIUUqV/vWnWh6
JFDOkznUhzOleZIpq6Fk3BYj0U3LcFI+9EB4CVM1+ewQOaoUjiI3JJR15db+GFg9DDEwOxXNlGCT
PEewBSwB8CCC2QQ3Ncsul9IRC7wDhMzC9rRPIsWwxkd4dxqUSfI5Nqrdv+98mp3TdfOc8BTmD5gs
xhOcsVJFxxgeXga+oKQfc8zbQygNQvjF8C73L3k3G5pLSo7qjtCseBlmeKuXFWAUmSeJaCMlp7VG
oNvfNwZHeJsAwb/Z23b1xBzjyZ1CpHeYQP7O//CTDhXyDTDVvtrF13mSH+iAYQV8wg5ryDNLdtQQ
IzkxgOwO57ego3rqNHM4CV3HzKrhZ5RHA3v6iFUvbxDCo1b4yeaUGAFc+GjvFTw3+jkZun2jCU7E
zJN6G1UZJEhPnwTG4bshoq0SeEatL4uSSUtFkWGXLxlbXzOjoJYTNUECtnB/ak+mKg67wtJq7pwi
sPGL2QBd5zPYigNX7Kk0opO0lOXnvOBPzCtTZR3Qh5Ma4g7jzY6Gl6+Y5I54Ac+oI3ydr54ZMj4C
Uxemr/rt2hV8yfLN5zODpyOeqexWVdMqYqS5aWMogUbIvI7HjKU/r5T0hcqE2RNWVOVUqW0qkgsa
MxvgX7YI/X2EKIQtmaBmD2dUUWfI2mcBqa2iTHfYYR8RaKpahTujYBBcjlDxdEuy/j1ZuSMazGQE
yhonQotIpBZ/oskyEIQSDGS3YOZANeDtImfuSh5Dc+8hVhmDBE5WjliPxoCJk9SH4gP2Yk5hVMwb
m1ZqUba5Mgf1XX4BVpJ1yQca2cZcZEysjGM27xGxfN9bSrq4c62N3ytVxcIYhAxBtZAnOTWYeUu5
gTtsP7V5X6R+5+rTTrXsN57Wi0QK1TsZL0iqOLHIjJX0HAbImsoMvUHW/BWI+sEhgutuBQiUZIgN
zd1bnG+eNE7QY9fQkiUm0yszqTEg00BDrYpp0xLbkTIEZdHGv2Umb/8S/VZTXZVmbwGIYx7SvIXX
H97YMgK9jL28BDypOo4xenUeK1+5WYoeJK0CNh4JZ/CVjcGi8XRL3dB5OV8MPvD1vOnQdm94AEf1
zk19DIJk5e9btIbH/OlrtwdNnLBq3gyUyGINEetK5a8S4el1bcTx0uQdPWrIc3bjw9Jxx5pyhx0S
hC03abicxcjYK3yjNY3M941/Z0QOjdvESmUvdoDdTp9HGWoX758BhEhTPgg7BvevQTiclbmgYH3H
Z8z4ZxAded1DlkRWb44XKM2puRWqRdffPNotTAgRaLWvahQ+kw+DsZfuqhuJM+Yx2RYDjoeaXbZU
V2SGuBj3q4wvBZNgGcOuJKcRX3a7mHMCUQQ4rGmJ68fiTEXoUHLPeqM2QkMeTpNoijaGXkBHTk3X
hMQaC1hgrE/MfTOfFY2VYzFK2DPFwmtpKJxVNcU0LUH93wWZT/dXkHv+w7ZrufY6Nae4H25rZCAs
NvWN/ozX3bQ4dgoxHP6xZT/lU3BrGoyE3W4HkSa2Gn10/FhCeWwKl6VgBXNHmu5NHlZtVypgW8Ea
YasdVxi/D0ek+FGs51hjTQCZluFlN3nH4qhW5y9J41H0wdOm5t/Wac9H9lyyzN1w3xobKhqARthP
7a3BAUPZGhPxfCQEVEiqKo+YO5/yEugTHAz1M2s2JMq5LNl8Brhd8giCV2SIz+v6xJ3BpHA1Ctr2
XqC3W2Xaze3JzV671gCYZxPygN2Gz8x5yuo3ct3NYg4boCthtqYTCXRtpT6P25DUxZOJr1eYK0jn
RQC3s7v0lnaKRl+QBvSxUh0yRJQ2MB+/JzRwlctocWnE9KmBZzrcNBjTo2u/ZdC2kyjmP00MmU4a
1ZhHDDxj0Ki6izSiTJSxg5zGq/AVRqV/dvr4+7p2PhQQ/mX74iIKVetQ3bKchHArubPlq5ir6lvE
sJvXpefUS24B6e6rnC3G7B1lDHdGluBWZTnt6eLA/KjoqDE0lTbIJcugVPg2+v77dT7qujDQlSVn
34PaQ0VbV0UmagwhYRAPmgI9TioAyIDkAOhFXd1DZznR5ARIl+JMJxyhDTQeVtjlmd2S+sZQ/0xk
VYpCj6Lc448H0zjbwspDGY1qnZDZHrGmvDI3y+aMMX30YaLuj/+vmbfzUmotP1kL12C3zwnh4PwR
8poJNYJwDF+WHUbWvXj9fgwO/DqGei71A8EcMPyXD1JuOGvYRBb7S/DqE+lkYyhNAvFf1Uz+o701
oAYgd19syTdcnzVSIm1uPN6iIsEfBdhZc49lWgqI6JuyU6y8P+2n7HzOnO/M11RurWmsHakyMilF
m9w5QnPeLdFvg/1f2hT0IbvTX0np82uU3VLKBIEiFG+oNd9WGswuvetkzH7XezMgYTffm75sud8J
QEnfj6o3q08JFAoyRJ+fQ/k3AH874cOdF49xgawp+iCb2m3srINWhIZMCvagceCJh3Zf/OPPFv3A
jxE3N6ThLRWFJAgU6dKdWfApj4i4bjCorxdjD2Nt4UNyzshPvrZ4p5KWIPBvMXOfltRzGuSjdVup
LXLW6Ic6X2zOUex6+N5+b/nzEHtiG0qOBGq2IFLm/7Da5hs8WZNe0f/7jGSchYnPAWYAq6bqABnZ
P8owCR6JgTdVymEUa6cuL5gCAVZGJ7jS77k5AAccX5urmjGsRsUI/EE+21Hp8StjgM9KtvJ6NOOq
gBysI/7nryoe8Kt5Z6gzAlxh5uUJaBw8qAyT8mhKY7w2aNaaWm8WxYuGK+Y6cpQSXkztmp0nXsd9
BNOOfSrNA3rgy8jUQj093MP+qW5bsZ0WyMbumfHzAs2y1GMDEEvxQVIISpQG3Zfwe6uxRlYkVt4D
MTPkewcSklW5F+Z2cXKv6yeOiiFmil0dg/oj2yLa5zIoypH6BoxVG7zpXxEeJEf4ZmFmX/uERxmc
/wv/M7sbsod/FnwsKFJfLSLrETo4oMrVnxJSfcj0DqdK53h/18/zDcjGIdq1+8BHmYddReeP7QDu
sUblisAg5EkxNkFczhSUBOj2YIm8DKc5GDSI45nZmz1f1XZhXTgPNs6Jmjz/wXO34Jy9J68P8qni
4nLHBaHKFcXgAPM4h/XXVZiMzQ6Q2GxzqP6pa198z/LDS+IaaBFfT8eFmYosVCgJ9q0cygrsedM8
uZDElCH55x33btglni4JZ4kC5BUoJcS7MjBJtl80wJjLIoLBMlH5U3OHff8i0svHGTDhp+iO6T1J
geGXEPgTkvUA66SSZm3uuagdDJuWZhYr3Spvad9yD2d1q3Y2h7eW08NqDKVn7Eex0HEk4no5z7Vn
m9i9uqvgo7/Xvj5xZLZ0JKfeEppgjlpKL9yTQPhhfvihqwUeJmXSrRClsHAwea7L4or7gmP94y1R
TViqMowYeJF2uquWOEinFWi6BGnPNYoq6uo9bxHpprW19ymgFSuHijGC/ukwiDUxYqHlPE6jYat7
X7SDDNhB1bzQN6NcArZrKwAV0XirtkrE7uiPAM/npw+5SEJVtj7Kn8tyUfsRYNc3OBNvm6HQqxgl
yYACVsDPXLvcg89CqrdeWSDzajsVdC9M88hzWgjLMS2PDXu91aoCKVq/E2PABcMqH5GqPVujC0Sz
OVNniUGSZGrIdkWg6zDI3mvh/UBjb6Ttw7b7xpAzOUL1MsVdJF+DDT5zBeEhWsYVdAxy2ewKGCql
YbUPt6nPFblEeqQhHbYRc4cEGNKtLT4uNzkwckHwTTBE0OC7rhQ7wjDJz/Xvz9yjhksojATswA6g
9ATe2kbldqjpPK12LrMrmbXqQ3PMHZsM1aUOq2LvenP7j/4OePjha42jx3N4SMPTVU1fd7fpWRN2
TePRSB8Wrzic+C78pM2YThMVTFJx4jZ/0i4GV+KB/qYGTfylTP+/JHmXbM/UaJ9rzbfVDstghOJG
evtUpQw6+HFg3G6OZeKF3oigVkhKpYAhye8z7BpL6xd2XsaK7a+Kbqv8/mJD8Dx/b6j+EwOnMj+U
7FNaLBjozM3/+Atp5Jp5uO37isCF3HDTKfoaX29X0YuMXeACrgnQpzzQdAGWufDdi9M2pQ0XgxQb
utxxf9DFXTLqcdsnhotilAIqRkA9pirijF8rhvwHVprdeainZOvEILWSjF1vTN62v5OSIO4SwCyC
MFRZiWrntHhDnrwbRSr3mrMgM39g2sp/YAXBHd7HvFMa+BAdhzHoA2bdO/vBPyaHAVfJYAEN6kCe
aVENn1dPOqzs96p00tEizy0lzDrep20M5qop3XOq5/gZbUi02iYyQUif3G9hZpKlj8wBAwWBhFNn
Q9iIidihZWHbtZtSk4e/4Z+b4TJqJmHtlmubkqmmV3JS5reP1Zr6VFV0jW16QAEja8jlLfd5qMPB
cQpF7jyaNwoAnOSA9R6Iu0WGBPs/Lo3PJ860oFiwTPt590KF/kgiuUQ8SJ7xVsNh/mxPZ7D0Cl90
nh4z9MLCjiFaQQ1v20ErUjnNgB9Fw76QdHGbJskqQxNpjchw29znzS+sjLPsKs5a9qhk3sqQMLOp
8yOK0JfuSEvosVim+yJ6EgnBoQIuHPHpmlLwS4QI4MlYp6RYR+LCKKi7tPQ6y2LPE5GgulTXEQ0+
9MoYgcoXayheFGLZGmiBPfGdan3/YF4yMz5TTSKSJuaaCYz7q1MCkBtKoRq0V7x4Vf9a3WsoQpVW
ZFZIkYXn+H6y/xv7RoA23wLY2gO3CtsYC4MrDSdXx0LOsL3iE+SGRnAfJ5JLVsK78NWR6MCcO+OZ
zRYAdJoYEJWJXl51p9wK47TVP7yhpHkV+wVTBbkL3A1ve+10pM4sQVDDNRNfbORV4F4SrCWu+lJe
XOo9bMjAg0Gqlj9hCK9onfEXzhZ3jbsSOSm8Gwk47N3EG4LxLsPI6cQuBAJ9s7A6DqFNUPyXchXR
wjXLw5uLeQbZ9q3px1OYZiYqUmAhfZf2XAmHCccCwSYlDBgvfq94kl6lmylMJnl95mATwr0apdNw
2kfidi+eRt9OUkYZ2sx9qCSghhZitSUoRzh3SB7d6jlWT11zVaC/XGkmHkQms5ZB2cduGpJxD+Ye
aYcrO0meWl9X5oenQOfWFvqRVRCuyoEKh2Q5t2XvKYj4K0FspC2C1WYFW2lLNuC3eHKt6+uw5xfr
Z0bZoDU13U68A2Qt0d1AIRPAfsp58DZ79MjWsj4JHwef2w/hIYHeGol6FAWAJSPY8DwRzBHhOTjm
y+7ezCX25UnAOGfEeOpy3MCbYS3gOsn5bbArHi3+Or/svy4dlrVtg6u8eV3SKwmEUfRQWxHnlUpP
wvmAwRQzL35SULc6ZP/yRk5NPfDAoyGwPOdC+GEjNCtY/Z90VgRWrBRHyx1T5UW9iZjVMlcUTVmO
BOY8W6moKFuojZ+Jk05MUHvlkpwvplXqL3D1DTjNqwI4pzq3FXboUNQ/ekytYTerUSLh+HboIbAD
r7/RuXJ+cdB5mCpwdqNYHWOW9dIofNxzSAlpvH0ZsOMb8soEA4j6itKcWkIEfZL/begavLei8Ylt
gf1njlSqSn1dGOhlV+5xC/egJWAzbJQN/X/1jXp43S3x1OAo437eEavcJ843hBI4KhPARMcUvZ/g
TN1vP7jXgpwcq1/WIqKK4Uj2SYs3p3Lcz4LyHHJym50RNsvFFEqSkXLz7hlmj2CWZlASKSNih/ZS
rDEizE9k5J8fJALQD4yGo84YzTqVAho9PUBhDjN7+c7znUCx4FGEVZuv9hIhZX1gJ2sBlJOU4Yfv
+tnXkwO1JQvEN191wKxCotDXn0Vm7aXSwFCpE+TsT4wBv6/TtP4ZeyM5ZnAUcYXUWSPqQEJ0GX/Z
uIJGxnm3J/Tnqb+Qqo8Jo8pgnXxKfQVVBbG+zQauD3fRC3t7LDUrcNMPUUxxAcrvrrTSjQxfv/wo
+r7KgOdKSg8UyXGy8RK1yDBptPYNM8waMTik11vMvZX6suQDEp0IthybRal6QNzsLuyLJkClcF9P
Q32TBql4XhIZcOuxRpKJ8fIUwy5DKshBMTImeUxM2q/T4BXD51Q+w3k6xf3JmzXfj7ewMj9MzJt/
JrfRAe8bCY7FRgrDtNltv0IpvwHP47VZ0T/NwjHKmmDfNEml16tANKPWxTzNI0YvZo3texVyEbbx
uBrP3GuTcb5uVGz2a4/gutGG1ZH6ga7KUKPLc2bu22HrHj2xIO75fDsM1lQgCxmo18H55zAr7xSS
UmWzW5jGgzvKVLCK8nufK1y7kE5c8Ry39WuANUP6sAyQLyZKskEakAZosX9LlQSZHfiQ5AvyvUuF
ucEJrxGJoNM1bz4j4L+vTvjcEsoCnLuuXIZ6q3upHFqtGPLEnT2ulQkd0w+4KE929ywlenQNldZI
SJOcuHlRehyVLlVCaGazgE4//L7aR/P7yROabpu2kLuQqSypNGcDwyNvYLiE0QOJSNv4I6xRj/ml
PaQjQ5xpvd2wNXIkSa2eWjQtFuoiKcjr0AZH64JMLlPeTeURMbeC7zVYmEiAMGK+sgE3+FZEFqdC
wQg+0NqKX+1ClQ9mgNlGd4vQ8Kss4YpCvzeT6ad/i9ttfWa7JEF9FT96Ovq0omhOVlPtjbgcV9S1
l/LfmIAGXupI/URBeZTTjLy5NYw+FBGTlnoV4FS7M5XKri8i8sgZqnUFQJojIe9Z5bWTi73+6ot8
iFzRmqxAOhqSrRzC27tTgdTYmqBKpjpQax1iKGfX99OgQtYWpUEGCkvICPHUBTDLU3vFuoPNZRoR
qcWtvJ3WwmCo9z0EoyvYBzxzVBVhPr3DLHBhkdE5bWR3wsIRQ3p5jyfm+nQ6daUTTjMn1JLDqc6Z
OJz1DWsYDgH9Ntg2yYIVJm80P3Mw40OxHu3QpLoIn5sYRAE/v38LPcrvCj+sJEW1+jg3K3zPYRO5
d4KqF32QtpvE/0JfZN7wQbCMeCOM+hBG9dBy8Iv6Cn8uxBWOYFpsfrMfhEEVjyH8jAr+NEdgLepQ
bYfl6F/AEt+KFe9H60U0Bf58FQcowZg/p+ammJx+hDJO1xvZftRuF2EuN0JmRryAqKCwRKw1Yh78
1EXouxQL2wwxAbA/CwGeS/dahs3yBbvU3ffs6JS774h0hSK3EXy7Hx++v8kvfrUixzLElZt6yqPN
gOegZHtFd6EpW5BC1HRZhqBbUc4WttzCWTlulnNtF5yVBoHtwYjumzKfFcn9Zxg8b21EJqiqu+Hg
WgFq+VNvRooE+renwELY+V5xnVsesXCA9I0cMh5IAGlWScqHk9GfkoZnd/X3/u2YG2RWpCLCrkOn
y4QgbOQzEha5f5hdIiNkkcJOjlKQTUSw62pOwFoO6I8D5ZAkjVBDPkHN64mEyk3ufR3AAqPz4sOT
2Yd4UAdxat2QLtKo/x5wdyYGEiu5duM9TRQmBpaGIzVuarNauG/vWgU0kVUJAGtHUcGUcIDvuUQR
QPCWYXrxeZzncvkGADem96rxyYuhbDjQChbW5pVh8olVR4Xp310vqIQqzKERODo1uWGR0ZrkUmaA
8gHtB9d3Yh6hg1DLpSp1PVveE7KrioM8JM4RfqvfbR/Lvzv1+LqvbKPmQ7o1xzhxFOsrzfI0Yxc7
w6qfKETsE7TmcOq+qylhWg1rVWK9W/fi+PHn/uW/GAx+qSLBB4sx7bADHfQCFXi5l9luj7GReXmc
yPqfPQaTS6kgQAhAcODou0HSp6ut6Niq7ZNsKAafMPfrFi7HhBU8xRFSBDKY3gIDeDpHumP1N1gY
7k3WA5BfQIS1I3g6qojeqVv8+7FAQkeY8OqrGm+ywSjX3gIkSwWHdCnI9gwV5GT7tLRG5VvNVM01
Ibwl4fF9RVVo2NDHn2YBfbUALIDrgT/0iKKcK/t2cevnZN/eJTHXAySYebbdw4yOz8jGGZvwRz+R
bXwo1hAKGvbOj2DlX4IncmjpT7vTSiT7qReqngTL0Ceq5likLlWqydW3+5bZfzzAaudkaDQiJnH6
8zyrk0XOI9mtQzupujsO/WQYdFOrQyoW9Q0F+pQfq0I3v1TcCi5nyj9kRhNxljytP9LZacQH8mLc
7mxHw9x6yAwyUDTBZkHKTRxTNrQTsXl1UOHDTXAg1C+YNdoLusUvqCu37oDpuXOl6Gc5vbhMqBK0
rM6HiFUu9B4QW18M12TiyrHfOI0zy/IsQHS9HV7CZXLirZE3Bz8duG7ifl84ob5PIl2fSMT+7BGo
HgBrWycC4pbqI8mPmMJORhUey8mgoEZBi4mJUqNhmYB6zlCPJuX/tZMlZXkqovxPu8Hj1JGk7Qcs
Q6Sivg3uAHJaK/OIpIRXUni2MGnpbO5vQeYYgDUxaMXtMI8c0tXDOgtrS7VnMIj5BBuzN0ZPa5ob
CtXsMmwcbr+20Yl3JA/3qsYnYZtbAiFC2iGFnH/dHnQI+zoCTVCXI5eGYr6HWuNxrvxGAfCs9pKx
JdfxR7vfcxE52qtwwqabDI083wtd0W9vJodv2ZRi0GCaB7UjBJMkQ6HlvPDopOMjbwUZIUM9LMId
u81Fp7S5MboBfFxZrAvDHCTTaL25BFILOtsUoCBcfOu+j6gtz+fvblHXzr3JOiNAORxSmYDfPVK8
MNjUaf69y7gJl54WTw27mxHM0ZODC0lK5I56EeFYj6ddT08PXBkG+DD0BgnYox197D+CS55qjWbd
5S0iPn2jHSB1ZEVXraXlnW/fSWQvGTUh6fHEUVwNsokxQp+5KP4FVe0VYn67V1zRYhEB18W38XIO
OKvYoH2x9W68WRoplL6WG5zstyUgsM1Zc4FRA8eGgQwye7IjDr3IDz+lqPG0B9vDPbyHYXQNcM+H
VA7RFgbIhiC6Tyleb7N3tXnM/6pIPXXZWSeDISRvTM//ETpBJM1VbjJ8/b1iO7tEugDIFJs3NuxR
7DNoMp2s7rduPwdTK8UQieAwnTBAI9AYyI/NgJIhmfsQEOgaj70vRwjXZbBPJECsaHaIFp2xWhcV
rF3ZhKVHgPApluK9VbFYRxBSnQkOVYEMDErfdC8v48g9Wz5B5p97vKxKxwigzvJi+a94jFYphIKp
mBORxweH39IFoGAF0y+LJCj5ayMvrRhw2vha9bxXAFwGj8jc/NWbemdP/bYTUU4wCOuzxKHPAVoI
x+5GVqLm7dMi8fQqsy3MLa1M4uiHDzMrIXzH0Ja8SXYgyJCgzj+CUy/PO2ccNESIuttdZTC0FlTg
DDY/2M01J91m1qxcHVt5NQwc7M2FKX7skyDS986LfrvQj7Cn81phC5L2+JuWADFpaGu99EkdqL8d
y33tbjhx6Dge2c5v/CwffEJovTEZcGs/wnlYoLdcPXa9YmBEN/2oo594ApaxRqgfYSiL2jGMQ37W
tBjZjzeh20hh2/yJcG+QGEfxTSmXt3LABGgEv6xwDllG5rSfFxDW04Ibeg75fPobmGzT0xQVKl5i
WXlghjlT/xoD19+AdZvah/fijwGdsrBfSMH/nc7HHip4iiC/D1MqwbHb18hMtiFfqBBQwCEhkpGM
PO04zvTotZ9W7HDbDfN7Lwm1rGfPgnDBPzkFRSY6kSnCIJt9oZQ+q8WupJG5OULjQwj1Hk8q5mQI
ameuSHPuYM6x7hDIZooOZ+JZZ1o7EV1C/GHku5QbGUtTJO43rcs51fOF8nDqQvKVmONvfkGBvN2W
64tYX1lCC7NBL/0oKJi9thDrdP/1jcsZnkVwentvUaUKg44JtvIE06z6p6zj9g3Wwxq5J9+edUBR
thYHb6QYXt9WrliHifgd+/P1rc3zqR5Pa05tRFCenB8cOOj0R4ZxzKTdHp9++EkZNucQ9w1P9/cc
qVWi+XqUS3KaedMqpgWd3LVQvLsvHOMATOblD4sQGr/Pp6rmfCIgP7lHR0ktr0gTCNXD0n05LJ9H
AYdhAX+5dKNBf2r5gRXQJes1k9M7Lz9ROx8a0CrfQLWUBKOXA5Rkk5Lhhi0vWAxn6qElmw5bUyqj
AsSqgmPf/pNi1OO7THdjtFFu+GXw6dS475Ex4IHRShZTtyKdTqMG8ttRfti2tcKTdo+1N4IPGbSU
9jQodv/gJShe97v5W09Kh9HL0+/zD0Q2gFL0JDc+66CsJ8lLwFhCYA12Qf6hsaVU6uLlLFo2NKvW
l5k1x9GQPrKe/WVAus/J3HesjQ/IGYOYx4N3VXdWQ4I0FMCt+7UJa4KC0D+Y+JzWeX9XHANzOHj4
rDdXY+aiLDRL6U1ekgFoxCkZzAVcDdxRYbS7Z1ANl6CmbRtTOgEiYqRC6HdQIe2KvwY0ADsMJPgN
bUK14xUDdFUY+qCcB1g3CxJPdfy2syzDDfDDATwQsmVXJNCDrTJ9by43SCINA+0qVhuHO3Id4qbm
eOp+zWdD5C7gf4EiV++gdR3kQanUN3jGCr6WGpNW7I33DtO7As8f3G1hWFyuSJgXpDdE9YO7ggS2
whp8JUXoI/DF3lc4McI34O1c1Rol8n9Vd3AqHfzDnh6PtHLsCZ68iNHvet6V9n66OmLZN9o0eMlZ
ULq+OO2721SnO3ieRq0VDbdFdsMvAi36kPkWGyTOiHofiuagaNH27m+9qyMTk95NY5p/7SIbUJ4f
IBEmKS6fpRZNA0p9tk4HlwMi9pFSynY0HgKKta0loU0ZF29+kn+QKLYvrINDDpXWGb5oHw57hkG0
XKB0LHKJAL2YJilw5tKf2SOlVNMuoemftxhKA4jrmULW6m1EIFkjY2iLOw5qGDGfQeKctx3Y0i6p
Q0vuRy5fTpaF5jRFyaeaWEeri5jmE7a5BlWc58FhM1cgPk+yZqptmUcQhOPCJ7HVsORHDEz0h31V
Pvziz+tW55VjurAwChPGaeCMOhrUMhIHOsWto/2i5PiongXlcVUxb/WhN4BbsfId8+hkAmncy389
aEQD3bbX7qlfRZ+QAL0iSFLukh8ASbgXBVFMW3NcrDKxMnBrQbvkjT3yuPjUrnDkorjipHd6Xdpq
8d4tzkB5ZYO+ErSSVhKxYm7lJtsYPyu5v7YIP0OycYgDoo8G+fw9akGs+jKGcDschidzxOgeGu+u
2W3zLPTNbbtGJU6csoBn9lwpjdhF9oggvdwrfyPelQEWWb4mcInmiXdYItkY1GYxRXqY+/eahRic
NKvMzuDDmPU5mMtfehsVTCVG6C1mrSdTe6zKu5rw3+TEErXwK/Vg/3Ut2RRsSRlzlPZk5MfnlBsP
avmN/S3UpmHUEHpFwfgicJuYyGz+2keC5nhC38pqeqNltnWcg1xQAPeFpNBRaohA3RFPNIYka/o8
StaLn5fVULbKbnIIOeTkOR+Y9Qjw/G9x4Qeq4b5uwGyMmCQXRs1pyee51E/2hDrIcOUQMziup91i
NnhfM6eBnBWAkmJxc7NHrJZgpHrQoPChzWQZ7NXXl7/ESeRPYhfpNcQeQXs7zaJfI88cs2jXmFbA
nfpb3kIwL9hu5M+LtvNpsfwOQI2jCil47EeTn2wFwdrJyDJvwMfRM578styvSkrLSg5TTcN9LFTG
d4G2jyLXaIwl1cCShpTeqMTU2eCmkPoYogSx9rkn0QY73f46xB2m00eCAljAuG+n+ynI8PMFZDlA
6xFEru2taT0+qNwlhLk/+hwI8g7jhvJ8LBvRwS2f1hKX8VBNze5E32YWNjdtWyHEBt0z4mL7Ngc7
s+dYmcm0ye4cGMzFVy+2KNQArqKMeNxkyzFvt9bGiL24KN51rVkIKFYaqYPpyQTzBGnZfn/9ejy2
u9XF1FFtVSLQlmemuNj1MlJP2iKmDrVgioygdINEW0kP3wV2UjlAOMYR2G/R8KF73aXW5uhiAsaZ
DrJenWx+ygrLc1+QLHrwbnnEzTcy3xvzh0yijD0okN0ey4nYzgSuYaF2bf87pSLwXFvzNmnlfTrb
Q/Ff2qwUIZjAJf5VgzGryY5QZNDkcWplaIEk9gjmKNSwLCTAtZeDN2bhYXEEoQl/JJrBBo0eRZqJ
JCc/h1hxdpWRqIDOmREN6p7SbDJ/G+BjUFrLBtld2AdcXOwrYqgsg1AVgdes9KtEy9chYdj2jfpR
SSXKXH/O6Hm+GVK72yyoY+31EzIKXh8kH+NRJsYB8SRny7qQUeCakYrsHzekSb1lC0GZWoLIp0IW
2rxBgcZYXyMNldYh5N8xpljhB0awG/tN/zZCIKsOmnLfVjax3N7FWHr0A/N7ftvhuYz28GzJiTas
aRKEV+wnoeuQK/EjNZvCsUzIVBKbyEz2+XwGDcke/MYwe2xY5fJpFvG5TfW1o2KYMjxn4mtv0gaZ
y4OtYBa5mN/Wws8GOfa9FJ/64SVgWxLVCsyKL4zmiCy53pSAXLcko6smOCEouAQ/Roodq55g+Pjl
GlacxtoVV+FLHUP/yIZr8v+hhPyyR7WuXiylt2ee1VbDYQ+moG01amerMtzOVc7rIaoLBJPiv/rI
F5VNFBorQc1Nz4bhMmZSIjPe2ss7xBMBld+AoNL1kRCl0M755RhUcJ5OsSLVlcHPFy35vogkIFny
VRVCrOStZwh5nYXBBIgsWeRhaP5sRfJlWFapRfh8UN9zyjfmBaV2dLV0IeLvNFr9uouW6/Xad8/h
FTsvBvGcDpUTgMBoJ7NkLspGP1PeuxSJsAeduehHj4x+UbTBJjxhDS86Q/uSal0lD3l2Ahbd4nG6
ev+udpp78aYYCXcaKAVbHFOPhbc9MffbCUbFSdiohgq6efW62j0nwEf+PDTouAqodnB+/vvKQ2Lm
c6GcGk+vgNEJJaNIjFHjE9rZy/lHSrUDtudfqcOe7ecjWDhwQtu0FiU/dgTIpXIR16bs15jc2k1z
uuKFcVzIe5MI3F+kd52jcgE9wGS/S9ECqTTO+lZESWRugCrc68EQKn7tacU/aSzh4jVuJ3lfokUX
gCdLoZ3nyPgMT3UzCp+F6Nn0/6zu3IWBp2ulXe4Ovbx/w1KEhQqZDeMB83WGAYf6nADPW/yiVxOT
AFT5cQcLKEMIRnnRY03R4kwwtiwBvPI4UMlffgj19zlWZm9/NrRIQoWSVAZHyTpfKJSRr5mbCfQC
Xy7Do3SwO5p/GJSO7IbcM1zsM79KzZrgBd7tUrpnomzlfCYeUFtuN1vNfLt14uQoNG0OnOsIVcJh
tmEmAKjcWjZCaJky7Tp59vSQmSnUa00cyVtvrdWFVHIlLglSasqMnggbqsvGnIvNM2BV7EwxN0Ql
xJZhOfBXnROTEU7WSYa40E820Q3T7YGIhPIkpcHJZpJRx2BUvKnGoRpXuK9LqwFHR9hgi5UotPpa
VjMstDY09RoekOWKZ6WbPF3wnEW9AxrCKxxcLLTDI3MPiVexGHQLSTydWjC/k6yihizWtdj/Jdu0
Gl71hfzGJf6JhmqLPmQKOrSXGpm6JbtF/C5mHb96PFPWO3Z38iL75elWG9OD/RZkpzB/JztvT/yY
MAhMcNVPxyKdjxnxUpEt+dSOntLf9sHeaM3bSj1v+fTHmIDMAnfsLzr3+CKHilAwdlWbj3f4RHPA
ryZ4RborzVqoMc4CXY4MRYid8e0AjiX34G/9AYKHnJlearqrSQ6Nad9j81RjrcCF/6PQ4YcWx6Ww
Qnfwhc5C/AYJiZ4LREVK4SI9Ffv/R1hzEA7ehPGzsrXVxOMJmXimHwvQkkiyO0BA0W3ZXexz9e1q
5uEYKev4RAtgTnzHrDHWqcSS9I8TJGHyEaZtHm0rAe+mmiEiM3koezbLO1WRDrtrEJgDRtbokoFn
0y6O8nfzRWZkZtY4GsHs9Jb9+DN859cfbJpEyltVbaOcuHwfUwNXNG1JpjjDzaF2BhdutTWx27ok
flHqzpRoliTH6jRl93vk/xFVKBhr5alSiN04j/kejaiKEU5YxGaIc5wEiKR2jlpF64tGL/Zk3uoE
DLfiwxRE9OxsqczWH3NyGj0MsRxUqsKeilbcyxAimMa2OTphaCt3DmwdRVIeTovPC3KIXguvJQ2U
Mp8Ar6S4ZapJ3Ez+gBxl8Eei/DDR+00IVFSue55mSlfzjbC4uJpWeELahEAgrNDFIKbZraTWuVUh
mc1eFzcqkgD+XssX79b+bIyiFR4xTL/SWNU+MNu57k93laRk3Q9S7naKofa8yU0yNLxMZiK2EH+3
9bTYpT28BInh0mkSJ21HutHzQo+w6Pv9Y8/LArHeIUqFRTRk+/fQXzL2Gd3NjrmcTeZSJSKOWml1
UsNjm6jwFSUVwjgdXjr0psk8cyPTOKYy9NG2T1IWRtkB41q9cxZjWZBwc0+b4wH5oB2qTfM6BQtE
vebHJX2cuxRSt4VpsrgRq/1N8Xq6H1iGUPiB9CN2XsLGY1pSlbctURZvsCTWhhunoau05G7JHiV2
/v/gOQlLW6xEqa6W/tWbE+w1nb6Yzop+tGGBy77GZazDs+srxCTV4zanioTNYaSshSiwt2b7/A9v
nU46qO9DPWubX6aPAfMIcCNczef6qy2puGpnmkHy7OFumvLMXDO4NbG/xNo0Wha0GdMlZL3yRw87
RrpUae+9RrVCuY2ZKyP/Zj+JFcAcz2/BZ02FGMCT+aN3uqpjP+Y5agc82qEJcy08ayiPLEzaNnxs
WPTNaHR/GPC0nZJQNTzXRI399DPZ1kgVFck2+LWj2NlhrI2i4+jlRW9jubQz0qFYGOA8OkLohYNP
VZ5/qQHxLDvKVgTUjuIqVpQ+/aXNg4liaIPp47P01szimS0L+7AV2gwIa2t5chO1KhrylPjSdtVe
HSHcdKTcap+DSw02+ef7NGX0sndJpO5W0sclTZWpyTJJCeSTYyWP+/mH1irWGMk7S0+toi/x3ecE
Jp4kyptA/gtw+Rs39bSCgUGCWk4Uw3ZCSUB93WDtVF+VM63Uuw4bsNk8/5rKmBKBsZMbYYgXlEDf
L//NglmCJ/erUWI9eFMIDEBUMQYX/OP/4HC0La81wivWhmlEvlu9zfUPCJ0uzE4KfAOHD8Twa7lQ
yUktseLVrjdVm4iBG5HFzaSXxIp+Vp7vMr7MsjoUt/YQascPU4udNhO+XafAuhghb92YP5G5lhjS
Lsx4OH1m9PD7a9Y1GAIa3XsYWVHUqKM3Z66gOO43ovkwSU9F1QVeD6P72e12Gdds8IxGp/3RxF6A
mWc+2G3BE6lYvay7POsjWooHcNnFRj7IqxiS0uAOjP9euquZxDtaeD0yB5o5lW3eO4G0F++8AsJU
pGE4lw0Y/gvfccqonGHhc+hw4o+YEIjxpWJYb5GeBit/Z/DrawUJsmz4h6Q+akF6GXEXke5Lll9r
a1xFDbR96kIbGIzsINd4qMoz3GgDsaSFfiCvBneIfPn+3qoP8AdgeBYloqod/lbCgcYz60wCggEz
g03YdFnXWNG60neX+NK6HMMk6nQxfSSS+6mXRAmSAC4Q69iqcRPCFWAi531TAobfhy/LgxwOo8G8
G2JKMdLJmiO3PmeNXzBFhQijZKoglN5J2C0VgusWs5ZboaVHRRCUE334gAy4adK9Hryl4WrxOhcj
ZcD/U73SY3iq+/yPGRftqBfjjt7vsOJvOED+bAN7Ralq2vIvgZwrU4jLfTy+7Nz5+j5eB9AYga74
LDADYzDpJSVdyl9+89AHDP2C2Be8LVnxRSTcGn28ZrmmeenHE/VPDJhRfD4XjRAPiFhDj+IGGefj
T2o5B7b19RnBmg15SnYizUCOi6PtRjyByACSY/XlJZY3TNMmDBPF8tSDjSFRmIDcKKjizIeHI51n
R2Aw/yndw7z40KorWZD5D4AB9OMRQb4zRZvjhSratwm1uUULRcGpDhZkU4TUO6czJLhHtdROtB5S
E2djmHDsUTiYK0URI3COihcT9OwnFnWp3lsIQe7WIkTQ5dbZ7LyV9xuipU+fjnWovr2Fx7xCreEg
5TItErlrin2taSIQlu5TnkcHYoj4vuC0UThJVc/bKC/TjJwOmNSbzdbj3zRPK2iddsBHpwV5LL6x
vhmwXfYnKs50hS8TOfhIwkopHbTHSUaqPYnfb2c9+6igbSsb7nWfMTegDn9y2nI0Aq1dvwp4EUD8
4I+BTc0RfcNCBkJF4fwAEc+s9uPj+CVZd0J5PUapzVqh87HgRoM2R6efqCd3P+T+f0gHlLk1IGd2
AFq4SFUVv9nSzFemBV/hT5a71Y59rqJQPqGvY4ncGf1ViwJUhnBtIDbZ1ABTLoyUE8SP06Ewx/eU
AbD64fLPjSL6/bqxa6gl7piglrPQ0bKmVBWA669DDMFupEWog95r9mj5FADEcOi7D/ADkH6spAqE
is9yU1oJBMObZO8Gk4cLRlOPph03S6zXuUIEqQmYUd+h+TUcJHkT1wZLpxb4W+1baqqbXGiFSf6T
hiFD9+11iFFSimWQRsmfQ7XxeZYqFe2k3Ri7Xm9VYhJnZRXE3moAdzDXWHmACpa6h1H6oRpAjwFA
o+CwFuvJBM1lFrSyWX5TG7/eurz89MS/cou4mLG71qcNx38vssAJb+nSFBLyiG55bYlfTucP6XBi
4ji06RXiUOKfCLYX6dukMOcohKvJTHJt/lklGA48irT7NJ6qzzZfmTvdW/Hc9CMzdmp3SZenA15f
Cl/vY6sBhz3yTgVWb/vgzMV07LVdhwz8LpxojlMavpVCLJpnMTDOBq7+UDhqH9IUiHJZNs6vitFB
357mlaSK8U2oOHNQxKNfV9pwPa1R8VD2x78a0cMTnTbOYhkBq3Ha7eWO3dtvhR97GPAcsVIs6Kba
F+WFMhhQ7WDrtIk3y6GwqvEIZS9ISqQJP26rSiXimhggnzelQOJtmOJlpshHx5bC6EyAECvGJLWT
L8hn7Qf0ZkHympKaxIslJN7mCJyTLcZ1pw0u5+w6uJgwEqAfPC2zfR5197T7gGDh0ol9NkxULpb/
K2dA+2aQV8fvmmbYyovnxX1FeMmkDWDLHIT5PEeXHEKi/6PTrhbx3dweSWnTleyaIvU46oXps58j
gRfGMZTicn6qnQt0OUu2P796KMfEqy0AwdR3Qw4yzsO83I+bIU4LPYTj0doPBnlqPYATrxxizO8i
EOFH5m6O84634Z4K+qbBjP4y2k5152FAmau5VBxh9WIKslON1IZhWDkn+5C8AKwqPs6yhZBKoTMT
W9xQddfpZMAurMUq2sWcyTucR3965Xnu7E9tLrQKkH/0bH7CvfBLxJSwVxbxJm5yUeTDnPSm7Fdp
8xtvZGvAxppNEKXUhrUaRa8xnG6r7OmNxwGQjjxLUQgISSLmX/Vuv+95SBgExfInFZ4njm2lu/TQ
99sYBhbsN61B7aUIiKTsYUGMQFhe7T4hYKtRKTDAxvWj1eriXKW4rH7eArF9goUsUJnyjPZBzWV5
E+hD4wQLBRouSa8SXua4qMSx4po4WrNWC9D+8LXKzFQSSIwqlgMVBwxQ+m170ozbHla4K3pDLTAN
9CKOzeNGi8NnCb5Rx2K5YzDjIbW5dYWeQdOt8Z7gCrIFJXuXlVBC5oL6cJzdBK+Gf7oyFua+WZ00
JfUjOR04FaI+F3vY0My+31LmuY65lakDSfXidcr6zll2wMiHXMroGTwuWSL3BRYztmy7iB2dro7K
vYKKBgAmOFIXd9ZWmIf4v9ITZl0pdlVDIzGixZzq/UbZ7gJOJcChVXjcXFC2L0p/0sks1CEXlWff
41FzANBE7BIcdvOFwjLn/vJXEgzy96d/Ft26pjiMKUtqHRblsZ2iqrW+1/s/fCdM+qDb26D8Il73
xdCZNK8rlcyhdGGyq2i63HVkESzB524oK6uqsy4CT7+L8TwLHPLpUKCqxx6eqgaoyk8qf17HLkfB
VU8FdBdqRrn/FaTjsnmd6Ykn/IQKQL3f0rw3xGKqmFJrA33ZpRr5x/m+jN539iR7P4GqOniZA4gP
2MY0kihl+Hl3eYUckXXG+Pi9eNFWaFFdwx32uX+uKJWwWFWCI34/eQL5KCRkZ7efENYL3PgAtOYX
Ut7Uw5O1BJlLcfhM74ftAlM7Y1PlzWOWxL/E8UQG3AD9HFp5NGLySOvo1VoLik1rXkZWJHFxSTZ/
8d6wZ62i+AZX+IRos5V3pDZKOnGHwkhvcFn2SjXkukmJeI3663EOrkYfJONQCUtHpWG2Y9jUGDBS
wIC73o0nN246mC+MXt1fphVP+fBcjxnDmxnRHHU2qMeuDuNMKoAO/goDmF9CdwvBLp0r5uCvINY2
vemODi2XxV5Pf74Ozf4rQBU5E2uE5DpncCi+ohvmxsTpVcyGiIfKOTPejom7JElPNaHXXDtuJWJH
W7xmzUeH+4oMj8ixVRjL2xpb+kSEYM21CuV8CF8qzZZs5/MSl6GF3UsB7F1Y/0l9wLb38MaaGXKY
vj8pjpkpbUKhQdPKisfttB34P+xrt1QyWMFb43FD/jzLcl6Uy7ow4myqEtxbFOx17IlH5+39f/FD
fcphhuYrpIBEcqcsDT7b38K8mEl+Cin2TOqvXY06b9PHhtYwNf9HBcH1ULVClpj3L/kBjzE+iyVv
5z2RgVLkSzn7fjZPHa6fL61GD3dPySkkweN2aTYI9+HdM0xRmDrugpTA4IPC1+rS6uTUcL0qhxSE
t/qYvWF+OGNf2bXW8t5jumSuiJlSNMqlNFMaFtG8yToFxhRWQ+UGoFwWUqWgnOmhMyOJYvAEd5IB
Q0jdEQM84zW+cYHetcFiossyl7ZsadSAVqjAqiVRd34kY2Kol+gzYZAjlhhO2ZOTp9pKJGlXNL2p
NNw5jQXL4+tyYyoVv736dhYK55ASWb76k3NBLyUUz9GQVmyjf/UAGRh6cOCIKf1Q8FrO9dWcg3n6
n8rc3NS34aU4kaCzY8qrZOMbSQwo20qKzwUiU+ld/xqFwgDdyI0XebZn1KuY7fzaDkPY/YRSuxUM
IvA5qA6r0X2QqiSPDFAwsa3QE/cpcoUOTaE7rUHXCBgCsChnSN1uyf0ewHvWlMhdJLmBgp44pabi
cl5WGkCZXFuImdOLnPL4ORy4E7eDcYJ+ksR53XwZUOMW+NkFi+6VrRuBP+h46D+Tppy7bc6a7kfk
reZdwWq2lY+CX7bbJlwb2NZyNUC8IMR3Rs75GNi7Spl7ov+IbSQx9LgiMr9S8cmK6oHzQZIJtr2j
wd1N36Hn39PUiNQttz3MFHOVoEyLY5kQnnLidxeMJeW0iSbvJJJKW+vGdVmSCrc4YfiiBz1Y2Tf2
4I3qt5fU/QoCoU6tgHxBDYQZHj7rvobP6Y3EWbFs0+jX1yBuG/HpTSdYa29j3Vtilu9yHIxATlYG
Cy4j7MP2hkbiSFeYh39o623bqVmqxm3VzM1rV2hmpk32yiZo8A96mUZtHuIk6GU3I3EO8UMPEPwU
UFapx29GJe45BE9LkGbZWGa49ESJmOo5KZ8c7G2jfgdSeV9aKCXnoe7yL/a5WLNFMzOzOp1cr2D1
Cdd0rThq/DK3coTZEHYvYykgEVV8U91VhXML3THr4pX4xVtf8pY6/fZZQfkug4Txc5UUrUUZ8AEt
VsRILP2HFqkdj5aFQNGdvEtLA5JvCECIHHzGB5CYj54iYaDUIZzH2f1lFSruXBuLXAS8mYdw1Dlm
h2As4OArfnYygXyMTxwnIJQz1NEW4QKNS76xVPj++FMaNWkqE2Ur1gtMVjnxWMKcmKzRXkONMZ6E
ZQyAJddlhERKI6Dr2FdcqF/EIByKGXsKvBG8yLMjW2VVNhnp8XBmB5IHb+tW0y19ukppby7Xn+g+
1cXoiw6ue8Y9ghB/DVMBums0sHbuj82MyWMA72bu21oJLdTGL2H89TeeT6X+TeJfqDVVw4A+CFTR
LYaJ8hHnAuAonJ6ocHeIkr9jA0Zte+b4ChtzMn3NWNvcK3vIaJ+juWM7pQGEsjV6k6jiRHiVl0MY
BX04oa3jZ1E+DRr8xuOdvgwVoL5VrTFm38NY+3VgaL5c/JHs/4+dUQ47MLhU6IUV5KNjPvgsWg2g
i7kE3aoY/8cHxeKX6CxhK0LuIpV3epNyQgTK3Wp6AgWFMLUoDyB0dKlAOTcubdpdM8xP5Nu1267f
/FLXtiOdefdglZB83xBjhQ7hIFn6/mbFwAasJhD4jpxjYUr71Tc8mJ6vVMJbhMXGTYw0ZIzbUwFw
Q/BK7UaM1F+TGwZMfcZnaLeEWJaruppQDtyfdJrYt2IyP1BWH+kssRaWSwziRqk2axwipFuzOAW7
9arYFFGgBsCh7GXV+HZbDD+qPakrpnHfBBYCL0zK3wc2OMB9IypRGQvkf4n3wXvpSXlAdb84y48I
vbcAD1cW6pspFCvIy//8DbgXumvA6GmVQQCDCJry5b12QVUKeUHaVVcVbmE2q2bJ5rE6EEDDYkI8
lCTo4f4X+8pk0cGQFW/dOgwaUBY4fJdTtFyTL1LijnISlozp3SXfgRZf1yTxAwr16GE5Hkkinjlr
+bgNwzE6SzGCFRsummqNdDgCLiR0fxn00IWzczYkvTY1J/2WSpXZKLsB0XrYZSc4xOatq83YwLYz
zuomo6Ep+2SF66VNex4OFQ92NKmIACK6rgXtdoHQuEsYl1RwlWRw35NB2BHpnxaiEkhgd1i4Wqpw
KX8dGYb4eD2CPbeOsy/UIn8xSYDYldfV4/cx3GRpjgknTwdZ5K0N/5sH9za3vDq/U38sWi8LOWce
kUa+DQm4Qt5DiAVxWtgNBxqg/tw2pp9hwROOORezuan9RYKhGyFUjxwvcKTvdbHgDG4p5DDslHsw
dvLR7I7p+3bVPtsuotXnOLqHaspTGb+ANrM58x+nmVAXxH9ePwwlXzcakVyiH8mfODPHiw+xftEl
plJjNkgbZoMGt/txqkS2wXB8RNoyme0KiTM4sjrj0PN5BYaYFDgU1wJ7ZKMwKZP7ET9wGsaZHipn
NaqwMhgHUY6rcBZ1SOXvWABepYMV/p3J6fbyuvQLSghGJ9MKbr8MxzAEyzbT2twMXljys4a82vSY
dmQLh4NrITLkrqmuTjTbiHIK7WZ5i3kaqu7Ib6dGIRt3B1Bl2Neuvl8S4942B+7ME83VbGmaWQ0G
u+5sXxzMTR081wi0X3hRDnM5BXcygYQuOJvkyjVS6BVtVwybR7LY+DnffaADMATY8+Yi/tAXiOOG
01K8warmNhmAmv4gTiRbkxVrrtURgqRqkf8Gw2no2oldU+3Y/lNDmGJq8jMldXxYRhXO5kPp0yWn
gqdryi6OgZaHUFLkcfx2H6PaF0EK4ejaYYS63r9UExBC2m8IodSKu/cJu4YEE2va0+lB+dN0n2op
4Cvh4pvsaOiFusX3hrnJO+bRPt3Kjo4MOtyHXxYs+aVRk+ucur2PPLBgEtoq1/fI8qckFO6PeHp+
1/pmK60k2x/C/mI44HuVjKb4RslpZuUJgbZAfsHiyStRhQ/n/CuP5CiB5pODikAZiJIaFgpLyTlx
hwLXnpjQ2kEWaTYppWLrUeaTyU0z5uR/pTjjKNFZPBgStemrA23bMlaB9UhVYISvJweWeiWu1TvN
nZEO9S2LleybHiD7qlw4arwEnHJmDTY1BOzzgKxPsAQ/vZ8KrREamEO4XLkpLxWDaehWovmoclab
sxwAlOmD3SwUshtPtp1rOm35LxKF0zf9JhxS3XDeYEM54y8BW7XyIhYU7ie4mjgnMQhEYj/1hZ8f
mdfW8B9gYqjDoT79vB22Y7IRR2MtUR/5vH/d7ju/wVspfqVZhxfnQp8Z1RZ0uy6JywW2CeNLbdOJ
HczITj8S2lBHR13XHvaZwEp+uMNrWWXZkKZgdYZDjvCv8DWmnNHBQZshkC1bCignSYpQOiW/bxLZ
1OHisF4ZX8gKgm5Lp5qraKPyPV4lh43y5LnRQjc6TzQNOCadm7ixYjKCgFoL3fH6cC62TOjbL1k+
dv1xu+Fv222we2AZXg2qQ4wry8lV3dPVl7RuHavWDg5tBe3l2fk+fhdjMJlOsAFyrZFu/hiLWKpR
DDlQProFPuuFoL2DchVoGj/GALYo8jTISy43xYNW6C8M2pE3fgDNk53jTa6zsambiGcCgqtWsHgQ
8DtSeL5tv8ooBOsOB++YdnkHNTuow2tzFwnQkD12NkNn9xXMdAiltqjlvn8il/DwEhVSwIw2j940
/6mtqjfmm5FfAVKbnMMGgSzoeIyuQrSqxmEfU11B0zg4UFPfz7rr/uuy/VLAgkSPdA0t0HXf5hl+
ZVSSQ7oBI0b1Y0bL4DTjGsWXBVSK4Rmu87JMD0GArAZQ9Kr7HDng+Tc5TypP7bxRfcXcHcr8XKvU
WqbwAuonwkO0A3V1HEtakYwX8r0PYmQhVrvKlMpJQOMfIsgzbCdYNk+jdQAI2CK14kzASPzUwvvg
2t5iSoYuplT1LA3aHtox8qna8yGHwh3haNn7DulZYpp66tWWHuDPK1hmxtICyguDy3rHl2SWQkvz
1r2JHH9L/cSiev3bypoYAHjeKn24a3vPnlEadaLoXqMq9/c2jQlC6v6sWCUFNnUB1b4ARPnvtmJu
lE8sPD6G/Kl0lPC85WR7y/aZuA636cWHHv7vuF0yZzsmYI08VZVn7t8SrLRxRHesrSXBtylHjMrw
DbOlFC5Tlh7fLVa7ltfElgAbCoVS5Eos3NoRqjGxJLd5eaj879sHkHiNrxOTyrVOk4cVZPiFiFUc
go5x/neAQYs0nod9K4v2Gh/TnKPrOgpGPmC/6CwOXHcRtjqxJeTFIVRY3vIi/zurrYSjnaSGs9mN
0BexOwjWSVUvFTfQyhkgD0X+70KqjLAzR7mhYsSoQCZd6KjlAu/yLFQ/7Qfe24tFrkrkPJoajwwG
BiWDN4VjyDD8NK4WlS2vhHgA1Db8jVLPblDdOI/mtZf5din9TtPPM3wzR88hmG7Aqdkb9JeqYe/r
z9x8yYGbVMu7HBgbQx/ogbzK3hrnjHjnNevC53nlPADicH5ZtafCX2JK+ISytshoUSvbMSekWr3G
Qx1qgt4ovIwd1WvcI0Pl3iHCOZ6Go1lOZwO3TC3e0uU8KOP3YBMXENM8dHf4iuXDZuOsq5jh4kxp
Hl5kXmhiGEDba9hBUDsAk7UUPAVLdx5I93F5I1XN8y7ZK9ZDapPe+1G4sdob4vwwDnsQPhQQflgQ
FJGUPSfBOQc4bfcC/zWaa3a/2+5Hh7AtPYIo1gOlVhjC3NQUuwse8wp/5e114CEJFepWPAt7Tl86
6o7YooeKRKEhUmvTxIoNAO9gVh4FSSgYrYUXU3G62bPk8suUB8zO1d3GSHjw3OlGSPOKDdLe6FaQ
XXJx0P4rIYKSy4bU+G0O29Z8kFS95xz91/oebe8tTELjtxl/ACkIaL9Tf7c6TRh5JpysF3zqoxv6
ntFaUxlJ2ZmJ2BYg1lQJoxPqjNmyfzg1/PLBQ+dAA1481IbgIT1BODkkf7v8HLgdA/0nYsUPyOM8
qeXV+ATnn/ltH6FZkXWf2+Eik+QUc9eIJOnAWdYDTXjjaubhXt/uOejV1rKT1VHuSET7pPxNoHNo
DgFXIoIW+IeBHWwh/KmLb/ScFGWEKdCZe/Uq1IWyU6+I3EPl/5Ko+ZPDUu4WMMTS1NVbp19fdq4m
JA4C7a2s13Mb/yPN3WVssEoUOoJeWsRfo74NG7TvH9++I4dS2SkIkUnKVuOidOlUib5WbL1pNelK
CsFLasH69i/kGPyiu6Gr+q9X7+a+NSJezKPzmwodext748Ly+k8ue4XjuN1ccSxTfkuVvl3fDHzo
8aCU2Rp0Y43lQ3m0rUjwhfbwkMf81xeCfxTTYtmrGCFRQAkZSOhQ+DkpSfS/injNzLQdGbjXuFKH
uR/vs6ciEBuKH+olOVHB4tnstvemXRuFS7+HWJsCffIVICxaQY1at8H8pqtSK2QMSUCCJ6Sdjoxv
XKmv5LjFe3TwPJ30jWa2tAe5QTvzikDVj7ChxYsjyue9M5Lppjz3mGkNPZgzwP35s7t7Hgfq8P/2
tEn4FrI7KGFHDNaKMyTWYXCENmMmcmfQO1y1MrUC7WA3WWo6GGKp9mcjo53qRBFVrqTkYRvEU1D5
i37ZmiHUXntnqxL4ObSyz4Os5fJfp+DTGJjIn/6i4blehT6acWwpXs0HGaDzRD30s+tTAD857k2u
i17aT1NOsCxC3auR+miHw4poDR+MW6nNN2GWyu6ubQQS0h0br7J+isIDgz8igcLejagE3SeTLFSC
YTzjtowdYNyXHs5uZUcBsgY3NpBZnyQ7PT67KHDZbDjKEfu+1ilPNj/RU04KmZG3/f8NBKTEHEel
fYPe9lGHDI4TfNfc60onAKYHIvJEIwa0+QzC6/AUskuGovfAYlzz2SepAfN3kO0swApgjYq9aDbC
S5xT8mTqtEB4QbCSPAeeCSsjuOkm4fY3l7IXuUJAptXVl6TW3/REtz9eT6dswzECuBNGG9Aua150
YnzsmcVAeRcN5y4HWTXQmZStbROkI0Zt95vtnN9Ya57VwtNxgFgwlL5Gfh8KuZu/hedJLB9aO8oX
G9Uw7lk/JkDTWYy4d9a0BfAs8asZUyWrgipEoYYLr1pCqTpw4sknpE9be4xYm0M91FWT/tlB08Ss
4OJSWfLA7IgNFdVWj/sJQBaLJxrLKPGEC6i8vRJlpxkiGMWCzj6zWx0H1FpzrxHMsJItE//fddQF
/8YaombIJeiTpX7n1VrMw39+WEnbj42EYGgKf1wDZs7jmDkTz4aONAo/G7Ju1G5k0tI7BT+assuB
JBqjJfF5QLLeZ1fm1IgjAbTrabCAHo2VsMmhSyJ3WhINY/HFWS8K+tvEJv+LGO9OGjpcFZHuR4cJ
GBwpFm2SWKmknnldTtbwd3krIv56LGjkwCo9CNWI0tPiCdJJVZRB8GxDk4C50RAyQxCsDkZYNBM0
BkNBBNsVdjcbe5ctCvxdFo6AdaQfghVXi6mJZcTFgEKArXsMsQJoQ1pj539T4EkGmE2A3Yn6qi8F
XdUvWBltFYZzSy2myMYJBlMyC4ajF+u5qcazPcAa+UlyXfM8Q6thDn/9PrRR54xyV+6Ll06DYFQy
/SHHtSDoAmB7g8OC6ZO9loh5lG4JtDiZZwpaYTE6SNMrfHNAv7Sm3t2HP6XuRKney/WnjHCXxTk4
fNrX1pdB2xjA2hAaWOiPKimlcTrd8li9uiT5YOdL8NaKWTHg08Fk3AX5Eryd9rP4H7rTQguPStrM
tdSDoMxTIb+mV4CiJDAQLsu1metuvnw6FlvZJUs0MnyAbx8aNLSVze381/5VoYuFcmjH1CAdzwqG
L8HqmTdFMD6N1pcDOWfLV2uu8dxYDTJrK3uLK5KMlCCThryXGeFw/3pAQ5HkqDxKia2hGtQ+VbO1
AodL2SJuoDrzKTpooN3o+nvpFprXpQLlznaniCCw++kj/g6gfv8ZfiiPLDCo3P8C/yJg9aztBffU
98C0/4M9VY252e29ly76IBUJIV31IynSlskH+xT65Z8VSUbdIXqVxwXlrFdq1sTfitkb9wBV4EVq
TSQVGnM+a/ubqhadey4Zgap1gQVYkpI2d0GPXrC7xlXcpMqiAdGiqsBeSN2timcRz69AXbmeXJu3
L2M5hKuEDd8iObv4aU4WhTDpyEutEZEveX3N8BoyiYAaveNsx59oG8ZUEtD3jhGb6g29S9vhpkea
65CY4F+VIod89qxWp5cypKM9Ocyivmxv+KcXPu7IY0qobg4NJeQdS+fp7ixxDtWM6WjhrrlLng35
/68y+dMk2ZjwGlatciH184BpNpiy8zRZFPwChdLfc/4onRNkk1KpWi8twtCu8DXsPS3UE6yJjkKT
VO4wjo5+JJ6cnpNrsxqOtVKrnO9rwc3zk4gXA9ERXF2isG9xF7VwmHE0+hFHqFDAOX9k1Iyk8a8m
XCVZVWxzTBkV9GdutDzebIxRqIDpIH2p5SJA+lbX4lj2mm/w+pQ4Ziof/4EDj4Fcu1a5JFBgdGWi
av9CWyCO2zkfJ9S3cjO3c+OC8DeFjmICyvt/cZV0Whz7cPytmc7OV6YFqH9v2C00YdHqrleGnJp8
1nEVTc2dMQpPBk5zxwsDzR2S7tkH/E08TNyf0A5gYOOcTJ87oaC02UhnhPBgbqZagr03p9x5o2AY
rgy1onTjUJlDuIOz80rnJZChgbdRbrGd5HZa45ALDz8AOQn/kR+hq0ipVFXYQ7ABnFyCyjgIq+96
i5v4kVairNAMX48nRLXrWHPeLDVN7FJe4Dp6zKAP2sduldDEjaFRm779l7EUObccwxEE88NJsVx9
l8ldtFWekSk5Iv4qI2Loc1EO1s7FhFogLnmCI5w+N7vnZO3KHw86jsHasqtuyrQZzzTvddqZaU/S
0os/5dMFWd2WwyJBPniIDuz614VNDlizHoLhTaag1KakLDE0l94y4nLSaI8mrgDfVPrBKiR1oLOW
cq66kYmIuOm/qse18IsGumcqh2zFH/Ibp4foDwc5cuzHe1R2C7wbp+Rv1Gzo5D2rYOefUpxRxnTG
n2J+CQhqXCsjWvDKh0GrprudDTJanjhJv4XyR6OtyVewS9YSEBwJgH2tiY4htM3P3hP39PHjKkDX
PDuzpGx5ZFRhzEUSZryde2MN/jCjgC3zWYa+5kdLlL+1qFhyWzzLloq+9sXSaiiqoxJiktpKbIUi
zLtwFlUgl0k6riUvgE+falE2fB4ENSM4sFWdv868Wu27849efX5p2sEy7g8tT8oQ9q1wvJqOv/1x
+TbOlU1hkkekqIoDQV2qazDtHVyaIUYtoDmPJbAXp0GECgPYTLxzSbjvByyyzaSmFNT6ucQXPvma
r5iM6tZbrwYerktrJ/VvUeAwlm3Pjzfw78jdRIY+r4c5guijrShgA5odWy9i2RkP6s208mfj6S0N
j9rwnmrUVjV8Ocw5LUedEnoRO5XUGkykAPOcroD9kHjHoYAEed4EZqxVuN56zYDjEpM2F9EHk75D
PtIh9T4eWRk6X74RAwntjyuSlb9zj6vuLEPaESzD6YnI5KKNOCry4iS1AfUTuiqQOrMFBybyau8l
lPDU5I+I3Ib6NQkblYP+TVlLv8W8weKwF5QoT4vtSGsCmSpQ+0/BfXb61hD2v4I0jjf5WeOP7ob4
7QIrNrbvEcBO0QNpmoLs5m4yY6DqlNHkBJHhnR6vT0uqA9+Y8bDzi7FsY0mDiZprUmLzXCTK42XD
SSP6J1H1cmKtRz4yh2arIeXFVoG4aMp2mQjTumfwoQTNGy1C4hGiQwnn1FktW/f+jR0j0MKsSP27
ByWJx2QVF69+q6RvSxP11prFf5OPEK5Z4Z5bL+CZDeUI+JInkF6w9rzCSV/Qjs4AwxZhgNo9P7wO
Co5c+N5uULoyJA748iQQxhZFgEF3dLUH5beFM8y6xevGpyVtGNZ6sDUl+mhmMPiF4m9PVQw/Bxun
9QaRMmlQ7TkKuf1yv11xsK+y0sKPHkL3/0pkLo2rX0qgNpIjxPdZ3GiskFp6KmLh4nW87REvYtdj
siw8acQ+Jt7Ke8YQ/j6Y/DtEa5Ea+YQxXD9zjjbJuKpi71cg2aRaPO8Bl0rkX0eRYakRbG150Nw9
+y/i1D1d+io4DrWhjuOm33FNOwuqXWCgu7swOaaCVLB32PxqxS+iiUj88aDBTAiFePhuM7MBFGZ6
0o0pH/b5dqGr/VnF6dipoB44L0dZcupiFeI7RWv8iD6DZ2Qf84m1WcZ2rClespnjlXC4rKNwPZ52
0PovvYcPXuvK3aMJoMsM4orlXTHxikGbWFNpz9GflbYGiWu4873zS+mB97s3MmTfXZoVqss8CCAi
biBfJ0HfqdLlPntuXdYDYam8YoYwqyvV7CwtQ7uyb/bgM1XNFZT5Vny/42JUh+qrlQudliLUo4vg
haCpFbYdLxw4dbQ+5ByCNrpN3bNfW3lnBS3vPPHhuEyja4feq1IYd+DARoN573BpQzUaaSTegsL+
p3wMGbHTE5u9AN2iKl7Hc8Ph/N+0SKkgipJLzTNHAQ9tyv9yBh2FChXrDp+e5kf5wIkKKw9FxPuG
ExeiX54owzLkZ/8InkyE234a8t6Yb4uE2UVcauQPXF7PlLu8GmkNiqs+R+wXAVaxG3DEEO8pj9Ld
SbWSJdcOtNnuWWHdkP1gA6z0iVXoHvG6jEdxLaYKlfqEkpc+vmV/AnssTARUjuG1S4aeO2M4jo5s
316JPvx2B1enTFETNMvJZwT8ysP+Ouafgs2eEI0TFoZ8UYLpH6A00Jx7KTsMhqIAu+9gBTRWIXjP
SLTZqryxhA6jcysTbRNTS7Mm32R4NI4UZMb1wUdL8sfEMC0Oe4wuu9xA3/jWSr5nW9LCRkZbXzPM
ABTH4E/sz7Et8TzkV6aSJvXu/hp8mtxqj8admvcYakSl3pVO52i8I8o9slINmmqYuPzkKjzIjWnH
XTgQbyywC8KtBhdZwu7IES6wZJgx/rzURfOByptxsoFdZSv+y6owyLoj9KAhCKkj7iQiw8Q/Ikbp
1/klyEyv2ypBphdhStsnLncqhIVd5jHecTZpnb2ZEwewspE0QdqjmudYvYLfp4ka98b9e5GAD1j9
RJE1noQHZSB70RLyJXMiWKX23kFzCRheg4ASlzogereS/QZ10MKWX+NNWJoNHj0qsJdG8QxJI6DV
A5HhvWmEhQNUGAu+FwwT4gCjKh3+1YSvW1QCmi4D+wAaKpUdBlHr52HizQVnhSFNBzUPn2lGjVMZ
8gZagrD8uYM0sFC002T6oYxS9w2/yA8cVXT+QXoTChI7UQYqLIWJ0EeMflOL2BErqw+a8xu94eTj
QUtiPxreBgwWq3w3KDazumJB0J0lZxy4SftgST3wzU30BMRjK/tqoDg2VkuOWz8Df3lj0DvC30r7
IVYOHVSmRozZAWiPMOzSPdz9sXAJfcGRaqVbOzT37nT+YDfDwbr9N+d9bzzfbwyBQhx0L80tj1uN
SGyGJu0lw7t8HuSQ/Q4oyjkyR09xj6te1RCxMZZI76qma//EPCUJltLj19k4jqPeq3+AiTziJli7
ebjYs1IDl69QZou+30m9hFjY8uC3832tkeXYUnJG2zI3G0kR2yGebBox+YMr5/q/pGj6LzptmPqT
JmXrQIU1rkWpP2/hZW3HeCPYWDNXoed3HlZZwEI9mRckh4FSeJHbcenPZp/Y4vSYkQHG/WIr804x
mpfIdlCqhbHahV4vKgY+OIq2PJc5qVkOozg9AFo1rTIrh60Pg2D4pz0LAwyaxieT9iy4hFq0bZFu
dCyDojKT5HQzseQQRwBKpfC2xLnP0xuhj1TAwAZfph/0YwKfR8pHcNTIhp85Fzp8Fox5r1cnWyFi
mKwjGf7K7ZBzLkUNPHgfA7k9IiGMNl+ksnU1/ZX0vB1x52pWUGrmCURV9vhlMz1qMSJFP6O1APKa
byC5Dt3Qqh5PoqtO9UBsosUTfPCuko4lUitvfmU1k6YqM4GRZhaPgkMwvM7vuZB5KxBkvu8xj7UP
BRF4Ycw5yvL3yomczZrlljo8tMz2eUOd70bogBa9XcXzoR9bsE/aUm6C/fEupMtvw62UCdGldQSv
VNc3xKD5feDXuG3P0hcVdaPKbgbHNe7RgvnpRp9TKZdC8w22XC65kdM6Kk6xIXBBfBzjcxd3dpCw
zHh5KQftiC4VB1kDp01jEF24xMEEqw46XIgomnCiidblZK7HjYr1AYCHTHxAb/NG+X0D5yqO9/Dd
DXetfmQQyCVNppb2evJ0u5SGwP7POHIzxdM2CEloeSfo/WOazwlMwOlTzljzoMfW8mgmLEaZZRCy
CHl6+ZpywR5o1h4e9WQPMhoIvDkvWvVkw65VEZSOXvXFAACP/nrcGgQXY80TQIN4+uMqyfNyJC3x
os0J/uXQ89tJK1uPcrWXnXzJgY4pcPY+O9xdXE9dHURyLJLihS+AfB37obyYLPTr1hm8cLb7cUXS
PbZUUBJRkok+WkRbz4SBi4SxtWe9IZ2UuUVhRRF3my/iaDjkbfCVGAg6VWhugq0wyZgFRYInNWh1
HlwRwldEZydWT0nUo8ZfjlGzhNXqkgOsWM9AYPXLUYmUeEs7dps45a4IQmktKHU5gtLjHZDUHD5W
9DDCpdtmUz2Sk4us8bDHFvgvXaGIyS+5AkyjkQE7lCQ5tRpX6UfDFyA0z8TNG5Mh6Qsz+v31fgp9
xMtIEVy76eN3XrmSQqnw75OxAAU8+xHmMeQAqT3QIJPXjKMru965Lz4IOBAgWEynel0RS4Jw64XF
l4imMScreTtJhH4bB7OX6z7RlaeTcczVzPhZCJfmaOqa5D5RlFvkNdW+xhT442gWdmMRRkeBhBbJ
U2yZGT9NF5IO8brgegT9ItZgIZcs1wX51QVwzURBeD/vU2t4RzkzYbg/QsMUtj17BLbrsxCbEu0Q
ZmIi95Apt2pXfezMYaXVqVwL9fCt3zoc0jNCK36d/QO18Uo1VTSYh6MOyo8K5Dbj1o5qugjGKY8j
01Ih5TZ3YHkWEauc4RT6W4kI2WsaHj+97+H7DTTAQAQmxriJ5QNX/dNTrHKgF9+QZ+/ObHAUpYAR
Q0yfvKz0HlWYycLxair7UsNVCrsvqNZXPdUMgNbXfBlZu8mOiVVnzYtQYoLH2vSaiIdGek0t8EV5
hBAP3hNKMO/e49O3hlHPpM1OkaV3hGxhVtbmynRflSuiwOZWI82aiMn3sutSilrHoQpCHScn+6jP
hlPNx3KOdP+5x9okHd3O4Uh0b4jarj4LSI4W5W61KEpYkB8SDydZB4BhkmVNgWPZ8OpFSO9++JSU
7K/n0woAWNhk99I+wIUW05P6NV4n4/Spl4niGZBW07ZZV0xHyfCWlk5XjT4wPE/sDYLliUTWffS9
J/vRm5tvoDiQ0kBKsm35G3jwIpmIaL6sUZM2DlDqmboqhVNJApgFIEZRJagSxyWxXyOdncDxvPN4
VYgvLGQSiY2bhLW/+b5tD8WiLGe1v0pM/yjGDyujlt8FsT5YsCbJqZrQnRwQAXra5MWSgJsIkImX
hq7T2gi2zioxtr4cOUzg7mZGX/WFG9AnZqRk4IKbln3fZC1atg6szLNPfaTtl46ztDakQ3EOMsBu
7gjXxA6+PqORkmcGf4ghQknljExl72Xm9ZHqHg/v9b8F4ueaN1HwLUPpKlyH0WPELmzKUCFycJxN
pxv7SowbSwQw2sSDb+ci4Wpxc1DhIBOOIlpsEd4bwt95VMRvFkTBjca8W38CPN3LLpVEszDPXODE
mXSdUreaYYQzPECCo7g+uEQzsD4lCyUk7DPoc0axzY5eYXXw/jdZKXKvx6yJfNQC0dXPeBASMceF
dZXdUyvAg46fKlgEjT1GLI/lJTwV0Ke1BOMb6idV1dI2JFoQpo6OJQ6zmtrcfHqTkCL4C10RNHED
voFfHBDxHiyRHT7HlQBEd9NHyR9R76yp38GmEcOf0Up28pm+nRtDj2cXjyGD4W7qiUCaipsgnxMI
k60eHIQ4yfDfqtBzRZSAV2sajLnsWypFNyLHkTLH2OtqHlatGOPLx5EWVV5ty8rdwjwT6QcWv3fx
lGZQ1Gd7zj7XKkh+2FA4dPNTklsW2O5cwqSQfYQ12lfSEPNKX6MAovtMV63JwGx2Rm2/MGimIM5l
aBCMRtisKMPE8WMzYm+CPUUbAetmmRogVVd2SQ8rF9Vp1k1xlvIvlPIrojRsOdHME8wp3pbC7MZy
5pNgPctjrRIem3ClOOs2qxjvKh3aljCb7y6Z7QcpkWQxdYHLCL5eoUpyftsVVZsgiBx6I5Y2i1Ux
Cw7s52EoDcjNbOQ0zRK5BbxT7TCNO9lV6DSicZ2sB/zjZvUFT0gNMNQW9Y2a4Zgir1FwG+2wYBLL
WtXkgzIQZmEmYwywsbmH1U7wSfPwV7LeOn5u8TYji8zKt9clSBTarlU/rJuXTsqFVzetyfzWmDvh
lnb1mb28GsTJ62zQJePM+NZat2N7tGkyvbc1Mj3pCyA0TemHfCOWyjs+vnp2vh/mfhe8p85UDP3M
8mX+TJNgmLROQxFFGLEAs0M9XUm02utrWl3SbW7fDQU68iSuDM3MuUEYxPzPnlyAB6zVpa9yviXa
tDJ94nvPOT5CXwY9rODTm9wcvyvE6FImnS1TUx9codFfOiwppOVTt4GOmnu0BvigkkFtX9PkolhR
gqBfBd6115FG6r16iUH8IBqE0VeAUnZ6+2EXkaiq6xSQVhp+womt6fl855XOWiJhlvgAgllPVxuA
ueXZp748iKhQMxvTRdBJ5uz81kkKVTHL5KesE5yIDne5dx93X04SOMsr1CR7AYALvbMtlB9POXIR
lyAHQXx8qoUUvRKWEyySlceXIbLlrQYefWIV47V77RDUFK1QliUR1g31dfCvbzuvUiJonIdSZ3Yb
a70iGLq98UXp8RI0Z7JUXXcaStC6mVQ8mH3bZ2zoRdNCkCt/L3DgZAgcW4PRRYabpm6M4aPrnS83
fl0WN5FUmEcHBH2JAX/OFbxgmIe3aTR5FezKGiKyhUKRNK4aYySbe0eSSZup/4EV/oO9L2mkrghZ
QVnbNJcFoR5YzfGoCz//0M8ZAAo01Eju41ZYiVjp9BSmaKDWuzbfoO6lxCtaaLaZr+ACstiKZzw8
p34bd9oLFpD7NbHW+n3eGZQ9H3MEynSzNojVV1hLzi631Bs4GLWAUwJneRn7uNV88gdTheS84ynh
3JQsf+x5cHR/Du+aaJcaHxmShzqEO7EPRxrj63FCMOpTGWODAxfNmucTd4EYMO23Hc5wvQ4RgGKd
pEc9M6RD44dF54Blo3Pb9rXvXqSUlrGFPAMRakFN9VsvnOa4wrKYC075DrnVWDyKoRFeK50BkZmL
UINbzYI7b5Ha4ZE79goLfwMiKoJtbMKAQ1X3MdGfDMe9qS8kngwiOpYlh5eQvK/OuE2nZbPa0kwc
Q54QogfQvPzWFxLmoFWScAvEyUbGFV1m0o4sHIrtHM99emSkxGLTuwVSkivpfCzPPJUZavZ/vTfP
789GHKLlclHxMnmRABJvbpNN/hQZJ9VYwK6ArppgEKo7/bgNd5wVlBns9FcvcnCm8PgU0e/d+03/
YWkwhDlj4IUL6lexO4IbCdQslAa3b70R0l6pLyTtSGvxqSCiFw+QzwaJO+f/jl1lTk8agOL/ryQk
yAIQVO8lbCfJbr+afPjeoO3KtEh8/wea8KINuFm9B7+gcGGCR1HpS8yZC7FFzbtdr7FbzaJEe6qm
KOVqdtPbniH7asqf3i4FXWFXkV30wzSb4r7Urt1zKICZ6FAiWvRWTXeQRPK/35DM8pICVkMKoM6P
4xvH2YoCh0+BXftHuhIxsWR1kQvG3Jizm3lEklznm0XYQYUVGPJfqDpQU4JEBoc0LApCerS1rh+1
hDgnWBalTEwMdWHozaLg1t2EBMr08kC57qCKtouS4rO2eEhvZvmTwvenUsnn6INFiCcK/5noAXMI
XmEmK2vdL7aswXSxC3inDgAlopzXtHBerVnJzNlYaa/ct12dU/0Mnerf2gjlu2D9m0LX2kyIOdqZ
BsCge+aRrKM5fEy3Ix6DS4NVgOcqDUr48q7Tx2iKyXVv2mgBgzkkcFhNnHfAySahT9jSJaVswfGC
lzmAW32xyc1nrhR43MZtO18XJUSCUlib8CxA2vBm/GEwsInMbzlGjRP/3oQnmxmY7ib/3AsySXFU
+VMRnu7wIMWh2ksxK0A88qIQESxioai1jXYOD2kGIQqjMVTc1SeymwL9HMzd5PyAD7OH0tD+5Ncj
hH5uTkJuJmmR208XCZYnJySvi496lF3E3jTgESScJTTsukPxvNx3/lKxL+Rtfmo7Fss4T0izE3Va
pT3HIHdV/GkFyVLZCPF3kie88ss5/EBRga0IWUBh69K3Tm4nTbM/2kRcqr7AWwFun47cxq/jXRtx
5dlzIf/G4eyN3AntjOM7T0zsftUQXu6jU+aEoHjBiROQ7wndJ8/6i9Gz6LkppTSUJsYGi1Lp+Zvn
6CjB/2NB93XZJEb/H1tcyVESy2QT5ryswsk7UDedW72DIbqpwwiprYscxfvOXwfALsj4KRMR2qvB
XseyJNZP2mwRk/jJBaPTQuMz0YZzesiKTC34uRAxqgUVx/8lssaIAyk2RVgwcmvRcrIV2WMAhG2p
rkEOqlYePAZdgsezgtMHBPqa0lZIzyCFafBgRBAm9lKru90HRTsOLVVr3+Zl9kzlh/T+UHP6fQ5b
LzG+Gk+5Ua+LuWGgWWcehK0hUGh97mTBID73uJIgj95PoTANHh9/Qp+9YeJ2WgvNYkQVGiCQ6esg
cR0NmIykv9tVn0B4bIfoj7bvIaIIPkb9n0JdZxJsTHjhEI6koR5nXKF9Wpn/8fpL3JtNJfqmpb/1
nNdb0irUJKqghQBKfgA6rAFtJxjKpAKlfEN+v0GB9Bg7EKQ02uaW7p17e9sndnIlKON6YFfpS6lf
EEAeqAjkBQqa8+i32RIJV4SsHQ2yvofqCezADrzXbY9khhtOla77dVWBKNTI3T6H2kW/u0tI0yPs
dy/uU3lRNrJNxIJG8IMKqC/29qiNewb2vg95Qj8aLAFO4TCwiEEAXhRRm9dLRFWdJUsFajgK3cVd
Vf+AJX8EPzhqFKQRs2C50BVXLuyQ+CHXhjjem3iuDmWrLoR9TJkExPPkCMXSZPyRYVdIgf6oOJn5
rhlfxR0BHgPWiUMNifhBAXTPyEwRRdzItON2BAcjcuE4D52Yr3DFWArWQKAhQxayNZG6uorAVzrw
OwNPelFSSY/9plyuV4TS1g79jR2Ga666+ZYeQInO05E4YR/BRuatzeKofdZNdWg2VpNqsPYravCz
uKhQ0rjpa1+BHmSmzsiCSvS31hl6LWzJfkBePdaSC5RZ+nnnGRsmW92644rDAswRaFg3Em8DTB7M
qsvLKvhu5HT56wYmdzcUJypDTH7QLpnxzSSCofJgEhVVwM55pilSBZCBSI8orO02YsfAf4OZF6f3
Ir5fM12ryBTvKOOcC2acSTkzf/JegmWlwDGagB69zrsexJ6kAxPPvJMufLyp6paPqXxdr76ulU1E
sEQsXzGeEFj/nEygtKKsBn7tHTzKgb8+gVJJftZnaX3YRTlKdamaVPftZWkHFbywer/bACfDUfug
96zfx3bU5eRy112LtoLmVbbNik+vHVxDqcKFu/dYzDka0qeLiQWnWREY+wLdqLbQXEVE3HQCBsF9
cyng/40VFiurbDmO+qlP4prAFaVEu9Z5sF0FRhe/3kd2s3iM1bXU7+PltAx7wbo6omfs6Tm+yui7
jfB8YkRtkohTLm3nxQUSQ0epngQKALSkg0sTy+BSLcyCmqyKZWFWei3BgXJAkDHejy0FNi+nz8hG
qb7zOVC7+XUloCcW/7vbMnZ1K+BCrLLMLlqWFm08iV4//cIfs1hqEhkofr9vbrq9TNMV48c40/AS
rVVOLbVQ3bSaliLs5iINfHGNhKrvF3wTWZvl9Vf1xCbiFPmzV+fEAJQi2NZ1utm7vuQChvsO7H/m
9zmiRzL3kh2mkAJOthMNS8TJhpzegxOxV9OnLW6Q2B2uoYU2NDv9ywiqFH+YbYvNFd7NFTHgnJPy
kLYIsaIoZ4pm3uB4Z3pAQ3XIoMi16jbHLUVKppr4e1R5XIuT43o9UOh0aDegVGVCSfHtu0Rl6KQe
tSLvewN96MqLD8bWHpYHp/Epyg4anEBd0VoVXrLQP41iSlZYtAMcV1LPfJF1msDtSDKLNSyf9bso
uo2mcbD1ASFOjES2XlDnV0gezKPgTOSW9k0K46pDZ+ugyD0qX4sgdf0Ea8tALL++A0OAYz6FdgA9
yfV/5t1Cr70gcJPsHcOoUvPvkbA335YuudITh56K4l/oPzXl8BYSIAH5BTrITGAOuwYE5yk9mFEQ
0xX/XlATb6EmPNJ3bO4myIdcmuuMlcifAiV3+a7W3gP1KpcAozEQ90WI3dZfHSSESdKFf72j3FlS
UpSpT4RICMeDfUOu0/IrwX9jZS40v0GTDGAsc0uBojeJEsgVyoIAauq58TfHxn3XrnNmMspwsvk8
AqHcnbsEwhLilj5ROvPsjrLpmaoA3Roqzi1xEKZgknTqxt5YzFEj5pakfbloWVAtvdZZYyRaC3Hf
bdN4GAJkmeTk5LoVDEUyrQkqZyCyAgIObNgNi2tg/u7q15T6YB85gyBNt03uxu52dI63O6CAs1wo
IwA0LDu8BV836JSCL3/imNG9D1YkZ6+1JLfFYS0dalIip5LNuhe+52PX8UruszpwsgL6k4v4J5YK
E4xZOC5YvsDGBwEEsrofJK+ZufVICLJrDH2qX4dYeoq6u68SpFfIuZ7/9joI5QOuxCuzXj/fuQO1
BXTFEZ0WSnf3evq/Xi9LW2ykZ7lter6G7oRJbpEVl3OC1KZ7bPih11qNJZR8UGowXoyNzks3HApH
QdP1/NoudgZqGqOtKx3R0ld0NOnmYfZsT+/QTnhf04pGen9gbosvvIyh8tvRHaGNnjJNl71R1CxA
h/5i4AZ0Elb8F2+xtRdqur9a7hx4v/x69m9yhpJs66Q+SIidTnUJk3W5DrLt9tEW1OSf8ijxj3B1
k8ZQVJylhPsqyZjHqry/cW2vcXk75SpPqs8hemZJJETPT3PagGuIr9uAwJM3X+ghzbeABELKZiLc
uoIk5FVy9c1hSot2jDog63g+tTR78SYrvgX4ZdOyXBIIqC0GzFrNtDgz5O20x5jk4vvQqeJHRR9a
CHg8J7fDeaMurB/90IfoYUjet4HrksPYluNuX6nIQsnNgxD4AF47iYYbeN39EMcklzGTJxQSp7gB
hiuorWwdFTQ0FIJQQHG2bh40yseRru+E6X9SDtw0a7M1Er14p48TH6Wc6/1u82gmaz4tcnGPoYNN
niRVIBn6AdAarfgSZV9yVZFrcNvALqJD6NIGeDi8eCKhMT74dwdtw5c0uK4hqLeQ89M6v+js+KOQ
U2nUnyTRKV6By25KIaffJdQLEFyCfZmEBa5yV2bAqXrfhJk0cgCCgsgGvswDV/C90hG3CUTwqNmS
1sfR2As13uEVjWk9PSqkN3id3/zBcJxgfxCkdpKrEc1G4ZIHdpv1QguEKUQRY8l0NNSeLy8ym1ME
LgdGmE1UQz3M2U3D8YWKrFIjlGPgduRj2BJvtqnAx+jf0HzEb3+JCI9tcr/qBH+KHCGKEvK/lEue
MD2VrWtzpKeqNGdzX84D9aOBPVPZ7V/jgvTUcWMnNm7MEQc2v2sKPho1Y5pCWI1RXOIHL/QT6Z+i
Bv2YTYGe/q2wf3Wl++NbUp/e5SOsgtkRO3QL6vyAjrKCEEjUHYiqFWZ6tU1QS1Uc2QGAIFGzAcz5
XIwKkPo7I1e/uB/JimoIiKFecazCqzROdf6ln961Q7cclbmUxsQnzysoBmy2XlK0mlK+IXU37adC
jsNfl+ybUny4c25WDWqqwXXem658wL0EmeaC5N1FcVFnTfw4prrYKEUqtDk86mkRBP9sxM4v/Vd2
TgBUOavRUHlvjHrKIdz/75cCradZDUzbpery/n77B2UMC5GR+zHtfaq7LEDXfk/RexRBvCf7ftF/
pZ5ETMjGu1eWeqSXSgWdxXWd1zBKZsVOMPUkF4HbXrNVEO35BVdtuSadkKspkKJQbZJ1uP91U+4v
kPwzNh55tIvPb7HmLaCFEyWu1EvGsHCLJXiIiWQvR59xeDQmefigbxiJjScafTfijL0hOK4Cnk9t
I/0Rw37Gmp709pPvA80VDbzGtGumnnUnKbP+PPxn5fIOMS8n7bpz+rOHUy7glYoHCFpzum7ElZZF
bb4Y4ibci+WlT7jIyPcHP8ZrLBZYF8BwBiiCLj4/jqiIMhO6NJ4DR0c1Nzw6GwE0YjSVW5+2cRn2
4cfAKDn3kbpLN11wWsyyDLvlEjjCnILlX+V/dThkfnn3AG6zFJWp0xof7qwAj0Z6Mtin5wV5v62Y
dEbzwmmod8KImyDrqBntc+fqztRt76ZZ337AdhCBNZg42XWlG/TglMogrWK5m533MBcuKV4XnpBr
/X0h5lJxLaQuvwy+Rb8hCjrajlvK3adVQSmf/vZy+kmtNeLxbPkVOLkSPvX0aHhYpvVQiPENGAGs
Z3qKctK2XZowZ5IBXawRePjBEZ7gzBPanh75VQnzFT1xO62Mh6b2XT//1YuyhGos35yArjGdRMz/
rDFRaCVF1pyYLoOITe7pGgx8/tp0XP/8lJKKM3z75/2o9tVAcauwI47wLz7i6hgg3MX4aVnje1SN
ugGjXDUPI1cjGLIw7SgCaW7S21p+PSm+ENylXXRMYpTMuynTZ5t9T7Yn6qzgVhchMW+bcL5qsGaW
PcoOroXlpaUNUvgcarHJjkzBxO/oWlM89eDgRgb5hoq373OZWVaJ4GW5X8vuJ1aorAP+jon3l2cC
31/354X+Zs/q7dH0vbxKhrauTFZbtGS5E+fHCC0/PlRDhFt4p5LEf2Nd8vGQxRTnRBrV5O4+SPQc
4DDxdvDCWhEknlwv68umV7DYH2J2VkooxLHiVVW9+TF8Cuxw3EMu6S4BE8wBMaF/nbwICGYQWp15
SDSwrp6SQDgCfLMeQhpXnpCS5WRzGAkxJ8hZS64bQPMIa0p55AFt8ue793uI0J7iIfmeVQAE/eHY
vNWkX2x/qKDzU5tlGMH4Rp3WfRx1OXc1WyH64E66Y6lc43C4KO7/rG4KUoKaQ33p0NuP+B8hDjVz
bYJIdAVhqyid22nxVH7AXjuZAmC+L4Jm7s1w2bacT8fIBlHkiAOYNskFefIpE5NXRJ959xPUcCrV
mEMfwpLT5vPoTAr2mFr1bWJJKBKGRBrAIJgXpljFfiOY98AsjbxxkK0Fpm3KNnoyAQ1zopaZfiiq
2zZUvy8FzjRpdD2b6fRP+cslPPGnK5X6tBwr1U8Ca0unyCmkIUl6nNnK/3uQrUKOYjWX9KeaSqfQ
6puZ08z60dOBnTzzNSRk60dnDcQe+ouC63R323nZUSxG+IU75jk1rx9+IyiiGWvvU4bF9WgwWHbx
pTf6aVeniA8hPjYJJt4gF9f7bbXrjfWMKhO/R6sD+LD1br1wOYaeHrGauLuHPxPA2dsFgB+IKzeu
YzQsBgfz9oLARQnEelT+n3Evn/azo84G80m+hvaDjNHRam3P5MKvxD83hdA95gyS6G81QMmcyvlG
XW8sPgUKcFGpBhK+G3BzsiUtmEAuyj4cNpYQwvrbprNESlgDQiNqLG1CVYdbz5RvwLU69lGF4hP8
h+WXnVgc2/TlntDEbsKI7D1IOVmBS55knYMpIDE5wnF9y5NmNoJ7Yq9FvWse4SO3nhjfsqU7YuPU
nq7DLEBFhFWCb3AF1A0XQUKpQeLc7bwaTziY59wcwYQdzDwTTCsxM1d8y0sWSjVYtr9E7WQchHib
k1cKiRd/vDD3iPKm/AyMYLyjBSmOVNBMNvLCmiB1VfavsyqmXEG0O0knA6p6MfTbEPXZD/m3FweD
6tpqz1i4fY8Ir2CEJPGdf1OvOuwTk0VKCcrd2qq/jfFfOpgS5yW0GC5rTtjVkkCkyXC2+xt4H1ug
GuQGXrT02YVgTmE0Dm/4u4g0Ny23I22QOphlgr1/O4Dhb4bWjvJvwzuHBLedFJwFEW1ASn9g3mGO
eW1KQtxIYIcaLh45t7Ua8lVUODG9shkVEDZubFF402LeMPOmqW3V0Xq3P0XUHHy8DVyYOxcMGAiO
3cg8cBp9iZnEAzV3n27qCu7vwcTg0v52oXFo/XB9jOga4ut0X17slddhwaBCSBRtkcC0ZL/JWVfm
qHvgs0vezAOm3en7Y525rDaOSn28/hUsrpTeJbbgBYiQaZPTuj6xHGyqAGhG9wwZyr/tiYFgVZsl
Cd7hpZvk7QbZ627RkL2b/ffpBFPeo69Bg6kicQgLDqiBzJAWqNMZ5Xr+pH3lX3L+mLFgMnMrDKGS
6AtaeChZE0l8bx/dVv6OQyvfPBBvRwelvimYxWqUnR8Sb6tygJ5T6+KUhQBnSvi/eqf/2gBFWUWF
/dae2TvZcm/DjnDpENbsy7NFJDvxeXv9FshcZvSUtfGJQse/CFM/e4xG89uqVarCn2jWrC0ckodn
usz7X6ecfZxxdZvxcGpEvB590NwkKl5814wzXAxKFeohC7hfFIl4MAQ7xMYyyGULV6/S9GBY1ev9
Mz6NpildttgyHhs5egFu3pzORy+pkz58zwBvcOAaTUg/ZQfpxuE/GHl9kEIdG19SU6Ru496Mbp7+
DINQ0vzHg+80s4cJFtbwQIPgyNnNL63TJOpZSAlj2Gy4yxTL5iyEUlG8Y1/SMyytfnBfZE+l2GyE
5vwxt4Es2B/gLydJJPTMfhfDqL0o7rk8EM3Zyv5Q+usod9qJmXlQFOlaURCq+ChLB9blnvFDQH49
N5Xa/UFdMzTBe9CTLyz1Y1G9V8yOkSBWxyZZJEhz/IvhvUxOgmwlq2wFwu6u+rKE82/RpOk2nx6Y
qDkVhj7Kmcl1+P+dZjMk8dm8pUUwXqk14taNIIsy7a7+H8YUUoCyM956+r0U04K2MoqpSQi1q2eP
09TtO4Z5z5dPH91YCN/Ei91RhYmsBd38EHT2bG/KnA7YeBrFgH/eTgKwg5PJmygdo6nSslc63LBN
Q5qrDgFKGc9Y30sM1Vk3Jrh9baMQ4WazqAxanSt8pHnXGDYmi86k+voiy7l0Oje4x0lIL4+4E2yG
mNIEOb6BXrXp+eE8ZJYUP9s6j1RixpSzXHfZzqltmlFqWkUNZbETeN12PkysAdp81olDyrT6P+ee
9tHhzWAdsqRs6QnwMr/CoMI689Rh3Vj7RrhN/XCenFXTf/6SL5Dc5GhAwI+jcuf0LmTmrsBbEwkv
qT3S6XMF6hcNXXbPDlCURcnV3E5r6YRLQfcBF4176DfDcmwq8YDIn3GTNw60r41HunBx8qfMhXnx
BKgjMF29HVbkyxwsD1zTtaI44+knV0GPuce+ThgTM30qmcVofInCwUOu5zaPegH4FMPbjvl8K3xj
9e7A5vZaUiVJ4gDvbCzOMM4ajAadNapzWCXcHYKYMrCEtTFgvULIDdFzmrXexXvT15rScYO0hBke
pMcqmzUBpB6bkg6J4wTBZtjscj3bFnws/QzDEaGdwTRzUSMwwJo73elZoHMNu92c9W69xc6ZnOdM
DLNX4cm5e0YYDHiGVcybhXW9o4lzTG5YlI6XVcVLne8/8TIuU11cRBOQrGr92RsyYCl1fsW3a5dq
+AfifIpSPi6MNS/j5gcPpRLAs1IXYFbgPOCLJi3qIq5S9qyMp/9GrPmTyjwlQjeC0uYrKlwJ6W6l
v2dD75rXWyyG/Du1Qzb/wS2y/2+amNYqQ9Vwwc0Ofw2pilhw7bR+V9WH5tJTkKJfUvR1Uy/upxuR
/fbsPwc2qob13oaX4npgRRLtPnBmvkUiY1Kr3ng+CasG5aaoRHeCF6Bo2cIcausJvgeSG1xyTywL
YJ2hQCO3+X92QCaDLiyP3IEqlojn+G+f56sAA85vu7vp2qBF31V2F46zyAvIkWjO4flDijRg0fsy
frwNBUwzGrNgNy1LT9fkPrhnb5WhygygQb5TKoAPcY2fftVnIPDMazg50S9AKEAhuU/vMfSyRrIc
HzCRIRrR5mGP4Np/j/BSo4aW2aLBoU0Vfj5xWLNv53AElZP8kdllBqjKTkDeBD978xRFyOSIB9VH
9Tgck/YtDBJOjqUPmIfISfpaggxZG12KWpwHceE5MxQXcp3dvKqlUhlvpKQelYAV2kws4YC0JCIa
4DigXyhwN10UbihXvHfq9Pg1JHlDzn2ftN9k7EFnBwYNYb05QUD6e9MeXjx9XAXCAVfmC1GLn+4+
WFGKHHIPB7VsnwsKFqxLk4nBazn4bZjRjt2EprNJLfvDQf8x//ZAVnFfWSFeKVM2oeQ4Kayuli0Y
zMuEIagau3AF1Mb2y0H4prWfzdJOKxxsWCp4m8J3ZNDnS5/JBhLU4khydqblHuXbiCdXo3vFGi0p
UECbrPGvx0lHCugG9A4PPApYyo1fXGRwHmci8v7SJullxKyB5sJxuYpPSY5sSbGz+n2u4t6tFNrg
aDipKdl5GCVdNfZXqNXXN7QDdQbBGDDzqBj2vBTAPSdisoe4Glqz3eM+VgrRfkGue+fNWdizoBcU
Kutv0q5eInH62ioMsjjJkxdyZq+mwxd9+MgwXn5msq2rMZmUUdsP8q0N3OFZdqUqqu+J67mBxzZm
7uLXXs1q+4JPgz2d3NBbENa+Cfqna+nscIw2KIJON+CBsrLQL/FbVcykT0LxR/7m5fFWxOusy457
xg22NlIpkVh2aujGaLqZTSjB1u2iVzlEGtJb92uNe3eT2Uzx3jHWTU/jIRwEZ7sT6xLlwRXYEI3G
xrRnizrzo6fJ0GbnEolnjVq6WNRL+3zqFYYqu0KXHY8BHOHo2mT56hgD95sVhiv+c/GuzpkfXGbs
SQKZs8krxsMA6iY2ZOtTFCh78MxA4JrnQs0JBra6k1MLaL1ZcyT+0bgyypcJKCvEJezegnbXiiJO
X1MJ1YxRzsvySLfi8dBSJNE0dDc96vx5EOFbBU4E86y1UigjrENNc2oVhj0v5m6W6v13m1FllDTT
j8hiNsxxIFl2cIpjzC8+yEicGy0CnKiImj+LX2/GU05lPcQwZQi001gH7BFPsKgzub+Smh1pLkPE
bBxnPLCbUji0YlluoQ86s6zGfZf2wWWRCkYPTnsC9eEP3WQu2be8Tq1AF5g3cWrIP7eqC476/CcG
ncsfTuVCkr++mzj+xFNy+8SpddG6eUnRDtsfk5LOUmz/Ch9WNKAZCQAu5YpNelJG9Pg0GAkDkZ3n
YqQKRjN5hBrUMDa5/fhu5DPwRr/oEQE848G++Yco9wfaNUWSCBZq1xyP7aLJRvjPylPggHjxhvJI
uDGf1BiC+MFHYwEy2cF6ytt8bWnfBzetKK6N9PCUSCiQvVyFH1WCf9W5e0jnSvoi3+8L22rXiSt9
IVHHSn5dKLCNeOo5jCFJH57CPSQ6NKjYbwhQiXsswMBrdgDVStnVG7Gy43Ytxv92biYim2xvG03D
Ls4MtHH6lydKAXBz+VI9fzlQri8hJr7Bze9QjPW9OiRic0d/xf2hj0Zb/uBE/qVh9Hw6V0Pd6jMV
DcIIPXFNId9OIabvc9eoZpnezFso8O07yjB/ePPUnLXwaWAzEmXVhVcRLlibulEtl6IBxqEA01GL
qx+ZP739rXNdc2IBWMKLbVclQ4acQylz+lsdxfs5D3dLXdWc8v0rg8TOcD/CwU3hsBmsBjt9T8v3
fN0zSVG/c6eDeev1rEiUtKaTcaRwcup+oo9Os6ntr7oZ5Sit3Q/OnhZjwvjxCmam+KfX261S79cX
ju2dU9kr0uOfSRWlEwjVBS0n9Eq3MBJRcs84Stcuo0YgK0t+XBODppAJT8ra640HCNwmpDmOauTr
l3MVxJOgNy44fXIAVtNQZmgJIHCeVtNSMByX27quHDF2RAf8SieTeAP0DGoWpNlo1fovFSES0+EH
ey48SSGg+6yOgRvYQ8pvXVJxUnTkM+FWTAO8g9ouCR/GASCLt7leJ3v0k0yX2K+s2222g3e5EZev
ir4qaNQj7vFJEqpWffMXXitOQHmEuzjYb/fbecgKWQ9uAxXBPaz2kDPleTJcJyOQB1SqlZtI6fJd
8r8m9oM5mJnDn2n8tVt4LVw+9VWG2xSwydstgboZCYRGfCAzTN/jrcyiJhMYA/wY8cKz45AszDYn
2licpsNeMUat+xRsNbzZpsS+JNX5U3yOAI4O1GaiQAigViUsGbmZd68q96RD7/W3y/DCn6Ar0E4l
CFgykboTFKzApDOK+l3e2hzLSxlAeDo5oudQMwqUDHJ83TJlCHGuy3/jK+AiIX+r9c1am2kRbwlN
t5u4GhNAI//sVNFqW/pJnPgtJsPPvmvTrr7cmPcklT5ODwfaihmdp6p+rVmCpTnQkOaH1xMq39BS
3ypl5C0Tm0lZgWLee7cbxvid+VMgT2jh7UG3ElpP5J2gLRAj1+baKtzRioXGqO88BMfK3J2Dq2fK
U/0WMCwAxn14Rnhr1qI7WuKQsVmOySYsMbtOCRQtVTSOSlGvNvRoNMpXMzKMt278r4PyOBXZLkBD
7hjH/MBdOXvtq6Fkjz4qykwu4hJ6L7LgTGoWz0RWrGsBspZ10cj6AIwclZHKFmfrjrugZRjwP697
Ec56OlokhTUeolTA/xbejq3CzTe4H4FjeEztkM18gbptBGpPviD8h9GEGcsPX9lTORFGOGlVqVRE
P6Yn0jSeLung8DDgZpXBMwpZvi6e2iDWpn075GkMtyuk2+mRYbATMEF8Z9GuNaiAIyd5cHG0D+Hb
CSOOz3dC272pP+TQFM5pOhZHVj79ZUUMR3UbtRvLey2/gnddaSdmjxofuU5zLFvn5sbgibYf7q7c
rw8kONEEN4+NrOoTSH8Or542f/KmW3cK26Mhjozq4RUNHHgkp0HKBGQG0kFaA9Xvr5kVDbVJ2SfV
6oIQFobdSulEKzOQliU64Fb1rB0VqQqfRWB21/aEFsKOojtWDad0mbRec6zE3SzW1vS4edTWf6Wy
1WJo/cXDjjsvgEQyTyhJPqiar1tT+VuHBGHjPha4LEsuxEUz5n2+/Iq1zR4SrIpPWuYFHF/Tz/Ia
v/fXiRJ/FnbGAYwiO31VUATm4/PUPVcJao486WL7iFtiZhbbd58NcrPtHhQ0e1dCL69nnYwceqEb
t0Dck61DZQlqqjh2pxW2Y1yAgZbUEHTaskXFNX3YU/ILnXv65wF9arbZ5AC8IUmUzNTOys4j9q9H
ytIEINS+m3FO2J0ObT4xZAtUmA4Efwobn9MZPZb5ycQT8pVoKKidSM/lBurx6CojuzAA1tU4tq58
Xzy/YzonI1MCWB5odT4TZQcamI8Tv00M5SbEdxTZYMyoDD1l6QYivHDLIkdV/sUeXRbwy74mpL1f
enHGO3f4MlykIevl+E7/tiqjvbXghieBDZTftGWA4l+Mf9viYYuuINNTFfBj2qu3cyCofNHePLcb
nSmJXLHjwD1IXGFHRxbQmHqpeHS9SjluJcP68SaVQcvJiBAxIYxMnKEJDu6wI5gdNp6enbRNM/Md
rskQMyJ6czUAflVfkVQ5mpXXSaVtqirXkmKatC0j7TTacoaMANO/TX/xQZvTsHJssCQhGzc5uTzh
fRp7NBSqz8yO/iqpXNnyA433HMo0zjnzK10RIeEAH1A5TttqK+06nsdwS6yVC/aGRM8Uk2uCSIYC
Z6PKnb9Ttztw5vN3dW7DCgkTblSRCuVs8pVBQsVLA5/QDOek2a7HJrW46ylKqV9QTXqJPe2ffhcI
jHwHbXRT7P0mzsOCX55txqIr35Tb1EHVEJTtAWyYub6z2Ow9AgIZiNXp91K+TUJgz51pQ16Xhpbl
2q7kq9+yUzdMF2o07UbWvSowsDjnSennOVJj92W1pv6D+6s7TuzAVIeOuhrU/64QBXDaS81ngfm5
yiti8+OdwzigOvtsAHGJvqSf+hIgXE5S9o7bUWcN4GMxjdLM2Lj9MsSZnH0QLjVy/5cbv0WgUA8X
b7IxBlUtPMSUGW+Rcsl0zekuu2mbrxVYNtdFx7C8RWvoS1Yvn8vW+TZA5ltgAW6rUyTxA2RTreJW
Yvca2TO73zv9po5MkS6L9r1N9aRu12jYBMU1nIzUJpuZhbxdEDh+tXuXKs7aEdNR+jdBk6tXbFyy
2orwdVeM5FzxptkTtEvQEsQNVu3XpJ8z2souaBbXRpXnm28q/xi3gzsqrOZCBq2ffxHOopFVKskI
pstOjAzeQNlr/0RwjzJqixqpIRrhZDQGOGAE+7opBPPl4I6BL/3ghY6OovXLFq0ssixenbXtEj79
rQ1q0U4XFbQbROM3jLtV0mtF3KD0c2LKPQdJoKd/uxq+UEVJwanYTWllCqBh0XKiLVN0RKFz4lli
50xa4odzsNNo7GXYNmXYPTQhgLXBjd8DOiehg9bTDc1isjkMCS77YNy8Y6auosvp4Rqey3c+EpGt
5XNXiz/53r92lHmlvxwgKRtFeYFKXBuy+tSpIesOcH5wPH8WuHSEdQ1T1gSqWLfwH2kdaIm3Ya4m
nTMAn4ez/JOY7utT9ltA2kzSAbItqq4mly3jloWmro8TxWmfW/pkkD+ezW4LMeTuZkhL1tyaABHg
NHuEEaco0htKHmLmD8OHyvDbLZ33HUCn9TB2cGpseTlhytNtpwcd08765MDVoX30BXQ8Sa1rZDob
l8g6gGLbUZ5qtqX+SLFe82v53Lix0V1INJuSrVOz0iLQvwuCBbZglQoHE5uywrE4RbIglrzOpHJs
SjVEm/S0Gz3ZvUG+/Sx9pw0R3lEX2SKyAtb+YWDZyuuq5Y9aMF7rmGDnuOXGcmnC+mjBXNwT3hB8
z675H+yhjjQuT6dZ5g03jFUYQVTQeLFsnUXU5UIQOMtvg1vRyQC3Jih7UZomH012CxXcth9ySrxg
l0Arv9Q+G6fhLch4Ph3Wh2gGBygSS0QRd764SjtpvcJA6i5AtYxvS/9V90KUuXi4LnOSjXJnZqLf
G7ZQzZzk0nzISyDCbVtG/uVUltZ3vd85ebeJ8WDouECuKkjSggtZRQmceEk1p+824HIHWK/zGkHX
JFDVs0Y0C2iyZGrtS7S3bMlXWphxfCNO68taB8vQFjigByCVMilnft2DMWQt0LvemjO/x43QIzFO
GLj6U3xFLeA4H5/iZjlF0KiNXvBg1mmDHAsMfTHqPw9PAmycEj5ukUkUCYPK7lVPxvI2+1I8cF6U
yF6uKRl+VdQPCMVoO8fBGJRMkcONxZzOWsMchZX0xZj3B3T23vRof9k+btop2W6xJ9a3IQIi33ty
WbbHRYP9FzLNyGoDdKc6aDrWLbUFGw+qYCLQaL2u/L/2yXegJuSHellVLYaHkde2ETx+ojafDgx8
NLp4rVlFGQ8Jz0i93/ncQYph8z7Trz+Fa864NLBUeGBCyK42nEu8oxUqYi3p6UItqg2Mg4BxnImn
rD0bhJKjtktZRyfyPvqEE/7PCf1iS5NApgoT99RW76fiJFt9qIHmjQ2n83YGSJk6rvZeTkMdfa/W
EOBtDUee6kgcJ78xCnMWaa1fYAoehIHZIA54lxISMjJDnZkjxI9iRiZ3KsY1S6JOPjZzidlJo8TJ
C6V2JYeZUzWWp7if5z2VlSuFShimkxa0pA+nHFqv/LPqcg8hECh4r6b0HmRs78VvrTkYE21HLyfH
MNShKl1WPrIJ6cf9aXrSb8ekzNnWNlcUdJ4+DA7925aAdb85SgMRaTV4TX8pm/eLmfxeTkN9FZcG
in/W/TKR6SYcwLLx8XQ0VPsnajE78pi07Cebcrom6XFZM+A0egeARmshJk+5IimEoyzyzQDthUDc
oB8DYMEwQS8e08vvLNTeHrv7rBKX0kxyiPmlVLyge9aCAw+Cpv9+wySJaY65j5kQhJyo0yOa3aAP
UXbo6hePVC8EnvTibYXy3JBi91neBfmBf2gtP/XAdrcLuYwnBFNiSiUIc7sMkWD7LkWP2LrNx2Hd
c/C88NKzMno0UMla4RL8gIW6JZoVqECr1ivKfUiS6AhBQhvX6hh7CHidN5kcHna2Uj04sXXdhTZj
9cb9JDWLQCeWYFmSDlAiy8132JuZuM4x0LC8Ei3H5rPytb5a30aaxccj3GwIBRvW8Rfp4N2e6uib
BG42zcWTLJA8U/r2bhagFQJDfw9xuX9oYOEqnsr9eBQa3HYUPlQW3rLGadF2o1qUD7YW3+QrBfMG
i346ScW2r7XqqYGa/tVKLHEp7IAHxEq5ZDiTqgJ4BZqaH3eb4eEZKpO0sjE6qXHwbkyhoImNTBja
V1SbX3R+UXlt1+Cmw0gIfTO0ovxnm/9JLV1qVZcNViNGPDpH66vcUmuu45y+a2IlTDDniXlyCHaz
EcsDWqDzjDsYH6tZk6gHjERUpGzVkSsxhfc4ZFcbuB2m3Y2lKFY00+kjBeNsfBFvqsk0dG1FlbmC
g2UV5Q0TELwTlP15EOwnMkox261NPZushJsCjZyLi1LXc6C1d4HoSDRp+qBmnpqjt4axkjgp91BC
XRQkz/B94eul2gR2H2GZvKprrlqwyG0G+EdtcA98wlMic+LCGF0CHBeWthL26owc1qFbS0A5yrJN
pWSkV01ITpZ12I/+BuHniTRLkwMiLgR6gnN40BCpehG7iPA3PlVKPTCG7u3d5QvhsbuRsLAovdST
bIy8r2l9e+YhCRvS4nbkMeSowLa/d7czVIHgLq/Ac4p3Y4SIE5ytdOXly53WQbPrBvkHpBOFcXdb
+tQA91CqlGjdhuf4PnKMp6MKUIPCK6ZAt5MAZFHBHUwWlXOpTiTLphIxmBwfqnSA+uRY439YFxzM
/NdYtwceeIbHOp7SG3AB4b7S8MLLkpK43uU+/NRM3FyonN0zxUxNmAnwD6XyG5AdrD7XoOnSpQNn
wQJRk25slHrGHFRo77qdBtydQNIpx87ICuGKj/LmwLVcb1T/sSwsXwnplcyM9VVgbgygv4skM39A
5SVYcnZOKp+eCyNoAH41Y+ivo9E0ZNv/oUPGU7lAM1ZOF7I1S/CKyXC3wAo/iMPnzPHMhYV4ZenV
AZ9YaVfi2YR30PqBP5nlktgV09x0+9JWcjE7ohWGGhx0YZi5RKliUErVCcVm5LVs8sJ2fsYLlg1O
aQPFzUnzNxAKNCpERT/GfHw3vhW6jKqdkk1q8cLPCr/vtqz0Csgbt95nwmoszrQsnbxaONdZWX32
n0/ihMnatjpo7dNeP9YQOlrgPZVMZu5ZTHppo5XfT1n2ndwwzv6A/lbYSAao24sLZMpZxQ1njoNz
ix5rbfIYzBeWdYx4Yha1pkC8hvdIYpBbyNV/Rs56goQPx98SF4Izw5ywjAbVAdacncmdHBvF2Lrp
By+yQk7Q3n7AOVLZESJDuidhWz9OzmdvUQnefvXM0jKNaEieuKwt6LFoKrtrfW25u040Wmiqmdq+
YeyIDkaG/HIA/PpFPdknbj5gEj+VO9IbBBV8bZ74EwtYYTJkWkUq01/3V9My3unvoGHHtmktEywN
BMJ+qvKKKu5B3LwUZymFw8jMQsRWSmnttXlp0gPwYMlfxJhh5od7vmQZIyIV7BGRMRoyziMrUqIc
Ntrm5nFt7AIpLaLz5e18X5LVGKtTZmI7vV4mDkrlGiAn874zMcNqwhOsvmedfiD0ZjOVNN2OMwMr
y7VD3iNjD0Jytfk5H02BffsB7YM1GAyeYH7qof15qng0yZCGsERlMf8PQcJWTMxMqXphA5SaV94r
oHjs+DA3g0sCBheT1nm+AjT77KBYrk6Ueg8AJ7MWXr/cPvaOEPauwqNC/9Ey6IX7xoBzWig4KpRk
Vnu177ol7nYWRLW5H1+5scpkZAAkL/OyPIXDprBHzWHshXvIa8t1hMVGDjoewvf36OBeijGdQ0zT
efhuU7E25EKgtOa+jGEVMRxM2NH0hEWddeO5VdtiB7DK+WrDW8SMPBRtO3j74UJukrFWYpIFhPyd
wb15K+/EHG3HE0N5yGOVsY8BT+EAAoRkOpfGLrouYsWkEEjDPnNTJn1potM8L4Unp86xix2okXJc
hhyKgzJCgmemWLjah4kdePGW2mTUGKaDHxUprzQEs2GBKxl4A9eOjxS/0Y/eXqWNxhDEn4vt6Drd
KpV+8z1+KPcKdglqGbXj3JinyHtfWSZEY/jg1GdwBGCZGk4R8k4d+bMXH6d4Zo19qR6DitTzUCly
xOHrHUzmmNj2gwqmm9qPspoaAzNtTE72b65ZaL1J3Zm80eW8WiVxzRHJyG7tyL71LzWofpI4JZXl
XduNo4dcxMezZy+sSWl6AYbcpFCcRH5/eqcPhcx5S+UfGyKgh2R1ScUtFU0tJNxz7y9GxDQn0L82
tnBm+wUEPVpUfMYhrtvUrqZhajKGof96kzOzp0JFkKchTICKoTunf1VmeRW5B0oyeqhp8GWuki81
1nYwEqh0gWwjOLQcQhRU1WsbNBnK/4M4LHwz70HbCW8RYO0XZgX/8iNpFYV1WyWEY/NnQWP/Wcjo
43WtoPYgkd6Z2RYuxsv/xIw+d3+zxHgh0O+l8lY8NFlcZVENNJw1Jh9PNub9Rn6pdzb9avxD7A+p
9GBItRn+DzaoTejWvXvcLto2ocR/rJnChQe31DTvdhwwxMjHFuUyNRztxFTgrR2ALGCagUbADKe4
rP02VcGobqfqinSiKXnZcNVyoWFqdyEqTyy4dIwTu8KWKrfGJPwNPhPqp40fHRYXpiUlZltao7CJ
gy/h6N9cod9kjhOhyL2Hzq+xHwhMhm7g13Uhg/JIr456+UZbcPngleacy+wRTWq7TlgSzujN/zDn
+YSIo9w7v78GuRHA8xBRay1zWRMp8uXi93B/ZBJrT9tdUKm5l7Uw/MJmHPC1PbHF9zl6hd1heLCc
wNBMIAJNXaUGBUV1IkNto9svnPWFxizvSwmZ6/tNPm4vQ7iWOI1PN2xevXfHqyp6sbP+sQ4dhG3o
Zr7TAprOaatk72fWybFt44Z48fe7kVD9X9XQFV3OSI8FkRrACRpRvMHBzobw7alJKFuNNlG7AK1W
X1jPod9aI1zZlr7Aj5JRXE1RqTxiDGjwNEgFUM5mjN2h3sPQiL4kKLla5u3xRHWPC0S2ant9+cEp
rg3etfc2r9vqxxRf38/otmfrRJPYjMBvKdl4CCeg47qnfFxSVqp7bI/A7bIOX8/Gi2WHgoZL+eyN
L7Xz27pOcZN48khM0Z02PIujFr3GEkIVn/GpaKZJxwOxqRu5k5wCDcTin1r8sPy50hsdxj8WnmHu
BxRXhrW2xi3DXDiDt8wiH9yaqhAb8QSxW4PhQke2+OneKVtt6+MkJU6tV+j8qcjcOZndwJDraqp5
OkhUagTKiip6NusvtJCYUMAE3galc/8GRg2QAywjU59uR4pma1vxMV5LEraWNJLqRXp/OqgRkzeu
6+ythK7cnFx7stDZK5xL4SC/w5E9IFwFRlXSauUqhAeUoiVVGewo6MG6OGy8qwK/km4O35JXdGX9
tNMLUWcZp6O7waMoVrd3zAZKphR8Ln0nmD9JKABhbQa9Di2Q8HxSq3+d6XQPB4cWfEAIqHbkKP0U
c+H/Ff3wuQXKuNN0ARiM3U2hO269rhbv1D7OdhM8gybcra+tEsScVDN8sF/9t1cXQLObyLzi52wB
mRYgwq/EWOK4CL2sWbQBR/jMHuWBrPIJANts6YHlFnsJWqFQeFEc9SYFm13jwDwqFZHEE5AjKEdk
S0Ipw31W5lI8lDomMI5tudk+k698xuBPP1iUAADFX6VxyW4cOsdMNCluyB+wLzABGygIo/V8clzH
Urv/MzVudLYfCqp6Q23RUxgWspC6SmmLjvdrIoIXi9EmhCnkCsFhg9n6Rn1uxspZ/NT1MWyaEkSZ
BeoKSW900SCDeXUR54FFBxZxWckZCB6DW9AvXqe1j20G1jl1nXnNR6VwKhlxe6FYxrL7zm264pWi
NaSmQTIn7bee4BI6ZMqNFRI1eALlc/9kbnvXK215k5WOPpxbXOXK8ljhCSTayKubIuE3l/UVC1MM
Y08EDEZ7t1HEJxM+3hw/HjDNvAZAWrkqKamEPNtV54uAKoKBdFy297qZOIMMpZn0eMuTT7TDAIsC
zr20gjR/MaUO5nRr6D/sJ/iuYCJSO0wMVXkX/DK2VO7uwqtUf3vktAWqG7WSTNB+zAlGnUfqZvuw
tcL7ncc4OVGDxRo6oPRkbvAeQKKV0xi4Q7l6/zkfA70P6zgOcQSoAmU7EDaYthd2ByYOP+0y3yCR
vzfh6hPXv+Eo4t6x9PXgoCCoHtPefHwQ3wS/B9EiXYX2biEPtrl7A9gpspvvwnvqIjydEXY8UBZm
39oVX1ah+GLwrwMU4bl2UHsIEV2tzDGW1i1I5FTqhawsmQDQfq89w86BFfBUDh0cg4emEbDf11AD
+zrcG4UacsOwo5Z2cbbYZ53jap1vVhA4DiPjKW45v2zMMyFircSf0emL/c7+0VYB+xZJoWZ5uRWe
pIKs1VjUHxO7GL1W0919drMLNBw2xIDvqhEW0rcXFV/WUZNjMtq2FohgAVT6vDZz9OBY1huESqUw
McclqBhYKJjfK48IQP8vk7y6svzKbHMeZ48h8NxtEM/K4uE4h9XJuXbJ/mv3YQxKOW7auzrXhl6h
XusDV37zEL5ge5nFVrZ63ssfV2M7bT4N+XUB/NfydMv5Ux0A8nLFXMYUwJCq96u4JPdKB/q3IHA5
zI1ECQ/5LM1O3ALM/9q7OLk1rQm6WS+4A0oquuASTcSDXNa4M3dULFWbeXvULSa2QLrPVFFYIXJZ
/dvop7aKv7LaTLjAvNP5yVoLifLNGAwc9k3S7z/r5X4wB+B58+NerDnrxEQ5dCgAY/MuXmDQ4iLY
60WuVkK31xrynF+UaVMieDSQTp4L1zLnOmHGAdgF1KjtH7fC1Lh9Bn3oEDzBzbdkX19HCWNENNtc
10fn1dqku+0yte9eR0xkmvbnmivSOfUnPdR721wXqCZ50jY0uUlXJbPd0GFvrJWMC4Wv9znCk2o1
gAZo3fsTTM4w+WHTfcTDyvq5x0NLmrC3W2OLNPz4KwZ0W/FH8rZl2WStNNh3C0PY5fZA60Ew47xr
Q2O9HH/yGZaAqu/v0Vxe2BnG4rSNFeqMnQxPZsAZqFwoGH2pfR6j4dFkOgSBShqAmZ0h5MeqHuti
9d/xsU5XZuTtLlCU6w6/DU7m141OX3BNz2wiyLadBTh97EFb1b5CsBg7rCYMrT1bXP+aCOXB/DIW
CQNKZoJowtQMILGECPOxNkz0R41agi346+AV5UvQHjudtF3xXMd9tIy0sKV7mzLuNqXyPs9Qgtic
lUGan5o8NOQbtZ8C8utKDlArmug94l1Q1usgc7BG8szzvqUqQnvA2fmmlbMofnYxJAsVSZAAjLxb
ANo5un0luiCygm5Oqj+1CP1xnX//AurvREtc851xwLbiinujW9WsJ1aDuRQ+vyiCV+3MHDkekpD/
XstquvJZ6S8rH7tl45EhWMtmjGpBZC91KC22SdtiRynYqvGKiD6DrbZtCoNalKrPqJ1kqKeAwsuT
y1RkhLQ6xrQol6pjCf0FnQy1ed+HfHO5SJQCHisvJP/Ja+civyyu3Y2TTAMWQ9HjDBExXAWhQD2h
DmyT0VVNsneGiHOEL5Fg9EjVuoKraWMazC4jO4SqTueh251KfvVqDBdihW7D10JiKRuMLJ0Uofl5
xDDiPL0RLBeaBgWnvhl4ho+uv8p56fVd1wP3zff4ew6BjvA3835fNjy9iEE3sFkNwrFAGZC1BaQA
M19Wq3e8KR+U0qyQWkUwfhMPqvJlLXUE6Ty3y4MYUbaEZbMn7d0/iyIhxgoYeabbjQYoQinM9XbG
NUg2pzyki2+tCTyaVyiBhEhnoP8SPITdPkc915wirrYViunuObFSQVXFzMALunxosqm9am7tpucS
fKgAWSqFN0DNFqUOy2rmLDEqz12ubQO8Sz4+BxXrloBXvRdCskr6PqBxdo8t/TGr0pMd/MzBaAxD
2ZO1bgxrchRMED3F61OhjQUcXHMgzoTSsijk7RFM8QJvvIKDSpebRS3QNxUhz1TUxd6O8xC2rguf
7G8yikXDNQAYL1d4qEtqleyQPaRl9GT9k6Usjg7NctHGKgi6TGH2H8Xa7UuDLZxKnyvMvbgUTYqU
herTzTAL0whVzVdfbGEFlTwj6kw9hGWeeszThZLO1WVQhCmYk9atJuR8QV2teWPxNkAmcOAJvAL1
1qFsnkQKURzCf0HDxwDNnjLxJApqklEj9sP09d9t9WBkkc5CI+/kHNilGfjf/M//i4GkMl+YQUCA
vpyHbEAJWL8WzUAycdvHaNWzUJOwx065/EjCsfahHDhrqFhdFMVcsk0pn5xjlhieGzMVKohuliqp
v8Q2Tek7lMxk94UeVpz/d7pkPuGa7ddKFXjlNzLkdj3fMfvW1qUdqFDA9qUg/HeJ0xCjHAfexAEH
RvkM40pbdI7YkIW9S60RuBHHx088gp3GoUdLsaslPIK1AUaQ+yvmaTuqXck9+fuMyfAg96RZAnXP
8BFkRg3Xh+bG2PIC6hsDjSCWBi2ymBWm9QPwRrDTAVZgSg5He1gXV4tgQWADZH+h448O46GavbS0
VNODu7Re40QnHbs5286tShjG+qVfxFVFppnQoRB/UcSNqYoQYBvTKbsIOwkQue+cEzbmQG4HurNd
GEpbSDHSZpAWN6ZuqTmNX04tx9iNNmKrEx63iSFk+CpcaZ4KGQDasREf6srUpiIA+9KYYXt1DoEG
/tjYUS07T6LqNqWji7eXUvqKffWNxJDkXbXKBwDDBONmKaGYPAr33qWrbKFhNDTZkMmzixlri7T5
QLWlVz9enjRvH/SQgWuOZbgBiVVMutrKOF/fhCjfRrA8fj1LiYfeTwHCb1+19njOZyFU0IAXXARE
9Z5n09VuY6SjUx83u30nwoU6Q2AM9+kRmhpsBljGuNOXB2K7ITy26HClWZaRCOQuoqgaStd9eNO8
Uf2jez+vCCPDN/KSW9hS0/EAiUSXw04X34jUN/UzntWFEBt5stH9ciRiUGF+UkodYtLtQk5d7bK/
AEfRuKQW7jCcM1msxIJCKb/Z2eNqyPvKv51stlWJz0IEbNtqwGwxOe1lmejG8Z8/UNpD/xb9usj+
WDXIqNz+xNELK2zSuQrqAM9HUTqdNIIy5f+eQP5ZGX5MLGMvS6uQA7tcP3IL+TdQbkLZS5Y220Qm
An1NrtFyJ9tZ7nUENpyx4/KGpOBs95DYsZpSmBix1MZOC5jyWhmmFFuFmb+cKOpGtpX6F7fBh+g2
PqOko1ka1w/4wVyeHv4uv9IwZFPa6p7tzUEN6yFpBpRYDXjlybhKjctDFYufgYsLguI5bMWqrbGw
bPZTfIJfm1W91TlSu2FqfjkZIcA0HiNR7NAcqYO46o8Q3mkuxGLN63NVVLDtyjyG+SIe19+PTzTV
+jlGbNV9/84fx+thFHv77TGK5rX6l/bzkHfJ6bRBxTgVpZLJP70F1zk0/0K8bx6nTc8mLZXbJ50z
lwg0Kn3n4tvM2H0NjpX+5/PWlZN4B9hZGN2FGIeGBc9FROlO6C/9u5beVRKMn4tIJncok7YGlFWT
w2StVYiOdW12PPXf90cnkL+jTHwH780TidKWlnbrcgoENkmGJynTTZ6wlcyMmrXB5Nr3UhC4DiD1
PapfBqd9RrlebhGf520MTgg47xginRENdAYvCkACs/vjaVfV/ZkHDL+GbZfW3vnrrradYRP1pFUm
1C6vDr+VaYYALfFNZ/wYeAiSU6vQE3nX7tNevZDL+SbvyCZeNiGL8cJAEfv+v+oBhgtm9g4PgZES
rjv4oo9zDJBlLTSk2PJ/TUPt1URvjVIP/nZS2CfIlvhFVzVcy4+ZVh6E1qLIJ+x09jv3M4l78IEm
uTVu0gN121Gp6Vl6JSamTT8THAUaFLDiLoXDUqxiS0fK0OpsDUEmxDYPh9eTT+EdUOIroccZKkq7
M9fSb9f6pUmiZQuEim2mNseAgSDd+H7Qj5hf8SWcFLIqOlKnGj8WjrEy36BFj5FJQisnDUfBSHQb
nq7NbDc5ri4bic8F6ZvlhcHm7z1894wghHNcA4KBcvDys5nrlELkDCaIKHYlli6ivOmx8pFWsEfe
j1Z0jfEGf4Wm7c8nrltrXe8153GJEyFF1AulydwDneBakbTmBIpLLdnEZEiWntI16ZLN4AOBidyy
aGzIZxWSKSoghxk0dPntp+I0qB3qtwkGqAdqJbLVHpbI+Ll4ricedDhc0D74RThtLW0C2cAXYe+x
vkwwa2NFxE5WEc+kZc7qvIiQfjGa13hAt9EPJvj8FguYU5+JL4wSfqNwnqfgH+IYf+Tg+2dGWuUi
elsL+peV5QXt/qif3OtQT/Giwr9pBgtDAKon8q8ZisZJWJY8hEypBpszTzw2be6aDqf8LijD2nz1
VQTUiYR7z8OWEvqKsz7CNLklGQc/CQsc1n1mK67K53tLfweGSUbAMfPXnPebUvY0gyDTrRuUk4EM
V5y5j8T3XzgAhQtEcIk4+TZWWe7uwQTeizYBmi+p1WYp38Y9ee3wcZbW8fG3OUhtzNcebfI2XJqz
Hd71beDI+NU/K2vgEG7aM/82kZenTeCKKAH6NlF36d9BWz92v/VAdGJ+oKTJ99LpvzRFM7a7YvWK
yq3uU3uBfC+9tfKP7ToImvrTS8hE5aTe6yHzBwPWMRK7E3oKVMkN+TNhyyGA9rEMEJr1j5y1akpW
otoJgl/m3zKMqbOKNSsZAs2la6n4k2/+kppF7lG4wKNJ/vEqiZDTIECM/tQPYSV5Qys4/mceBHuB
Yz+M1f7SiptHI57f6JAqN8JyJfkbwo9lDl0PxYI/w7ECH66HNeOTPu1gTv0PjUahCjy3wDy9m1RC
Muoj2YQJ+Lq8mYOEs4cpnMqWcvyZzNUbna6eKwtdJ2MD6iNOeu2WaXUTvBX4vJRLnk+qkUNW+RX4
qBP5Ubmb+OxoS16q7eRgKQSQmQe9XD41pNyqhYXUu9bhz0NgneLPvVs/sBE0El/zSS1QHQGevlQF
u8uwg4l8hS+/Oywi+z9rzdSQ71P8K/Ef9aijl1srYMGw7RM3MZsyIyx3SvUPYhBJhbFR/1732aq1
hwzPhuQyUbXHZMD+P9A6SA3UE+2l40mDAQa+imlO+flDyKtSpIGHGSalatAG8qKTeSNVTFSL84a9
SRL+qRpHJitLujSwDH7t1irc3JXkuGLHlSmKatFluRCC/k8krEHITnBPPE3tECE/cbynxnWZOYXF
zXWPXww1Xjr+CczEHBgbQlZ3MXmRJzFM7zyPbROCdoCi8KRAa6Ym7EwDu04plsZ77XgxVAZAm6nu
f3SjK1sw58pgY7AtdB0BFUXiQswCmn3UOUDMx6w0jHsG/b2FimJxvKy7uvBLmFqyxuid11tkNfDt
vg3ZCjpTYmI972rCkemEHSooTRZiThbEb6B7C/TtKsdFrPdSJEFnzyRicYuY2A17ZyU5eWCxeVUq
m4Mcf44YbdrtCHQnmXUpnA2EK34CbKKDWKFVYw0Lnltq5VLFymYxb+t3qNitVNAX+0lsYmNJo1e8
M4Wv5WQWW+z31uxW/4LsFS42dzEIEJSfTihj88pdC+y2+bf9ilmVVyBWwqOUA/xhKoja9IakD4Lu
xqsD6hpFwluihbSkW2YVGgaKZ3JtgysAjY+FRKhubdqdWeoo8pvjO8pmofkhutskgEOBEN+vNFbg
kv/8m7gXQ5L4qSH85KcN53f829XYfXVSyr4s5j7eQeYdsu/kiM2W73RMJRgIVXi2ppMz98+sOTf2
WkaDxu9eGJ0+Wl327ipI4kk5QzcqPXYz5Q471EBfUQT28OOsQt6K5St65sG0kjwL5mcezuafyk7t
Pgx1r/4UoVFOiq9Xt1e0avCLjKz6gUBtYVx9y+UknoV5uODqP6lShvF0HPfBXSBppcReCIvxkNt8
FZ0O2Q2h2iPjyd0r1snScAhA23cB/7rAP2BvAkihwBpmheLoe/1zKYZthvZ1LwvEp1xRAHo1efkS
pPAwnG5/4Yw6awf7uU/+qluE9caGGrZXDaixtPxEhL4CSklIKi7MvwsAH2jv8Nz5MW5mqvg7NBmX
tPS2WkM6xeP2Tq9gQ4JiEB5m79RmYsuyeXFtPVW6s2GDaPPC9HB/kYqmWbVW34rxhfBbCoMUZznf
9FVKzDto7euaJqkmte3hW41FN4VddCyb38YKr/dtgvQ9DO6aYFW7alhY6I+30s56xfp+bD4dkMAD
GzuzbKT/wwbetVpRtJcQCt5SgY7eaSB6uFu5VcuOqP2UAHQv7+lpLaEvPRRSFZWek5YUhYW6zu9A
losp5IfnuAfRpeBtJQqk5rsgI2kR7jK+G+YcEo3J0KxoccEUiMF2Eb+zgBRii/ibO5rXtaKBtjBp
lRJMNEbHjTrf8C+w2zniha35PsAKlQkMitl0owR30aGPiRmIY/b/yL1j+uLR68gluZbQbtAx+BNw
jaJO3BGX6LeIuTNL9tqIuCD3Oz47cWvtd3iOrUBVU4GwO0CmX3SE1EAegziv9VQD/0AFgpsCQW91
GBWWOwp2WWWlv9gmeellqipg+bKn3MZ79KX1/4Fvg0LtYeLNhRaIttoDnytQHctANV+itc/JXU3b
ZvvVfbFn21v8V8YsjJqpfinoEnMznSbfMLv8ihxH1+ficwCsMYZ5YVNqiLR5LowIZxI04Wh4q+jo
3TGAhJ4tlYgz+HQ2EyCRwKevKhy0XFAo9t3sVKC0ewy3Rrh97WgebVjMInYEnyI811ePcgy++GLt
Oq3PC+tJRdPFbUDHVs+Ox9W0drjX4w+omfTVvLXqpET3lfuzBcfo0X30CkhlfWtUYxTZBvXecpN2
OdH74far64VmMSR8HBRYGOoXHmrgvsTdrbQzkK6mCpk2qHo5xMidYgvcP+wYrLDKtkBLL2zAV21S
rGTGp6PiS8jiCKgEVi4Xx+JzmS2wWNuJ4Cnk3kGH4QqDoZTlcz8KOiDdMNKi3YM890rp/q+4guJB
OOc2sO2XtyxzcIjqEsfKVq3oKAH1rbWzcJqzMe1FCQTFjZG34Q4BmLI6bGzrLVqHSpbobMP+F1L0
iPpoPhpkpBuyusQah5hTB7RsSfa6r38VdAwkEgGKBagEakcnfdNuj6UTVFukGKGXBghaKXCIWKjF
h2mfGeS164dl3LILJ32fmkr3lBS77hNxByI3+pbrM6uERIz0XqEpnKt/L2d/t4S9+M41Ne8luMFv
jTwtPw8LvdOHtVCST/eTHmlMAYA/ekm5ArfbzEDoHtpi+2cxtAWQ400xzUzoxl8yLWAj6Dlm39Hb
IJ/OePrz6codB7psLnrklo9a2rLlusFRHp2LYTRuuoryZtUfBqHU6dGYgtBgu9nx6tW6dC9pQ8kP
PruXkPaov4mvZN5cSo6ZAupTXCj8rEbu3BhVo8g8Ed9z/TD7wzguW3eW1PECpxS8NonPFb6Igw+O
rUa/9BpJA+kT4ifXlq0h5T0jdkh9hzFIyB6PS5HtupYS8TYrf6GAegMgT4YPMp66rtuVmS5NlObm
wjUn4BFO3t+bjk8Fuoost34v+dReHxapLB7WrJ6qnWmndfcMRX+iOXNw1y14Bz7Czi3UKVqHYNnr
HyyypkftyGkdP4ozCiBlsGlezu6kyThn+Trfi1h76GilwxJXRJlqsqhkiu8vydEblZ5yo8u+GU5n
PDkP6b9kYkPnHAkok4tGbqHC4/+/5zqVCt++XFjSpbn8Xiytvk1Bca3iSec37l5WSjYZY7JJqcPe
9mkr931dloemTPM7LHHJGre8CW0azmMHkO5gyww+qNDYwnVbrniulNzdkIlTCVqSg7BZZcKVcxRY
z/3CDK85WplMBQwPkzOMaVAgC54X4TG0QkMhYJbVY6+GD/4CSF30NcPQYbY4v3WVMxNt2y66Uxji
NOHp7vA3H17SM9QR7MFOTJJL9kLC7bLl6gz3JSVzYvZx8JIuMynJQ5VkSF/ylufd68VDr3+XgNMl
mSmwur2Ks/1HvpGrq1N29eXyy0tT0yaGx+Ki9EwF1IZ4MuC/Hs3gbGPd2rfo1Fz8o5d3faj2jGpo
CYYeQvLuoRVDA0br+gvT0kriRVuffzvkckEMHCYgWkm4wq12smW2l7AsVvv2Ze+58Alt3oe0XMH4
YnZqlT39L1lHpnFSo0U1y6sJsS6xSHwB2I7tsxBgmbZaMxIAjv5jwZ1By7arIBIuAGLjGlulSLP7
zFhfQwl5fb490ID2dHaTai3ihoEY7pbH/2s+2JIj8VeWSGhmD8IACDSVRH4IFf7qn95WFJ47UWR9
MHaA6GrOj12ydbvQUs+3xNzTISTfK4JPHQ+e6F2LqIzQMOmtLHiIBbdLAweXHKCild+Qcv5qNEJQ
7NS/mYV0qW+w8Zw+tkRrLvLnpo0nXKs9UHBnrBs5sFoZOphJtgdM/+4LlMRnrcb7BM0aZzA5jqDM
MsNCpHtcR2uvLG62FoZxgO5WJcYCfCIGKZPW/o/tVDxplBIdHJL296XAzU8s8GtqPHaPrsuFQ1bA
Un4NjC+Mr/nS3DiI+MJ5I3jXHUrbulN5UK0RiMsiCKxy5Re1xGI/bf8gEAFy5rKWizeXb66rXXyI
dDtDBQMJ6MNEVKgqurpfOwjnxJw0qIhGRgVK2eoJARwTjn0CyV26lSD/34rRO4QL5eJGVQfkoQVu
//uAAPK/NwTB65vTGk4qZ0iKO5Mv8TlPJKX3TbkILJk49Z/mk6NXqUidTlxwWB6p5pmarVaiCBUl
D8SPBmVD4BkogXBfTmF+jpfc/4Qe+V1ofQjQMTeFuUQK5uJdnfrZX+L0ec+EwTSLCvPUY3bE+Q9/
j9bT9HpS/BmRVZVU+DV3u7+MFoquBcIO+q8otPpkdaISGHwSspect6W5ymI9Bgeu1BeaEY+mWo4L
VxTS8a2cMbWWezXEtIbKulQEt5baaSXdfSG9X39V6fwPE54442NJnG1n8T8q7HXntuDavG8m+tIB
J0KfrxVwFARLT3i+xhqUDsKvTH5zRhKE0ZpGQe3C536S7tX3L8ed0j+iNlozAu0ZvFkFhosqdZH4
J+eBzdI71ZLwMi89JywWbd2t6jts7mrrhoeL3bf50MRO+Iz13FlWR8PGDEkfKrb5vaE9HiBtuY0L
a2TBd6aglcg790cTf4y3BHV7ck72vPtLJCKBk/qrhxN2Ci3MCfAXLR0XoR8rvPdlNIYo41sCOYeT
2scC+iCxoL7rsbdMHqb349BQugx9obe2PMfLDDhXhRaq5DZNoA5ldvzjb6pGW3xPx+wC3Mqf/KOK
Ln99PP8/Ydal7OTeTmrgFQlkUPtK0l6OjEWTtlek9j7KrkE/d3q/gLqyl1jN4fHB6y360ZO0Y+BI
DOAqqg0ED51XIY3ij3UefELTQ6WtNxjxHkQGAhnF1Pv/JHbfkL0G7zIg4Jos2Vt83zoKE5C20zwH
siCEn1HCDl3ZKn+KokiX9WH2xKKjvPRKtb49gQGzIaT9xiUDDYjWsIyORXkO7ZG0ZPNhz1Tu8GBF
KCMiDH85BcQdFBX6LKzTovsn4Kb7F9j3fKahJkNhjQFjFohlaloyb09vJwckjUvUGiHXl+7/oCOI
qEEbvBf9HWvB5x0zSoWIhqqB+Ug7UEr0eX7aXvJxfOAhcZUXsUK6uUD8LP1VMgcMCkd0fN5qVnsj
OKvG+lHrtwPAtLBbtMEl+VMBXL30N3GLL8yYYMh6qic+EjpA2DhwvBssRimvDkzeEjlTj12/tbLh
gveEJANidQqmzCc8dtudAJss/iaGa1YjdEtCi6q1HTTBdk4b8nNgT9pPRiIMzJZrL3NzQd8pRQEF
WK21nTdhy/LblSKhe9iM1zGRyoPQUQT12FHLR083ioRlwDhXSssS4oXXXtZoBk9I8qDFx/3+nGgV
Rop784NZfAfuhbxl6URV9PUf5PZQX/z1Z4Ev1AHW5l2hoUXZVYkNXHMznN6yDN8Jbv56vsOlnvOw
ZlFUOM0RwiUJbbZWE+iZspmqOiErkLUYrmCnBCvYi4P1v1kUV6DzYhE42SPxhYbawtcBvn1sTGPs
Qkd2BG3Pqw7iE4LLQ994/FzcUEyYWTbQRKTmPeO18ScUy4ItzVyYIerJdQVcaNajJaSUsHavUhq8
f0aXrGm9dn5D83OVsyrUFfC+uqKmg8wjtH3g/rwiN/MbbqTRX4M/kLuYlD/beQE9pm5JNhOM0jcc
4XKZRdxZqdK+RHnjXKQFbGYuYa3w4TVLIl8FKCzb02eXhvKpmBVYAH6dzQf1cxpkAB1SuQRtt7Iw
NJDPglwALUkn64b6cJcTKCZf1Bx3uZJhqHWYmWbDdaNgZZF/1noZ8eZViLjLnIGXmog5yTekIqlk
P0yomjAG+UsQVZQpifOfjKa/1XkiAM3QspLhHBN/I3agGhhbslcJZUCNQcQHxe7z1fFp/ND10+SY
HyU/+YqgvXZpQz36Q9l21HFaDTcnfpIwerhMaxLX+Bb3PX2O4Lf0MyBjDBrqg6E1cp8AQleA8coo
UODCbY7UWnmj5Uvv8DP8PE9kMbSjFaDK7CpleHWNxRWCDjildD8EuQSEeMMjpsJNmK4zjp0cbNxv
PmfnN0vM5S+mbYuRYzJxHQr2mJ+CfFh6lkA4k9gQK2BWYlBWw407vwcPBbpwc0sMEFfReAmr/BnP
CEzqf6V+F/a3QHcbSzcYE9ytzvBfokweRZZ03ThxpNCpjR1mPgQcnN8gJLK9i47YoWA3rAXh778Q
f6Bbo+sPFbQTbkk/TJKABD1s4fLEWnbh9m+Ugt6VSETO8l9KbI6LHLptFKroIbVNLFChy02T6J84
zitfKHHs7vBqMAUJWcct3PwMH0BXFGWXuvGpXsDQU/4E7Y87r/M7bHofSZIyOurhG9FIWIW8S36s
zRIo5x2NStpB2iqbdV4b+MZC88Fz1Pef4F4peOjgmF49kIjaBFOkeGIfxOpf46q+1CRi6tC1pmMZ
dCHHRyLMe4bDV1Wab411Rukn0nmG7ne2xS8UcZGwA5E2DyxbjRO6p4SWhhZtqfN6s68mlfXPqzsZ
ngYoY+jFbXG3CVHJ+gWzUncnTVaaIm4Mrc3XVrg7HCYCoeVGl2nMrmLwOLOeFPdXYOnHC7I8o09Q
Un7t1fAm5AeMswkIBnNpvVf/1w98JgojjH3NHkXvEgBQcyfFvCuJ8KJgYa3mnQbk8HmqT3VSGBr7
IguXP1g29d0NneKR1fpaAzgHaPOCpwozZtDjwGKpdD081rW3k1YqYbipqvvYTs14sI8ntQ7CYn3W
4CVWd/+CWN8Syjtn/t2xqkAKQWfBUwGDyVRP4YNTSv9Yqx8MsumZ/AkRJDcCs08qWTWiZs+hsg2B
/5A3qfNXOEzKXIAMkGxAUpUvLg3PTbiDrxffh8tTQ/4mTD78u0hCuYs6AL253yAV93zZwbhsaFrp
G7WvgpuihXWGdHfJAKehumklWYwlgqIN+5jxua7L/OZSRvd20+qMxJkcD9WuNr1iXKloRACMbG/Y
OrzdbXoZPh1XjUisMRaEYg5+HnJjysrGkF/wd/h1cXocfwAx+CjHRIIoKFCTlIG68S5YbTI8Um4l
YwioS1GHi+SVfoEtT1+rQtEtflTNlHJjG035HXqGdJwMCFYgGWCYUkgjO41vHKnpajoSwhQ+shqI
JxFQKE+YsEoFmkebFeVpiIUwNG0YfrU8B6tu0qUQqaDxf20/2VYM1B0YadNt08A9+NSBFvZ4mBWa
2swtimTkYVQ2yyiWs3yXKyyA8KIlIaIMBAh0k9V2FKJv+jSC8505icfdnIonCZNYYlgn376nxIRo
XYefM1vm1O3vq2MrhMZUYZ0Sd3xPUi07VRn1MQ2ezqJuOC7aZgAm/9pZ1b+Q5JSFjg8UQ18Tid6r
FGyB51uSBUW6zinVM4wEXtbVhUhTK7qS3qaQbodwLGzqpVgBz+T36i/guNd4m/CALRqM6mz3bGXq
OQZ7ervNTvVNawaZ34Ig1V4NX283FM6vQK+k2QZb1iODHV2C55WmatpX7if/DugL1qg8Aex0mneQ
Z5/P9b4E94q5xwG502t+vOIh4eK6v6UhQYPrYbTBKTxXu02VEcH3Yz5sEvFMrixg7fujVomncDNi
ZsTqxcpFdN75mDURM4kn/uEIAOynyyBN2H2PqIend25zSsOFZ18xvU3lNzuG3RFqdDFP4DrPYraQ
jg0olUg/mjofNeQhTD6995v72ejaggSkaG6N0xvuOMS/hj8n9utJ8QylyBPvv4E1Ndq8fhALy6yc
qIWv4ojK74EEtd8mjgLcJ60IpaSjn3ckro+iZIwf9wgcuHSaATU2wRviIrhwF20qwmhNFZWvwpZh
KgNwsFwgadN1Z2amZ9tyZOeG44Tab74fyh1uGeiw6O2NJPzp1fCWrNx2bY8gJki/9qRl3aOTXJmO
q9usFpPqwkj8UXU8fU+GJTyGqORZAsJUwhEhltz+3EAzSoaOgQvPdksTtitrvz5wW7HMH6f8xmax
O4l7vCukS3fpoAO/xZV8Q/sOcFdZNjZyNQdjLK2vE/pOnIuz7ab8YEbRV2ZrHIvQlJybzuM+Zmx9
nb6hNQRDPK6RE/Rpp0dNqIwh7T2041pN7vJl7OYJ0L5bP/roUmOX8l/DodT0kyz3Vb3uheqOC4MN
89QnQuQUFpFKL40rDd9ANNFVZrutsiw7eSaxsTEnjaqadhesG3G5tWy6FG8uB973uB9wfUy2ZAE6
qALuvNIGjbIXX9nP+c6gAoiiX/eGLQDppo5zzs8IskYt6+cZcUFmKO6tygv7JfnRKv9LCD+JfPBw
v4STHEBS8yFbsAGw+WswpYNKVtWhjuY0l5Q/x2vgROjIwqKOYPxO1HPp5hIFhTjGi5mw3amvfgbR
Bf5OqEXgDMDlGGXydDPZlPbz4mSWH7mr5EgK71cURbi5zzd8llX9juuP1i/mcjcJfeltijIOxTTi
+pYYySTeF33yHGJTuW1rZfQxoX+3UpvaXLHzfAIu2JcTaZQjJe32oBP8TrCtcF9E9qidQAQkRcbC
CADRbjYd0txQsjodQrP6WvlZtgmv8JAsoae626n4aqov1NiHlfgkSlySElgpVSU78Udd1h9Ei7lZ
UYeC2/19+lhbhGgEWoHpyuPD2fnXIWBtAilA6/d2Yn8snLzrQr4mNqUuwXv0bfsI9KEDE1+mFQoz
607w9fA0NQJtX2VRVMbY/8CXpv1Pl4E5JMkay0Di7qDlgMs1wmysU6cYhPg0gah9Xi0YVatX4WnD
kaFRQ0LQXCVEfybi07nnuGbwujoPaybsnYjbE9VVOE/F1xk383se4ox9NHx8z0TRGLhAknUhazmH
k5TWFtS039cwtkU+9fRYfSd2ajL6RYtM3EDoxtkwqUCHtgt0IVwuSdDvTma75jy2rvJoeMHig+CU
ZTz3BvSP5QWVxBKo82cixPvCBNBIiPFyNR1cKlOhu4u17Vxw3qq1qQomadMSncSHjsqVP17S4Jjv
iib9nWFh360cUgl6YN4NuaD5iAoQoXV+ltpo4L2Sho/L6A2Vzs7dzKaeJ6hJy2cYnEeMaD0lmUnc
EQoiq9FpnSMOByGH9nCm6jM/nS4CFRGW9/mWQRHTX3mFs4tr3XNjixfabVGfquppU8/+NHw3TKHg
PacFBApFUrQfh3BPaub7O8N/t757FB50DiHJjABdcraicF3/ICqyZhmkH2mdhTN9yq8XzpV/0pgl
3K9Dv95G2kEwGR+uI6p0ss+jHzB4w1c3H0poM5oAbva6EsMiONvCTp4BrtYJcW8F0aPlO5v4jdBG
Cflogk4YBNud76/X8j6cuWDlHO2fMq5cQPCnFlhG7fpwr57zPYJWU4eXEaZZ+JkaSK/uNtMiY0Lg
wFQ9fMpNZpTqniihf1sYgbL0+6TzZFvKa1cD/k9T3GdhwkmEw0mYM8P16IpRyIklpU7jIIjlV6Oy
Q60ghJVJiB0mhGWarTQiYta089RGrnUlIXbsQbOdRh4D0yVC/s+zMUECG1UPRvh/ar0e7o3AuJwC
gnkiRp+rzk5mmFsc/JXId+SRv7Q2hlHkWjtpISq+ftqtMy5N+EHnNnK6BdNHIUGFy9p3v+YgWZ7C
S5wJQyQ0s/6X1KzXIDK1zYL/B/5zTbNlUE0YsbNJfD9nfrElokCunfD7susXtdnqwcupNWz+m4Xv
Hw1Che+zUCjaTc6c8SwgMIdXZdlWg+objeYq/H6IS1VnZsHcgqa55F9mxpsq1vkoDeHV36/qH2Y+
1Nma6juF7iJH3Txn7zzgmeNwPHz1vL+oq5THc35cmGYWAcWUhVxEseyXMlQEih73RubOqQo0tsXy
8pYPa/gw2tZ04nDDXim8whMVGyFjQ+JdZmd5nv1vDzm+SwppzFYXUcc/YjPncnnR972GBQcRtBYd
gQ2GgdzvTK+HWY2Ox5EpgN5oypsOWn/xQ8tSTgPBk1eRfRBGcWUBGibjhyyL+rjxa96pBkc8HiZ3
kP33zNQYLngVc9nRUfCx8rijV/C/1lvSagSYUWVQyH33vdd2TaqME+LZRFlJdaUC9MwQ+Lnyigp/
9kaY1ZWqEKNu9qKH9c9NzmN4Kyi8DkhUqHgxzQd+0rf2HMno/b+X7W6dokIYPIZbJQVDt0bTq5bU
z6SvL0FYLN+DPVdr0mTkkgSYEVfkyhxvAUdxb73vtnu/2EwiTX0gTsZxgmqz3gAxFSRXi05Xaacf
uOUGTbHeuf0/jlpqrgeuTY2Y5rD9AE7SiBi81yjfoD61cW8eeNdXLbk5J7fa2yHvuzPdkOt5dLgX
Lizl/Eo2BcaWc3SHuOEC7azoHkvRWgOwoTNRi+cwcq3Jpf+qdVWHFWKH08hu8ZG8yida1mgJlQFd
7FMw2rVbeSBDClN4u+rjUoICb0kbY8QCBpk1FliVvsSWSzO+ashZX+gbWQVNIQvW4lbEZXVnVben
TUDTEkgbMIAiiJW06sTCGNfOQonpYYSQAAqagvQZgXXC+Jf1/Bpo7JEZmlhH07UOL4TPcjB74ofL
BRhKAyM22zQ6225VCOYAiNeMHKdtCa5iN6W1c2WIF1waiRKzXcwDlXAbwNdamRFsYzWfNiGRtmEs
mQVkFEIYImv3x8O8QqS1rEH5b8EppYH9LaLsCJc15zDVFTKu9pRl3a1fIl9I/zAd7kNWdl0TJnme
1tPNnCpC7bniWEO5mcWocpW2H4ku97O7hfJ/yNvpTyrA8C2tBdmjPJ/p6osIaKHISviOiugKnvb3
zwOu0KSPbYnhIlDBCyz5Cp0shIo0NFdj3h3mWNefWNa5TfjYGVRQPayvbiFs325OqPPBqJ6onooB
Ow1sGB1jt4LfraO3YEhDVxSvUto1htsLmJBEfsEGR5ygkysyHbqb9rbNTTQWsEeX6VP4HPi4cqSh
eJxX4NNVy+3Fmra7tBOk61pwyIkuwoER0UcdROpZKtsz+4VdVB9p0HJYWj24L9T/onwFOl5aOpy0
r+B197lZRuY9bYLC8dvDfOGBDnXyoddNCOEKoviQqTgclPelk85QbdV7iUUuBrkHHbXGpE6jClwx
dEjlwbOPbjYBeBGzHAnQNDG2lDjqFMkD/lgUSCbNysALb/VsN0C+5n3xVCpEGGof+wyn3UQkia28
wtuHsG2likRJPOhemlYkFkMrtU7mVJuhgsoO+VBiDb8yOv1bLm2qEDPH/lG5Gq6r4dxWi34rBxh0
UC5+HZ5D4k3/Apo64lSIn6R3UhSbfZ4Pm6VU1q+CX+TTFFN4kHAp/AeMM5S9MG0GH/J/RCZqSkI3
BG9eGwRhGuITy888f9BURUo81fjP9S1LkFjU3k31fp9UO0DLgX0Aa3s8n2iAYP5fxt6gyJ+gnTSn
a0koZuskGwcq6Buya7K4ZM01kyG+DeQ5SH223y7gHiMAqdwljxLCvwAAKhn8qRZjBeqh2B/vwm/n
b67mlo4tK50LDtAydwTMbFS02A28c1DkkdIsn4JUfG4VrEdKnjMbk7++TCI+/OFMXVdSljfjg7Gf
38BdscFHKW2oGuELHbo0HtfcuTJiVpkvWruP5Kvpext4s3zMgTlNQAH5JrUDIukTskYPNHKccOrg
SKO+bXlXOEJ6aatWRUmtgN+TASdHrlkSouxV2fHdUtgYetJrFsHEnm8b2EDOXgjpvvtLOwcvuUzP
Jfm5gLypcukHycm0LT6o+Mrl4wuYdvIe2v4WYFfJCDOyyh1NCwiTqquNlgVw1CC+yUD3DHFeoq1B
mgUyJx9GnTlRoTBcqzKTudKr5ibfCE6HBGHVNJX/NxAnoHBYBZAxOGN6wGCMxwZ/hHMq8hsatVDO
1Pl+YKdFiS2aIn48fHlp7fTmYo5rP6qajCBPEvtkvsOLcxvFbu0i0Q4aaFQ3iCSbhZ/le7evDfJx
+aPCieWJLxf/HOVe2uCyq8+GpzB3rlADiqsbYiGQNMURMTs31PKlI8vvCsf7rxszDKR2YxmAgOWs
pAi9vmch0h1Jw90TZnTZ8FucQUsoA40NZShHi/grVRrizJ7NIvjBn9kM5NjNC4M/x5+yuAvO+j6U
x8dw0j4GHbKMg3ca6klKQom2ybTEnnE9fRIzKNcoUozBs5ieVAlkxKIZGJoyjzVCUi/FZ6T8YpRg
aZq1iTLBQ/IxlYSPysFVbW+baJb/7EXyuRYyQBTlqUzUgt8hb29kb6YW7BQF7QVoS3/e4vXEOtSz
aPDX36I/pkXi3XDgfRqsgFIG1gamIuoW87zDeqdNDRr+36F68Q4i+zV4m/sJRzQ5BOqG2ajglCTJ
DYuUA1XO+JkezDRR0GNS5t2DKe/J6uc8+lODj5tgmp+xCfKBCSSK4cURJb5Abw8ifMgVnOSUuUVB
YVnTei9fozEEjq0+RWsV8YnLgDoRqTJSStKeQN5+X8RPQwTvcnD1Q5epMZraEHhksOPoDtqPLO6w
kJBG5bQpKrLALPvSH4VGAUryBFHrsX0PrPhxdw8rh77/4kta2HnDu4l+Mm48bvgnDitrIjVJFcV3
KPf2W5wFRakABjCeQfSlneRj5A0rQ7e1bGw37kNgU8Bwyb53T5Gi/nkj043X21I1w/oOTL9hug7H
tnVsq78qd/Dn2kBdvxjsqT9OJFFhW4ad6hPqrenbIiscTouqKuIicxSkviP3ECyERO7LBSWeVh3T
XNiXIhcIZ1MCIgPkd5b6KOnpyaJBO4b+68lri6th8ImxKmS4DaeFeiypIj+liYkqNBD+SL75+9z0
slxRkBDudDfx8uq0d93VEwbPRWhycHr8qtTHL6kxIBaiIwDI++J1MNhckzzQPIGuoGGuXwdsk4c9
NNUSK9db7TLi3f8bThU9F+hYaB0HHXRcKrn3/xkBTDvOG8q1S56jpXa4v/LI6sgMNVpWTUQfX8X4
Pj9GmDt8tfYxWsT57SLUsBh0wabXcvgCm9h+4QLFGKqc1NajVMIul/mHyoENA8I8x2ZYI6NqnN69
SM01XP8sy6qZSBCfBYhXsTzUUmiuGjQYgJZm2nuAm0o4YWdQx39rtAcWAKGI4mTko7Wmw9a/lbQB
CMsnxE2qG3T5c8o8XZttqON6t3q5Qz12usYhpluM7rSvRYzJomub5aY/CNxkn0GoytKApMX1Ic3e
ja/Sm7c2R60jcg8BN9P1WhZNXmXsADHKuRcdu1KJvyL7++2VbGuAYQnrAGH6Vx0TFYVxYGX7nn2l
Bb31lpCGCciBd58yB1F2x+xZuBn1FDqx0eVA0dcsOQfJt6XsrF9vq5W0el3jcHwEwiDEGDhIvZ0j
TzB/0LoMJ8im7V+mxKjxTRgLMRk0ogrxZGMgIRy+sBy6uTUbq0XV5KhiizAGBsXm4bY4WGiqtaqT
xi2DOltS7Pzb7Alj8CwouY4YazQpuQdOM9OhBpa2R7TQfvZ5AqKI0P57yWW5p/WgVgA/yhNWxns9
9FdeUHfxvGqHEJKojnjM8WnSMdS0QM8naF19xbSWsLG1Uf32pGje7sM+2bQzGjZ4pbMkseYaExnt
uK67Z8d9x75AQbPohkz6h/uHS0Fo4ETI7nJvLh1YQub/hKR9iSmjL3zwnENH0KCq0Wgw/hXhPPf4
dcsN75a0DN6KGRD1JtGqXwPaHndIV3GXRhk2rloTMT1ITtcEq4ce8vf7iam3WJ5FgwoZwE0m4kCW
M/t2F1pLGCh6DvxRYZM0qb+c0ah/Sjr7LDfc4xSMX92vxRqvqJXHyW6fNuHV6y9osjTPYKZk7KSH
vvvUlvKQ3XlEV2ig0SzYcxM9RywrJYASrfZLW6N0qwsNhQkjnspXbW6eK7Abhae0j75JZP4q6w4O
EEvL4gFqVDALm+Q5Yu22kO/naPlzx4wU1rhLdagffDB9tTL+XGSkjNnlBQDoihCZ1TuBfyAyHDXc
/e4IbStwpNMIjs7rA6eypRAPkETgOCRn8Xopz9qStAEm4w8LAotZ8j+2wKIFaqaRqd8bhe+XoDTj
lroZmyxOCy9tEdXMowIL3RAOzkYmR/oHk3LKrV2bvyXw71NycZNY4JoYWirzETvi1ILYqpUs4qzh
+MRlCNr+SPC9nTovqFQt1c0V+4KxQsCm0AEUQPuo+L4ZdY0OvdxRe+Yj7gf2weB+sZrUJlgc8+4m
i8cWHd+ZLVIIj5dyw2CowlGadjUVICxi3MAuBdkARw1P9cybGoIt1p5AcGbcVlnDMnF5NIFrO8An
U4aSh0IHJQ3GtJF4Dp7ff0rc8WWQxIUXV4KhP4P1s6eFRoKUSFVJHqxItrNHCgZamkA4z7rCsE+v
tNYjwn6J4ZlWu0UEL2j63hNPVG7fwCgMejxydgNXY/FhoJxZLYJALe5SfheweCVjWkcmaXNPmolz
znbuQO1CrSpSzh5bUr6i74pHJt8gxt5GkQ02NcqamkfLQ0FzCLG4bBpEjiT4KBshGAjM8WpDHRHp
S79zhyelII4Ten5I4XqosvwoBrYlvh/IGIMnHe/54Jj0/KMNQjzF/K+pnzT2KPxiMd7kvCtCbU6I
icwCe8QE6BHw56E98i+nE1Z14ppsNuRZVKR3CR2qhn9vMSon6k28ym6mOf1el21WzrcFErmJ/qHb
bao8SPvlQ87Oyh7w3lh8SmabL0ZIoeBVt6M0JeXCSnaYNQdokAi7Afc+6MtOSQPjfRrU5fOTPxXW
2MiUlD4Yqh8U8ur7aw56qKtpQ6suWKlQnFC2DnYjV4cmmv8l3SbqwZgzsneqsZPiVexWJlevx22W
PKGk++xT3h/7QN3It4xhGCbdokqiB/vDpgbksmZmct6Fol6DLZG2lPYZ6kw1OCgSHxKBgUYFA/VN
vYpUudHqIz6YSgQpR30SSaCHWpRMa3E5YT746S16YQJl6d9Kkjov+O54zHveNfMV2K7n2MF7hN8x
AQiOONlRb2WWMHprrKfBrrF2UzSYKxmadrxwa57eDXJJiex7iUV65Lg/rITbzS2hWj6nwcc2ArMx
eYmQJbN8OdCd4ZxcoEZr3fsIX0Coa96It8S9MOFIJRHPR2EpXf6XkixckQyHOXIdIcWjZURdOmrI
XMp9D4wEAaNZ67b9uh6A+DwjfBDHVzJVe+unW9qlvYXOfgCDoLta1NpHyGnjxwTGritKCm9eU1Z7
z62vgTc/JH6EwrJYlMQDAhe7hCcnPVwkW1uJDT68awHe+yZ1I+95LM9VRbXFpYgnSrjXHkIre925
vKRQ/GPJOv7lM+YQTo36EQGg079OpLkIQRoZ2Bl0yIcaBL9MN1wJ0p6N//+k8FgxrxLgBilO/IGI
etsIjBwKl5xShF4saXH5ShHT2BgO+OvcU46iU6x4eD+hF3prJcrytPpwllMa0mWLG1i5er1N0gEX
eUVlQUAPInSwmMchsYC7p8kSZK/CtHgG5KOHprzoODebw2vrpbdU1nNRz9diOGZ76S2Gf4/vGG5S
9To3igXR3GrM6PVz6+9Z6gHrzaOUfaDwrFShiE7nhO13j+TNkFPhDZqAmtTDtHFyvosxjXNzcm7S
k217sAOfeLtx6VCbvZEjj8WjZkBMWK7nDiibgibiI/LAW5dRIlK2sIXiIt90jFUPT74isus0vrs6
33Hs+wam0+hXtgoKrvu8pUiUecwVNLZ0iLCUQHN26VBFLGXerg4rolVvL1aAI1Uy2LO3QRaH3E97
JdrmHpME8xoxxskXALpyA7lboUF/H7pEM51M37bsRMRv2IYrLudHEttTNJ50g5VduwGTRhPhA6ft
f2ezXd4dSngvSeYDkxLSO2P16ObR8zGadp2XYYYqWboL/lZc82+v3mdQJXqA0WCI0YobebBVRukG
NcMXNU1ktyqnWCGKcq3vCekCF7wJ3Mc9w1TjRHcJ6Tr+Dt35IIBijIZIvOMk2sxwfw/udNUZQyIv
QpzReMMkXl3vRn2MA9/MhLliEXaetTH0AR7CGzf+ZLjDpeO6EMJ1wL8wWy3adQvdMeF0WqYkqu8i
14pohpBnFH/W2M2m7y8DVQiCsMVKtl746sP36q+anYXJ2wP5sv3eVl8g8DEWgty8mm9A+qiDosXZ
Ds40pCL4l99MOHCIvOA9JoL9+N50GWBdI/3xgvQhG6MG+9GJgYhx8e1klyqUb3+2gXQIs6szXFg/
+k5U1r8z9qq5BEaL/aK2a3WZEAJVIJySM4vEfTD5ntcF7npAghHyKzG5j71b6StRDW81McUG21sL
OXj9zlYNr7ymtjEfHS+VZdGRYSVIDnDmVTEoI/vTJJyksLkaiQywrt/3l/bp7j/IQjoWUzZFzj0w
fb8kZAZsYC+8HTJLRBoqF4yJqAdV9NNkqmo6udZKYDBDMs12RPE8Tf8crcMX/ULswKWPY4ttkh6S
orSZ8TbgjkzLqkDYDzUvtOc/ZMjrqnqfz3ckFU30c0VrMwLOqVkv3XSMJ0KCaCln3pID80wlCy/n
2hMImXAJZ3RNJu9Pp732U5FXIz6PdNSbnT+18XV96VoSM5yP2DK0D2C+e2oB91ULPFbUcI+f3dAO
mE5+gZ/n1jQAf6P60B0rrZrxXGCZhlMvzqgNxE5S6w0i0FPz6JNnxWEaTOZhqlyYcKUPr4NdVI8/
7bLxsRGFqiqzgZlC87JIBqtJroqI/sbDN5s8D+2ee6RLTiqGPfVUTpnvZ6SIUA7UpG/ulRr3qEA3
pxLL1rp8+W79U+zvNcbbNMm820b0ht0o7O3kiUcvbLJDMsjSz4RmXCAbdpab/Q5UThlx5cPs2Kjm
Qqr+9jyzLv+ZV7a81kYjpqieSTh+XsjRzX+N/uACNokAj0MjKG7dywiSSXHYouyi0AtSLS5YMH4q
Ej8K+XtUfNZ+PG3s9w03nbJBFrG+tz8nqbRgXsd/ZHawXe8WE8pUlVvFxGnkBu64CjYe1QMSRUoA
mmMwslV8/dq1LypzqsNn9y/Zhz+L2tUfaT27vkNt31yO++VKaCO6kY6SwHfAN78XXyVBp3zAVuNp
ZASMigY2xPpOYCUm9/Rkwe/BbawxJWs9rLGF3FQUznsRyT6n3a1jYqYBbpo16B1Sl2TChYTfSCD8
9YU4iQ9ilF/kF95z9GCLD5NBzFEwSiW+CcloK9vo+we9hjwEXu+Nxznp12DohUQMwpcZZfkImSxb
uJO+iqhcaMdTdqneCTx0ojtA8Kl3kCzB1iVJFnL6g4DkhNm/YUgQ6S5VHpNfb4FUG2VjZfrvtMDm
2yE0h7ttxwIPYHh3GHqwtDjAcX+uHKaO2eCE3ysFC8Eu5iPTrOi9406iuH+DWj0J/29zbZwFIrf9
AaFIbCa2s3NN/OjFAFd7gTDesKSKCnkCvn0IQIeMf/z596LMWnFhfu7FsPppbjf6UCOnmrx6SvhP
QDMESf5kYCEZciK6ucNbNvWM1+/jGQ5RMVUrjW2yFfNUItnuBt7/TMVUTjttR35d+ubp6kQKs/oU
Ed+8xHkd/eJyHfqvPDAdHTMSfyh9IPeskIYhBESud43bwXp9ADtA/mDzanuPOyXA4nTAEdMLYOyv
XxyI4p6RgKDS77ibrkH9S88NwpsBEgZI10ghVbw8q48DIlc3qvWnucTufB4sBWrPzabFefYxyNyt
yqetTIwP79NsnlpV3xzVoBA9go64xUz38jGXVeWXmbCDeOoL37YLH84MV85iZ+Gj2239Ad2n7ANB
r/8rNMP2rvwOSlho4dDfIdfKjzE6kVUH/9JXIajn+1zKLvMuh8eYmWcRTGWZhWnDQC45b9DB6yf3
CEiox6TrQMibFDoogZYFuEB7L6Y+mc9+Lm/K98dU54HNDfuUO7sO4sUbE+4cy1Y0kigGDZZHZGcw
pBLGOcKUmleDglcPZgzRJ0kBF06yHziDJOke0xMZ1G79ETTGk7+SqIrVAeaoZVyeKCzp6vTrdRf0
rW9/iOy2BPjf2JrJAisyAappBAJg35Sujg04x0PMCNqsm0YXsj6L+AsB57Yw2sGpPMdQL4p03VbL
UKXEdocurT+DCd5Q0wm9/9CMoeMFxGuP1Vbe2DZ4fGO8Yozy7iqfX8gHv5j2wF+ZFwt85Gfu8sM2
46tgSx4ZWPwmuCm+wcpbC2JpkT+TvLGxV0wOCL/bdzhwudW1vH1P2UYD/YjaZmmCTe/E5xfpcmB2
YjklDGKsOBhsLkxUOgvJWjG1wyqPyBd6NZd4yauNx8gPivq0XJBKGo4PUrxAPN4N+GFgy5+3u5xp
Xp77HrWGIGuPo19qrP0mhO0h3P3bzSrZNtsLNMcsuu2ETgNlJa2EpUMwciB2mAiR2Yy5r5yYPI0s
6pyfh+R7AFiyveQkeCKqr62vMI1+/NRxM19OLoB32lT1Mdv9eVHGr1LrlFcnLgXGowwXPOGHhKk2
TTrfqptZ890YysGCo324vSDp0+sy3q6BozqWhb71C+jbp7oPMfL4uPUBDdyKBjh81LWTw6Yt6mVj
4VjZPnpwTcQB943kTQmL6Um6mos+Q6wn/ygHX0BvtRLIwCRN/RS+UmlFzf9uqZGpRT+epvJVN4kt
NjYZOsfzUQYJ6vUpCmQW+R7eiIOZS98GnLZi51f1YVnWEYgpOgWUUu3fTqoIAbWTVd1wCrxS6w4s
C6+eRnHnT90YNq3WBl1+xy8KEI2IHAfhvxIN+R3gczOxoZ6bzy0a3tJYe2X+uWyZhOoJgrLILbnz
Ody1ocHCeetWFgKGJzrgsTCtvyfSSiVQTLqyOhHRSglHhwOoXv//QQCz91Hn6p7Urs/hS6CEiYEB
7RhheuxUPYeUGt0WvAPhvgzbD4vH5u80g0x5pJ4cDRpFX8mGaPsDcW81y+3cBfQ+L1FkIpT3qET1
n9T2TxRhckro2JgDekyGeLbsAMpux625OEnSGJY0xPSgiyXdSZU8gzHcupqZhtV1YW3tLjD2GEJX
qwdvHl0jpJwyd1jHLsCj9+RB/DDfevhHboItKlwN0mELBTT9cdScXN16MMGMf44vxDLtKN6XMlA8
YMl9fIQRai79fdtHPzdbIX3qhXxsn503f7S7drXoCRjulxltwJJYFGIfPrFXA10eJ2wCYxdMnjAY
AwQ3KcVxG6//HL1G2+q2MgWu1d+LbH6fi0NT0NlJ9CcEV633WmiYpluzmn4AMM4BdGOn2g5RzsfU
SVOgBc5RnLfHtqD1WXe1RBNrmhSPyCNXfOCiGDhV8WEZEiJbUUViKyJx3odal8TxInkcOjKeBW9B
9H5hdVZpWNFl88f6xC0IwgJr4DVXkEv7olF2or1xfmq18JNkoC3gd9di/ZC/jIp63K/WX1PwEC6C
0N0USiup6c81WygmpE9P8T52NVwqBZoxl2Dbc1ZxmDqG8meR8PX5Jg13Fp4cx9idwLl9Idz+YWrt
rvoi/NPb/IVr97cfhR/+nQjju3V++YqtkQ8/NFpHBYAQrGUgCzI/NTIzCW3bMpbqaLUy7NlZ7E9W
jI8GUqCpueSN5/tankT3lFD+1aQk2X7cy0vdf5/ZZ3SqJWSPpYu6bJATpHLYKdzzOmUebpCVaE6T
8+vfnB4dSg6ws9Qz7MQ/xs641iNO+alYyzE9sED5hbHSX6kzfBY/fzh4NStQYmSvcfAQrXDfizvG
/v3iCEodXxqxFHteSjzeJUkwvSoJBo5zaxuwssYf4Vl7BPeOHhta6augdCNslBJR1ya6eCEx7s5f
9Vctc05jgspOOVw55USDt77pyAGowJ7iQvoVPuwLZSvvdz8TuktiMfesuSJwccIfITHDekmUmE4O
D5bFLTr3aaQfioIPmwyGAdzRPGHvhGJamYe1dcvvzFWTdcLAfecQtIzF6cw1/nTNwzdEiQXKqzUH
Xv06MK5Sju70XIbsvkdfIO7FojL47/MehkC0vE0j8XGrKfBV5of120hWKLsJzrgv6m54hZeRk1Ja
NaSWQ84dB59GzgvKufS+ehhrCTya+JhYmCU32ZLF7wBplOYHjVFwk/V91/pZ95GZlBOZXyhdoOp9
D8Q58otZKgviIq941gbhXzbQd/EJmyBpIqmxGmOrHbyVlDXpJzmdtWyxWA7mNWaeJuQj/GjWn/Aj
IDCuS6GN6A6ySTWOSGkdpDZnNt6RNdfKFlDDUQmJtv9ZmhLr9K4CS8Bc5b7jUwvE6t+SW2XX7XLW
DyH4a3ygtgvTJTVPk9bTHNnDjlX7kqfzIbS0H/Cb7n9T1neQ7b4XRKogaKX0dl6rjdT+USKdobBn
1J+sOGgIF++Vg0gggZxCBtF7CcC3JZhQ3gUe88rFmVor5p/wyrS33Xa2+3rVwvi7q/kOdHp+Nihl
1zVOjBeBAOcD0H7aHkD5/9jeVzvQxuBF6HjkfBXPIdsEIbLFBi1xPPGFtntFKAzciaW+kGoc3f8X
uOVfcqmDU6nXKgTaZyhSX/LAqnsgCtRaDlNciAY0hqSOmSxsjWSAG6ikTUqA1ZWCIvoWAzYubItP
bAAYAt+CI4FGi9BvW15ZW6gXI50gJjgITz03JV46whHdUijQwC1UjlfjMOpiM3qWx3QLAv9BPtPI
lIixUpbb8X+wknAke1Gp3H2YiD6Gw3wTYczXprTB4ng2rxnfCCaQDnV+ExsM0zlSUuNb9A4Yc63k
pyfKEdvENezgywrDXWyhZKjttVhzIVX2hWqfUuXmUsDuXFdlqPmWbojUha6kVcIIs7eBioxTIruP
I5b+xubgu+QX2h+p2eiQaIXbZ3lHF3dhugjHUs/phyzX96+rxfSD+n0YglZnCsXUJe89XHJxjfOd
etfPXUJEh+SZW59SLcSnUKMO8oFeYTCibV1s88ZTtjK0+i1sSJbey0NeL0lwchmNw94O5dAG+Wn7
bUjXtrsCBVdM9fT4Q7akNYo0BAtCC1U6+s1WeMrwrN0hj4Sb2gTmjeM2SiEZ3gw4/LxfFhyvGWJ/
/QhJ1TpRAM5HDx7HAqTJ8DRX8TUB/w/qjOixv6H4ZUo/KovO+De9nZaNyP4cOf5t5JeXAI71xro1
+Mrp0QSlrfmmwfxWI3yCdF/tPKV2xRjkd0B8vCHlEH6BIz6aps0Y9k+xlXaK0QfJZV6AehE5Oddx
66ck/XGuOhqJ8n1N699XUvJy0xLNoqfwO8zS0kQiAUL/pklqzVvIgU49J4yebp5FqwZMzprjhups
031kd4LS3x5t0l2E2+bDGdFSqRP9xQ8YSg2+KqiKj6bkgbXqc2YeQez+1UjeXo9n9RSrgXAOwDtA
dKG0tKxAmm6WoxbEkeDq1O6LzyKl2OAk2ybtBG36qeAz8E+jrw0y/9VxJX7VGlFwmzjBL3zO0eRR
Ix5htRxm549Kn7N7CymHWeOWYK0aVr6xQSEyqkS0AJ5rv2w+beOrpBfthiQd64LgdXX/mV+k6nX2
hIHUm6RMTCFHPLlm8qKGnXhsqIsTxXAyBpM89Ru3R3HzWXPyTND497tatoX/tmDCE+wHv36b6QjE
zj7EKofpIV577e7xBDL4Iwlp4FYIy8FApdaQxmoIxlWeQvTdmN6HCmSZNyschLLGQhhKsW9LCHO+
Q0DkLt4To1CgNHolqNwL95TFxJ3YEKS/N/gWk5MxcIyJWSvyoZtfUq7QrCz43i+mQtxzZLZUbWF4
HFOGf/6anCwJ0OBVCBsuVsNvqeJJj2u3nMXnkF5CY5OCH62zmjyq5jtjp3Y4qLvr9aBqAQt/u6BU
JKRoWtweCx8iJbMJUE7g+ZxAcsehhwdhM4xRzfasEnyZ+Nwo34D5ELLdwo91h34OJ1iwDESlxKxj
pE5OfFzHc+AAUuNos5mBfCnkmF3AEbpj/FMOZgc5sJsftZxLWZovYHGvSJK4x9MghQ8haclNQAgC
vg65ofAyWZLDFFqngC1QdpokKkCVnEP7UiX8G79dg2kgQrPqZ9qCljbo2HzzVGNnYJwr99d/Cvdb
AvLHLk9lzO51ypUqM+SB64KzjULZ08OOQTBemsEDqJMytLUE0qzBpqVEnFo7tNrwI7+VS/4nsfxu
vMlfH/iTSkaDDM5DeOep8awRThfjCkKxsENuDovDYfzcZ+NBHTkeDArpGhVIgti2AEMyYHIwLkcc
2+YZX4GXS7QtYFKLRiEHLRCdzbZd9DaeQsmMqefsGX0bgyEXAWLsjWcxK+9Z9U96tl+7m+Tf6C/K
PEiIC8LSzZiKWQKnpCz6EHvUMZfu4XuGJ6ARtiVmpVD23XV/ILazVowIRVP7co/jS+jNE9s835VT
HBa4CNAawkEcTqxa/82FOc557jyBqFIlG3xM3kAqm5Z9PnZMvl0jkNclZzGKwASVqhGLrv/1I1xz
L37JaMN/9CB85vEbR9jigWkQlp9wWmuUqCg9hE+m4ojYKYZTi64CvAafIHChH5CY16lsRV9ydyP9
ZHLlm/kASl8jq8F8sM6E4MLjPEFKBR8mwI8zEr2gYEag1nImnLYrTDyn0Evm9m5aS8cxU3ax/snC
RYWiOfp2/Sw13RFGDOOLl1oyIaowsOSWuNvBOqSXfQBBtcgeu1Gw7H1fe4Wyu3anEJ4OuZLGYscO
F2hjE8zFTqY9yHLG1FlM5FEPYJrPBV289GOif/RlUuiKJE6qZI2cG1ezG72yxUc5VOwRiLoPXvij
dRLIb0fniMDqXauJ/J2dl2JBlex3j78rSRzkRHWniBrlyo/Tda2tu9rbJgEynvF1WPU76ItXk83G
a//32EDct/V+snQKMIeegiQkpk/dAkkMiG9uA4NDZFxv+uJ1C56FrdMJt/YbqtJww7pBngPEKTu/
5JVPKSyUY3XQLautjPI6AjaIO+I6Cr58ZS5NAKsiPU3463X3Ad7YYsdeN1F9IFB//i6zRlN6z92b
plZTwCwlFYTaDemVgeWHqY4vF/Zxxr7Yvoxjcg/FXYna6Dr4We34qdYditWdiS9vUcgqhe4KAy4y
tUA8vvZZfmxh0/8/opRYbFxT3d82YYKLeBOnZaNlo2tJTg9LToC11YCO3oMqUI4+2yc4JD9tvFu2
xuuPBqtkKuU2CbWao/1UeUaYOICEoRxL8azcbQ5XfZeVjnxbiEUuBCXPpI/3w73lVDoonlqPb9Ch
vxQ/pyIkl6KAjvQ8PGe+/XddoyjcVji+P3k3gNmoKrpQ+8HqpdR15gJyiqO8OvgJnMpxFmex6f3M
V1t13WCp9CIaWr9NgxsDz78e3Lfj7QEZ97rRvnKbpPIl6E3CGBj3iLdSMj2Dpj0sztAUQuDIL04D
wWhpd0p3EqmT3N3447C34C6hpEeTeiLUHcpNjHyQv15sod/419Yd6ooeJ1x8vdv0qwfk8NVtht5y
vuqZG8wn5qE4Z4pJlNC/RMfh4EMcE1z8q2lLl+uAr4NRAmYx1KSkXO4EGG7Yf7QfdDmARf3ovv9o
lDVJtHlHjrWXhEeXXDMcoUjNc9CbrPTldMZeM+uU7DpSTt+ZPTGyCwGaszD4yH7TlBtqmIAgon5O
vRAhvBBc1vapQOQJilV7Znyij+58IwRS0CXg6DFJYC9iRVo/SKG9jqBsEEzdfoaHDni1fpETFb5X
p/LbjZ1P4ntWBFCgtTK1kULZXDIvA9pmcmwkLbUyAbFmpXUD2eBD9NIa+JP+YakW2fBMqwFVAv9f
u/+3tYsz5qFPOB05JZE/i/LbaRmVpq0Pl6lGyXss86x5jd7INhme+78Ee2GoPBBnIDOWE6Sck9Fa
9ti1X4ikyLxh1+7Gy0+uVN4Ue/deLHeak+pbPTBm0xGWddJC7U6pOON3A0PKDxQowL6TSo2ipCdc
FHo9Y1dQKTWyGTIGbG0uA9sXXJASsQ6r3GZ42k6pOWPTG5vrV1YeB30iy3vL29i2RTWfUAiTimgg
qzn6iwfSwOLK2pK26mTFxskG1cPFCb5rN429NoWUuiRBhSSFUjqxaz10bAWEPLjw0zvE5YZOat9R
nONXTmbfUUoRTsqOdW2eJ8bNCPWnmixnSbQ2SMKbFEGAtLXUg695HWDIIsUIIKs3arI3YngloZ5M
ycytad2jaI7Hxz679QYzUfkPwd+pz710qZKfZsrwxkQRf5lnetknHGyUMOe2rQ4f7XluKcK8sjha
PsWujkboZ82VscS1UjjvuchWVqeMq/UWZ51MVnnkZppBh1L4WRvqZSE6mXGgpwhaYX7vsqhbmx5g
z0E+2eLXYtv7i3qOCnKEVbEplaY01uVdFOa91FSKS7Bw15FNHfokLOUpnZD9pMFEF2z6yTGL7y7U
rKEa1cyhqI4869WYQno+XS2IdMbbj69mHttECWL/3dGa9O4LmyRZrGd4eO7YKu5DXLn3Tkz6YkSh
l77MvY5G+oz9NsMi+FJ+Knq7HnML1W5wG3qrOjLg5UOJcgFp+8fKadrc0DlBiRLI9GLOMpHMbjNG
BQszh1Y29+9xmdTn8OWV6YSh6DwbN0u27MqSfsBQAepQmkoUANAh1pE6J+3/V+Dc5xl5ZGo5vTXW
npH4IeD+hakCWHyaECYYaDC9Mq9y/83DwTLT+3tXsl4mp1iwZCaTBe7K2hdoqRlHJ8jJfiLhV97V
QmUC/oAKh6uO1lpT08pSwlnZ6qKhuR0AklXwBdpRR8rmdvwrdLIrMIT9EZKtvU849jEMdKoJsyfm
Cb7hK6jk2O/TrbiiHmM23Wb5B0iUctdlgy4IrVaatS3hD2jEHYmyfUISHA8lCh9QwsCSVP5UT6qP
yyPhUXJ80Qcy3nDRCao1WphGf/w0Ud8SMPT8unDAClB59MNnUFg7gGxopdw3t5IbKetV10Gp2H1y
IglH/efHnOiHL6hew6MuJbUibDUT151hlKl4lvegVQmxTYID9PVxn8cwgFdk45mWXzcBbjm8E2DV
rG8o4Jr6ubZqZoiDQ+F9ZjPubu7vd4+Al88cMDwQ/nG5fLos919NUQGpZ4cpVKc8SgirzTM6G6By
uyuxDGz59MP7WvCqHhy6YnwdnlzBqI8JDfb2c4PByrNZue5Z0bAmJVhIw+AHptzt7m5jL4TCOLS2
KWm8B/sxZELjBIvxWqQa9Krcw7Ok17P6Zkw6QCHVb3szmU44sE5aV1bNB9Vb6pXhEBeKT9+PhzI5
6PVhdhEmYowKrX2/NOzuoX6sDsBEc8dqHcC1KLoJ8MZK5bRVeo4Ct0yRZ1gJVJrqG+UwFiJFfXmB
Era9laR8ETRMymAD0Q6t33JCU/8+ohOXqJa7B6UtLijdNv9ipEIB8DY7rhJ8L1sO4OUKaUpyI3NJ
OMBzv9SfPg8+WuVkVdKXOcNLhc5zdIvK02YDPSdwIM1hL4Fml0BZoa15x6doyCXOV7xk2HPKl24D
gDiAluHwzWuyClMWD32wUhUmpjlMeP6GoHRezM4zO53frFjkPlMVRTbtRzyKgFtMX80fKzhRCZAx
WVXvyeVq+dBCFQrmx2KDmbTwd86EzEE4Zir3JahFS86ip6fxVBYiaqHFHtepMcSBRr7qd2HkG83T
k1Sd6vHB0lwJWFVqmU+pmA9ngm/bnnVLbALBH8EiIraJspI2pqHdQ812MRIdMliBPB7dY5a2its1
PAnwBNDzzUJP1haEhkfKpsgDR4G4mIaOiXwj2kIwn3R8eJBTisH8fQiDrhqE1/wlwhKmqKMnrVOb
Ur96ga6hF5tVQX41QdwLWMTjUyhZMweThfo63ENru4GurNz/VzbrUTXXmqfGRtoPZfNGiur4uhFY
nEhBEHx2DXiNzExF72pZVliTuuLvYF3M4RctzAv/zP6Vw894J7AYgjIMyIMrll2qhxsTWvVx/E+y
wFhU1PBXxoW2Z6s2RiDVYK0ZzGXQt/AbflM4tODacm+xODsG3gAL5YakmFGAzsg4Un8kdixFqp5r
8+nvIvX5jttcZpdGPkFTHLtwQQW2HuYY3j2UY6f+0zHh7p+NxruB3isQRRWGbOGXu8wpzf0POybN
EZGAkVQ+hFfB9h1C+KU/vIGtDQcRhyBIn0HrCtF3yrOWDM8F4rC2r5G3qAOXbrnOJNYXtJ4g44vP
jDaS0M1PdwBGsPAMvqTIo2ZMyElvHzF4e28WxMu/5AO6ByrCDRgSKbx+BlXyNA4Wvu/yKKfCZlRg
nxtvuwCh131HCC7d5b70VvlwpgcgQpbxvH10V9ARBdgWf2Gt8+suXb6s4wLNj2tw8hgaYV7bST1I
L7ZRVnnYGAW2CLJDp5dyoXxZaxFV2SEIaSQ3OotBkNjiegg/oj8M6c6tGpOKTkKbx7ldrcrRKWYJ
xEwTgknHe8gNerH1QuGpRh45C3TfE1WkA0OOsokwZqZCpzFoiGj8K/UMu9nYzFQjoLbwLIp/vTqH
YREG07EXsgwBAxYkUY5NtevWGHELoQFKx2syUgUJbfkgt48mnrqgVtd44rlO2/uvj2gniKksr/Da
D6yTQuRYLrAyZEKnElKMrdZ5ejFfprCg41NEYnbLLLkaF2bMAZ3pLPERN0ZQN1n4NFX0c/m8+81V
Ta5PzRZzIMGezyRl9Z5qX0TnyqCansl8S6cxYP2WvTu6D+KkbkGh8wschHdLbMqKhaerCXBtPd+n
BVAf5xmmLuga0NLsPv8vO8noaRqC6fUaXb9DJLyksw4xUMM92xs8JLMGE4URPDM+ajQ872KXms93
EO/ThyICEVoBVu8gukxqczDaDThY6aKxTOhfOPhuk447Yd96M89M6zP122u1z/qpiDMz1vacy3T8
UN9cXuB1NWzv32PqSwpeR9q8BJq+nVUTYfl49U7Os3QZf3lWx4BrFrdBi/pAJLmL9h5hpumcySGk
/TX2hoKpzV+BkshACh2PmfsuB7LKlv3Zs5jCahuCcdfFlsHFXBA4YKd2qt6LxVRs2FpMdokU9ulB
Tky2+dAeR8/F0sbiijp04n/9LHkIgtNoRIA1mAVBEgtCM/UEzoZpeMfwXXUjQBdbdQPBiKr13eSD
ZSiuDx9YLhYA/n/7colxYL003QrChirsFaPJKCWy6OeMAngfMpDLW41nUIpEjH25qBacLB2L1zor
4nUCOnRi4lO6XeZBP/yA9KmGu37pkI1voiAD8Jk1beHDWoIauk2yRD9jrf+zNB33NgHBx5iUs1Y4
/Jdrqe8yaJN/ynyJOtbsMBx7+LmrKz1rMks2B2nbz+/ZthOaw4oIi5BVZmP26qod4Y0gEWGT1Vnm
h0pjJHzcUovJuXuBKRIZJ/UXlOI3sJmoxASkBECRPc//JF0QVeRgXALjKqr071ku+/Bh5SL6aPLh
Lqg/Kdh2fBfAf9zPaHO4o67THgyQdYF4t7m7xoYNu89/M/aLZWVsGOcdRAqsk9eKmlNUoV5EY/j5
LnW4Fa+Zaav4ApmTkUc2tDsncFcebShBvpHLLkQ6retP9mSj8UleF69U8QTfMeR1R2dQlEzV1MOB
C/ZXSafHXhyM09gOZcJb6gQWLq7KD/2K6t7UrvB55VwBWM7SBEGtJonPCTYWwaz0mOb6uC3YLd6V
GXGlYSy0cSL1n41YDvsEP+DhfGFt7euOazIqXl0/P9SFDgVkehVddEzrA0wDityt0VGjUrCsr3k0
aXat0BO147/0N82/W6RZMsk3hRy0ItZE7CSaWrmMFxE0fgFmWfAccleOiLLEuACyGxfnnMDCovD9
bx2+U8BsifYgjrpRslGL9ixO1P2eWeaUYIfy/HdnxDkVP9qrPptXhRa42DP533apsDs206XGXeMd
mA6LtUz0pCyK7NFxUcRLheos/y70+hg71UQIODfa+zyhM8xkaFU5BSRbCEdom+jP5fAN8pP4fM3R
uJX9+5xPJ6CiHctgMFbWQdV1z1KUJv51yo6y4/ee/7I2AVA6Ek9XiLpgGiaXVkc0cu7tKH12D5n+
A1GFhEpIWy7f9R1XEGciB6nin3vucLWIwap/C75fwufJi/s5hB7O8mJkPm3zMpkiDwhsvpnxWbDU
3sfvFJilFLAX8zqUy8v71EG3hicbo0NOBuTzDp6NFNknRc9mHpZNpDz108mTFsMMDLZ3JamVh8br
oiBSD5BoYXHTw6vU+7GYXvhtv/xBUrcLV6ptiApAElMv2uWh+Fi+AhDMV0oARSlhAZGCDuBgD25p
ovQNwK0mFFzNGFduCnOnYliuFPy9FzqaORLCF/LpF+ZJdyXUDMfBCLNJzQHZONvJucnaLEacb2Uh
QqiRw7C6/kFPBl7+n9VWWwbcnNTa3WMfcb6eBVqph0G4gLqLO27RFLEt5DUQU4ymjpY3BC1IhGL1
RW6VktVbJwz7K/i8oxLNVm/Fwj8/Uv9Sm5YwTXybYOJ22pZMKs0/EOWnTo6gZKXAhSXTWvEw0rfx
IFWSDDZgAn/sV7L1aZQVGO2npHWd9j8awtyGMcdBkBHPkp5cgbSWeee27b6kM4Z9TT37dbLTymQV
ygcfuJF5sdMP766XBG093QA6jUf13DofckdhDkFXR73hI2+9oiFgaTijK5agtR+4MN0BnjJ45fTB
+xiVrWrJVV4U3AjCHYXbzX+1cMajvRh0q10f9Ar1PLsEdmC2WDK8WJlTGDLqhADcIknXjU9PJcCW
WYp9YsUcic5QkhizJ+qDU0aAnoGiDNc0YVWLej96KLVeVCd+2xVp0huUA3cxn0xWLIjBY8TP4QoO
UcKRwrhhA7DIFSdFxQZDsSTMR0XmtBawbbZgOo6TjSVQk5yrfnfhE0ZZmyJK2KILFVUib9j0NeSU
pw1YBqTLkC2bp4vd7i19tuK0+tp7YAoYiyAlq2QDxW7ny5uZoTOHqLAgRC4rvww1nl0knJL096u/
q3Y576EjVPI6Mu8sD8eqEgOz+80RWubMAgl9mavFaCyg2zTgbqaCU0Da5zIydVGPEiKPRhHSK2Dh
Zsb8Le0aFBhHQXuL5d43xCBX1mUhBsnf/Ad2ANwYDqMx0mtvaoXq2LR12YPirDa2z1aiFDOSazhg
U2WJDsBAlO+huJr+NpMZTknZUdMMNGbPZqTEV2cR5I3c49tiX4T0QFHw/iaAnXUDgMW79c1o5m0m
rL9TsGkGxLr56tI7fDrltyOaPQot9/AbpY8MSBSo2BZHi1fV7/h+XNio8QTiOkFATPsKeA9HGeeb
D1ahsNRHmIPVTz3yqT0rUi31VAT1/TZG3D3FT6JrvFzWqG9dig7wpP0ihhNEr5A3qHftjfClXcLh
c5jNIzzjI3STwLa2+VbQdyDUG+VpmU4zcuR2S+mZ2zobj/3FJK8Y3PSz8y7UGpX6Smq82AM1ebDv
0xT0QrdWTMkQD9Y+mitmcz26gm1Bv8N+SxfovJnMm8NhhpKkRH3hDCZ2CiRvrp0D2aFdOKDJI/G7
RrdYQIN2j2dSWq6ANo+6R66j32gOHJpbf1KnNrvGqHtVdCvZAs/EueIB+vTWhvs3TzJcQpenoHLf
mZdWZafV8wFmyvbDnzS9XUBt8dnBPMuQcFA6rWXXau7x4AiK3bXqlmkz9ClyO+3whjp1Ht6sDb9o
MgG9AolhcOzmNYzA9UVkmoQCrJJloxl2BFIGwI+tSrC2w0ZSuwE90H2F5fNP3ajuzcJjxAI28xTx
cfPmwdTcydu4YvrJpRODM45815j02fgPrK2VzN0De+4enfWqMb9fvC7IdMOPRCtmynEpxrIU55ip
1ojXv5JfQb1DwmtqmNhos9jSSIoATA4DO3LtJF7FSkJDSxF/ub28y4tkE0NK3GwcapKLP89UkIv9
AoOChnNvQDADjGBRQjjw7hO8J2huZnfgVer7cze07OHokTrL2Bu/IWsqljayobXP9wIlxkzcK5DD
MOlrG7f82Th0AZHm8feBlIGIxPFRsK9+qyxRAq/Waq0T8iTphdYi9SQtxqZFOdO3smtuKgsivHyJ
OMEcilKXg0jEYnpBPAG981P+Ctelc8mdl/Kr01vtWrnQGEKoUvqSBhSvIkbI+DR5/zLn/YoZYkjj
Osbkve80dJxeWPxFiy2lEcre1ioQo96sXUD41Mn8zKpZXBo2mooJFJ/Ur4Rd38R601ddBf4HeWob
dREAyBcWIWKrsfyntnsnYtBuTo2fjfCEQOj3vxbpIe6KfGqzJFo0iHxvc7Ix8uwix7wyqwVj1MIG
c74lf9/VJJRe6M/D2fziLwkzUwE/qUBH8s6mKHkUuO1hEGJBnoNXV8z/OhyZS+MIFNgFoZZQOXwf
TXf8do2huTuS5frqKXDbFt1CUtJI14iGE42vm1RIFAE8a1xoEx6GZDCq6LIMlbLHmnZ+XqD3mMfT
8q2zLt4kM1Pu6nQW16S4o+lMSuxSgdFecgPe/TJEibp7ywpxWsxW8VraQ9hv7QEg4zaUS9a/Drx/
Zaz9ybb+shVQpwUinDnZjegsnd+jmrXENplzsPAouM6+HfEFix+v6YrGx9krxV5q0nNUxMcTTpOl
U4L49vyig2Nk8lOLYgpLD4OjZXQeXWbRLT8Ce++BmTNyMFd545L7DEF4heE1hE9caVO2/Bmxhl7H
VOUMpp2/7ssj/2RDVT+bMBAHuVmY995LCYHbSHP6W4lxA5mxz3YCeVFV0bMOO5XeCyjUVbepOEmm
CsUJQiBUtlIewWab4fYHO2ZSpEWY4HXXwgeJ2vX5uFzsMbEOevpadO3NWs8gMbVsKvP9P9gYG930
COcEccQShgMj9qHTgHD4L00nhe4wkKcFmii8rgJMeuWpP+nWWTikrY8Jsn9AZE6RXOyAY+DlpGgn
vDYXUSijgdEpSn64nIG0Z1vQ5WD7IgbdgJJ3B34sIFCYuBaJP7RSj5Ak7aMS2BP6VG/WSia8MDif
Gslfj3xLTt3gK5UCbixrwmMSPtSQ1BREF9JrvhVguJOGNe5Ql8Pe1Jf/SJJOSM3d3sUhrdh2onjQ
DD91JV2JkzUBtF3CVhfehfNhGK6RNWnEDOelSNdoiZ5deIk/DB2NTJFxaACXgZM5Dvlul/Hr4DbY
ngh5BBuxBrLQRlRlvO/CLeXk+qi4XWoqyKZCJpCIahtzufb1IxE6AAdTaGUHfbUSDKIzvSlW8sWD
tLsLSRotGkOcSMKDkWXZPXEpiYK4LwqypUnzpSFMvEIkyKP43F8MML1HIgSynFV8Lilv/dW/8fGo
xOvUEEg6F8EggySUMaT/Sb+PRdgGOKSbPkYanJzxPZjvHcZ7vhemDdkEUHQsp9+QFSt7Pq18n0Ba
LrcmMhLUb3CWMntZ3fJXbtoaOcN9D9NC3L2Avzr4vtMKHIRY7WKMH00mbold4RBTJ5NUY2GWM1iu
TylXj349FOqBnqLQdMbuMn1JxvlcvRHwC84LOdY9cuNYclc5dXR1XtgRbA4wo4xHtmOwu/8fsDU9
qa3CODSrOpODkvGvkpRFfkaEp8EF0ABG135NvVvU4frTlxUoCjeDqBozHmxImQYgQXDgrHFLEvrl
4od2VwKpehXyleglLZLelRIla8wVM2MLUAnrlP0WJmoVjIiHlAB44xHP/UAAFN39gtVczmY/qTJo
KENo+7SiaGOHxNNtCcyigDxLF60r/koEZ4RlVViXvP10/V51dIqqm2PMudce6hoMqp62vWm1dX35
VWTJ4uE0spw94on0K9pcgm0yxCd54PoLYbeE41ZbCQDHnGgFLnL68pwFy0eDbIPEdM7N2t75RMK/
CJfvzQnnvL9E3UTGV27cRK6esOh0nd5qtEiapN2NGLzKRiXfncqx/FoFZ8Lh8LO08LWGziKmXulp
bScg+ukP1nqsmf+GJNJMV5xEAiGFmTtxAIrzj3BwJeZRYsCzjVUk/1az7w1OfRul2ox8vSksJHmW
QzkuafShJFD5udDqaMzTZJkypud+k0XohUPSRT7l6M2HfAIugj/gLimlDY3daMGq/StGkd/NB/kw
brkNEveA4O/8nEY7j5ZIH/9xTftCE6apzvj7/uoSB/avTAq7kQVJi2xbav017vgJRbASkycHSCTH
3jYNIj7maWC8F9N2GOgGSJ5oy74AWWb8+E+GrKFXC0mySa1WZBFkxTJGHJUOqL9Pxh69DDMQ41Ga
xcX1vPr9PBJvDimTaQoHx3hjSF3RqDaeTBir1Fozn3y/b1IGcJyvXlxlRqkMcewO3iyOYyI/gWVP
l6wvtxJV1LD0WwLjvSJoMysRbu0lLz6e/uXvSc7ABTQffLhOpVXwedGSw9gnBx59YRNYITXYJ7OV
9eA6fg2OtYUJft1qqacK332/OWgqw6italNNykztjKaVEg5scT2BIfubcwQlMS1yCTq1gm/fYO9P
z+VNYsCU8DmNx/jZR8FBSgKexAwm+E/4rZ3vpWOKPlVVGbwRq61mFevqgSckzJyi3NF23NPeTOyQ
twM4/BgVkNAqB6/bN/jZAPkbOmW/81OfUZhfW7q2uGDYCpH6F9k8tjf5Y7lZlCNYUUbyJ/bwECOJ
LAa7wgFC186asgklgnwRddaZ/na5r8C7p7+9+Kwt6dc0HnbYbuJycoGn7lYNYVRhboxnP/iJR3+N
B9Z0P1G7KoCy8ttz+0vF+O17C484LPhl1oE0GNkh1aFf7cd4AwU8EuD2DNJ1Ntq/WOr0cYL/VPTH
Dnuq3BNn4m3wWA/P4Y3xZmYcfjLloC6X00EDEJlMsacliur5dQwMDUbUNFlSVTaIwJriTWRcxlkH
tsBxI7fxGVw0XuicyntXBthW+K2M2onCs2b62WVx/nBb63YVBIhEmHG9ML45ge5iFVahtrkZAWsb
7ZErkPZQ3KTfFDGBjZLKtdFG5IuDraa/AuYVbd/p8ByVLFs0Y6wSRjNaYriMqElAI1XUlCC4RaTr
FzvzCcMoWpKqDRNJcw8ErUX+HicaRtg/6OxaVUYmW2mUl48dfe4RCcuVVbm3nTgPMM/Kv14BLldy
7bYtwfXkhJZjJYzHNMS77y1E+oPBaPzkXitWgXaG/dQEMke1V/ewxfTfeR0+27+Obe5FlkKzh8h4
fe+NVF3YxBzRsO9nhnUBMiwjUipXUAgCklXMKgmdKX7nVijLILqd0eKuJpwLzeBMbpS+sXPCAKJY
yfNDqfRrcV8OXNcX4rmdfFvWev4zv6o2+gA+v81IBl0UMShQhZ9tfOQnvLGMMtalPNPIEn3ufNm8
MJ+3ijVPtW6X2892DDKFky8C7p2+Wee3vzBIuv+FSl/3dmkLD6pSvwd5ySeQKTHWCXB9ugOjRIUY
cBZ+dMiXa2rIYmwAgMO8W4LOsgr6Nj5gpsDYGjtG9z93NUzSCEGkPhyegoz4cRGJXgDKTDXY3Qva
pCzIfJ/KhNM9j6Dk3KRtTq+rxQd0ar59YgAuIOZYwFqPhBJyFiuw9BZ1SwfNm8pin8A1Kt6ganJ2
gxE8RBXKj33e0k9XzOQDjulrGQ9w/h1FqXiodlS7Xf4eLln3nXNsw1s3ntaFj66Z6DgMr2sY1XTn
zcgegTtRT9rYt1ewLCFnda2KuTsf4Vp+9zjx0hAkCoaY7trXc3cz1gJpa+TOj3FZ5rg3TSNlAmqY
y03s0wOFNSDkUigRMLwX88aTJlOUjHJ0jQA9WoYnmAK1m9G0HM3PnVj22F8v17Tej9VReldBaH7k
MlgYnDm0fTKK0PGwMuwRhsgNL+KOuj7z3ZdSg/iCoRpus63i9fFuEAb5wvxygriY4EH9ocT9tI6I
6/mOUjlxiYhd2Kqwgp46/GHFmN6y/KjPxFy4YmArtQwG7tPRdkSvXxAaQBqNqWQKkdnDIFI0idjD
1z1x6gF00faEOPor54wgolr6OnGovoZV+K923uX3edsPrzxFmmU2FEFnrJxeQwNMzhAn6C1K1ZWw
FAfZsmmx79DZuoSN66KTi4udqdJvRJKx0kNzzyJjrZSLLgKRBekWQvihmwAJPSfqHSyqAS6/1/Gw
5aMqaYQVocCNTlUnIQmlkIpWK6Vgjgjk7Lie4qAMIXe2bJGmwbNIEqra41Qldk1PusLFO2N0ogeq
47fi65HfXOtgTpx2vOvx1LzYOv4BBLWighYRQnHiDI9hiwjaB9ZfgXbOO1To/TEza1/cFEh6kaFw
V+bEYw52FX4UrhZK+kPnqFWjBjsV7c6Ckz6mrCkHU3Rrl+4h5oUg3r5GqA0am/LK3T49WkKygMpn
dwzSRlHxvAAcEtCqjO8ioXt//bOswh9dv6P9B4Ho/sMOivTP+wLJ0TVJK7b5V+zlSPwjHH6ddctL
eWpK5EGS6vyvPTca5JB0tQoQcmXGe0JAqMJ949iRo1MQTw9Ovog2J9e8pgJVEqpfGMAYq8OVhnj5
tK/04AZZWANPqlAbh00BK50oAgNIG1HkYvvhmsRTInPgcOUjS0cgMmVUZZ2vvKhxXsMtqRayr9yQ
Yvj1pnRdNk/5IX0YdgPCMxGDCca6wyuLyFRYL3C8NCwG4fSabQWJ8uHc9usYiJCLQMgcUbCB4v8E
QGu0BTiEktGVFLZZzu5rbfKipaPPH+EqgES5NvjoXdg8pRqMkqDslLpND8Zz2MtOlg97UIyGWDcn
/+MIE7gXlF+347/uBXRoKWylX5n73zsmFwjcKIPTj31MK7IOtH2Fyo3MLnkRgZKqj/YXLhqLlbWi
hsiHltfUcNZwFMCcHAXBdDmk3LIIz0FswqOYoN8YGkcLUpIMSIZVSy9oHdYzDWDv5IA32OSqYLeR
NJS3IQnKeYoZ/+gxkUr8NMoppPoeTPgGvOkRhLXAbHas01UXyMBR/rNkFRVT6PToCAeu7Qr5w5XL
tjqQ5oQaUBIuN0xyRM9Mqu0k/DTqNClaGUJGg5khVRemOhtDRg7XzYZq8OYHYGpvnonlkRfdG6NT
qXIIKhfBoPfTHm1kAJNocvDkrmMKimghMZRM9/9XMO079Z0ZYllmrXwoT8kNs86/qC+8UqSON3XL
096bz4GkzpE6/EYw4MeUKaJ5KZRk2OV7L25AXuWtH0/zbqw9XMfWiH2pKTC+yF3hONOJhaCpDlP6
0tOGOzfIo6x8WmLGBsK0uvXcFMX254W7z2t1vMIJenPFw3bCE0titVsyHvCsETRdBviuy5sq9EuR
XORJC49mUovfr25M1CT8kCnrvlNKU7c/EcTcfNHGOQti3GKTJ2/+WGWaQSby/Hwq3///UrQZwQ9q
bgfqxUCzjVkn4yxMB9xnmIYmImtJL3DwpZtl12k836swCCAtAdhc1eNxyKzOSkyUhbn4qIpSQW/I
SaRcu3kp517y6QpD2FGntrPuM3u9r/4JpWq/PDrYfv4ubpmejwUviacnEbi2gQnEjwYF4B5BmBqy
osjNdg/bGdUBBkokALnFR0HTexvApQfxYTGn/pyvcGf78+C1pdOJJ78dkrIJE3DNBT8BvevCdb2M
XsrCXsRV4OrI+UkMElOxpgBxtZos5hQBwsNJ0EK88CxQ78c6OrDNKl4wssFXTgjJp5i9cvrtP9gU
warPFWMTBWAD1GjfoRP8LkWzp9jriNr5Y0n5j2tUVmSPt21sdD9bFlAImSIxnkawpLmYw4lucLAY
xvetvDBOXjYLg0gWbjYcNYtvNE0b75vsA/efPSZ/dWjyieaorIQZAYjQ+m8LiqEKRgCdox+OvmKt
Ks2PVaxVOS0cCreHKS60BAn82GL9rndp1xOxGksN8GxQ0uc0x9jiHdSgAY9AuSTXaYqMwgPRMASw
1q3IR/ODOYd5qenX3NLr2fmnnBH1C9B7axIJE+9UlGVp5WCcKcSHAMop7+GLxk+yguRqYM8w0Xyf
CQIg974B6LvqDZCeONZHGum1VRkndeFpiRCHFU8HvEkDZfcHiZ+5Yt8ZIAwvQ3xQ7JdngzZ24TZd
lviA8GvIh2tmiNQvRswOdCQo55pMcpjZtJIgeGJ0gQRX14EbLmQKABBtrWOqEfCB2CjKyXG3IL6D
oAEJdN5BIondMgBo2gQSgXKjrshJMmFWQ651f1z49/IbFA/ZeeYdSvaPbigEZnhSG1CC0sjfU49D
bzY9Sz++B6uyB4pJSKxc5liI0IihJ332paDapGYoFLpg5qtdxgJ2rf0TEgwdGvhVAEQjAkveGAwd
rIdDf1JkHN0U39mFlyMWZQnqAGrkAXF9mBFaNe0sMxaP8VJGWQcKA6z9GvbunBRaqURB8F6kobJc
byUd1N183dbLd9nHIU1ah1RouO4RlgxkD5Jg5ANT8QAIw7WOVWD850Efg00PQqX6pyuuFAfJdFwu
UDx45ZK/mOG7B9iyW9R99/qj0GudIIHFt1IpTkUHCiaqL5Umyb+/sMUVC2AtPYvFPudpDGlUsRxr
zG8R3SuxYtcB2QSOHy1PEvHnne+zttoxchrs+pfSv4x+UsD1ZzRBJ/gbDyecm6wMnkgI5qK0dvg9
gurq/4AlifuuqWVDAbiiVsZk5b+3dcDrE9iPEqo215xjQFVKcVpKMgZDtvt4MWQhIVDTb16Wd0yY
llOEkytrRLOBER+zn/mNWpak32hTHeK3Qe2Gm31VXL9mfXxwph10uZYeiAj569EWBEmYPe4zgitQ
hwieAr+geHM312ZyazKGeuFYbqAcV6p9PTHgVUagmo8NCtmL2w07CMXtaFx8ZB8wnakGCCa6C3VU
u7Hczl5ph4UWeq74RlfMD8lpglXwTlip6w9gIRtbN281lMRln/1ZK7nqo10Ma1YMILDhMBhApqcS
4CcYpPt/UrZsnsOHYPh/fodEhdY3mEFKwaolPjzikiir2c2dA4mfDc2XcV/Nc2Tk5u+5/36J25eT
9KowzzhONzee6ETrLyo+c5ZvTcPonjs5/e863dT0dshNS9tGXv3LJkpUd1P7OZKulM4dAnxU4TeJ
+avcYD1bsVvOJD4XkGuj4xNrNrnHt1QEQhiZm2rIefKL/NyXVhA7jRmSKZBPY4faXuXr62is6dQA
rgF/oV8dF6GNUixVESzPsRMNvW94sjK1AEH+ez3N38RX145SNBuOkvJMAS5gEmQ9K3GeKqcGQW0O
V8ZXoI0ODR3t+eKfV9qfKyBjXEHHBNzYknvu1Fe8pIwGWhXokjFHaKpD/kXMnFSPzg+u8jvPTkTn
PLOk3liPYo3him+r7gJxyswvnIXSQ/D9Sr73AQvIlMkqXFYCWeeuKC1QhJF3JR+859agaiJ/2QDE
tiTgA+UX5DHE13m6PczgVAEeXrIwK9Df60MXwuZ5VH7yKjzdILhTjB/SIprz1z/WvjUNvN+7JG4P
FtfGvENY38UUu1GcS2XIV9Lhl3nDP2HlWK9FwM/rGPYm088bZHXI+AcvPtkE81P/9NMMuhLkazmb
EEU9VNiUCZGpNTvJbXdk5t0sRs+bEcBtG6RcWwXnLY7Y2HmyCmtk4QP3rLkGi85p8JoktmixyppT
tU06W+EG8TIXlPnRXJUaMz8jv/eaXmZOdzAjahqb6rNJ90rDXDGGdn0V2b6EHFfA0JARXCnka1Zu
YOqCV/VRvGhBhhN0P7cbEDfL0g+l4xDBa43TPikdqrLnz3/8GJAHrcn+uUsGpTcQPUDgz3jZkPI5
PJGcauwnuECRL6p6M7xKD7mUDhANB2BFlgIsax+Or1E0AFc/dq07K0hklM20ImPuVxdBvwAs8jno
JCc0vtuBSnNBF31OfDF8WmlX86QAFKcQJ4Iwtt+TwKp1Netv7BZzogVcfTbaqbCmiLsKkbqd6xsi
+ACHXtivnyNCQ96GTnR7uE1jzKMf7kS+DHsD1nsvTaQjscdtZK3xgXmU8jbAJeoKNf0jiUH+xhU2
sj3kkW2d5IryjcFPVtrMz/IIp24G9YZHyAEOxHZ1cr9Hgd/zngw7sGQ9SYxFgX3T5zVqUp3ZAnqm
v3LvV/ORtbh2WlXZoonoPnFDK9U08lqlzrDdSjmmpkfLkmvT6HDUDE8znw2qhnLo74YcMcKQikTA
MkPF5QFoo2h5P+sVLEIVDCJEzCiLmAS1noBXqLRgX3TWSuNLbakZlTCbYJL+fzEO17oIvEoGxzEV
jtePsBRMarh9cWrVsjq74q3AUrvjTmUbeM7WK2ysJ63u4YYu0ozY6mz3ZpYS3hcUEIrrU3UQ5F1Y
KDC404g3CP/wASw9skFxRAXX4CpSTXTpqOPYpDSWfR28wmxr2BBNYhxYkCP7m32UpfJAaKwwJJ9R
jDBo59veolgzO6fRuQwdMF+p739sXUIP2E9foqY23TYgUb+JL8iR6zcgUGIrxyS5jiPMrs80Tcsy
t4uRWS9gMrYfwT/rPxihwLCG4Pb91X/CmK2ZNV7623+hLEmS4iWajo92v1OLXaoATDeatKV5Z8Ef
zrKt89mE+aThGwaaXsio3FjDZ9KH4Ka+l4I91mmnJ+ro1TOnywAvg9kEdE7/wX5+Ed2LJlsNnvye
c05s1zEoIl8wonrwlx4XmCdwIIvuNbBxAxKCHdgggd5pvtx5nY6fi4qhq6SZCiJsrg1GYKGIzn7M
oXqstTwDtSgBAbrRoGBEK8t7lPU7NBLwrsPi68qWTKXd+x2J5AWQ9y20zgW9vGrAsJKxwJ47svK1
Y34eb7mFksye1jNO3Gb0BY0o0w1Pa0XmOsQbuPts6vy2xSNYNOn1do0dXGapBVVUugS/EhJ3hjl3
f4DBI0qKXTheeRNbTzNP1THsjFmqh7uTdNFvXjZY78PhuQ+dg0AL07GxEvzue+quQWZ+fd/SX8dY
SFhHix2MAINrN7GXcLLR1/eyyJAbklUN5E61VHXl484LzJ6KFdbQSbSsi+3bQSCjlTFORciwKRX0
0J2/sWSO0Wk71zZC1rd3Hay/dRQoS+IlzmkvVmkyjb3pKIcMBfETXbQDkQvP2lUB3twXLyJKZ+ud
L7h+v7eM422xY3M2sITvjNlsbIUiryxOpXEBRaaAMD8TwctHmAlXRiMe3raeyCNHka+8NnYfIR4C
ISAY/YUkm1ImTgvsgIruj49iQnryjaMjf15Ns0NkG9UfaGRMZKpvv4w1OFXaBZPROVO30i5DiDmb
lvlAz8qCE/3Yoxtwujfl0BnEAJEaxs59S97XdhAcjgutWiP0MPX6aBJJ0kx9qrC9jeoLgbr4bueB
mTBzJU8kEmbuQ2aYmIJ/3t/rkGlrxPPF9qzdNmqrHVyUFL9tCSlClBNfVvTd8qTitOqNR3IYjTFG
58C3U1oxaNgLV8PdQE1H05Mx/co9cwydH5N6aVzh4KklIAGsphYl88ldsSmd9VuJX2AePDDWsIde
9IBYXGzF2BYfUEWjXJLWN1v+TfRfAWc7FBX9x/VC5a1Kof6+UbdwMOEyDv48zDtoVQcY2zZzlrG5
EFLlI18Z1ZXHi0nZVLwXH3TT+twMkfeoCLPpUP8WASypoY2TxMNsFhzWCsMBuKdF/Bfmag4nYbX1
GkEUoCvpJ2Xjr7xtIz5F0/6a5kpXqXWMzsr5WtRC25p5b44Di2SfAGt5aP9CknyaLfvt0M0YuNDN
rbhQuRjrRxIfElkr1to5b870wSDItyfCun2yGUhPpKib2vg+izBavksm1GuEfaOE9fjPjskTDdZ3
jio3Iq4rQZI/wi/yFDkVNYf5oKSqn9iN9L0L8M6PVWEN8/QLgAhOHZbS1NnVB7vH3u/wvokfwh7x
z9P5d/1KmhJOO8qTIL56nLbflDFkGXQpo41c3C4iuVAndFZ3+c2HiDplBdQ46W0AJzbGPLCYMLF+
GUM7PD+KezFgBuOsB1P9a9ulfF6HEDOmbYbR8PzZEfhGP2wdRJmEhzcIQ05bBO+SHCXbm8wcpbtd
dRZJEADE/i/U7/1YE4SCb2LvcnnBy+BHNa9DuZJxuh7dNojudVer7hU5I70lAgGlZSGq87RQxjOH
o5K8ySt5QIdKWMQQKhiO1wlolZCl0+ZJZjf6hkYu3iv7IIdy7DqCYjW6Bk4tgxqG/WJgUXoWHodm
Af8MAIVXHUpwp6HKy1ObQmrgJW54vv/gX+w14iFJQMqwJ1F+3j45ICdNq0ufrlsTYbBpaNOwJJVs
PRKagZGsEKhmcE/GkOiu7gwA+kQqVwf+p6Zc99s/W2HiTznbl/ti0+scsxcf4v3AbYkIPIg4tjvn
vU5zcqTM5wo3GZNQJVFfwOH+lW4iYHeK/Dl43CEEyzFWIBEmL1U3/Lhi9QNbNONNZ8VlkjnkPhnz
Oo3t5RJ0Tm9+TehCClbOTP1Yhq8Jf5+5WDiTCX1727QvNQnJjT2+KeNZKUSz7FhIUeU9o3ETwVRo
ZImIDELlhScWwE7nFeHwAs5vd58w+KaZdVeaXh7slQRXu4/pMPjLCLul6M21DoKxwQ9XPkQM0Bi4
cTMJUWBRaOLMWmKlDk0wAHGkSmtWtlZIJm9XHUOcfp25ACPZKOOI4k71cIZ31qW0n+QB4ymIQXep
aIPPuX/NnDuVQIg9JKjPTcxoOMRJLLjwprNJ1/GqsqBEv+JfAgJuCiCLGp7FeQt7vIc7A2NDv2Vs
u2T3ZJbcvPlKN+lqmEDHcbwz+eVURm2NH3Xfsm1WpIXh40fXyqi3G+m6AQDenEueMmkNUqZOMZX9
primHjDnSRRWKlqCo8wmP0LJmzWYv+pWnKtfru0xGN3+bnMW0WRdYfcajuAbrUt6WR9cjdPhdoMh
xYUQ8f6K4pqQTmEoWXeSCuUZOarknazXFyAG52J1Oidcn5fUOUSPMpDj0fIy8EkZVZEnVXbSOGRB
717KUujos85Oi6KBMNtIOYPd4bIrIQGKjTnvJfi9EveHxi+f8n7eHCU6zLI8XCW+mDLBYxxmHF1I
KoymrPcK+ku4sCfrPl8ToQgiXvfN93arr/FZx5DLrnai9ubuhysBYm85xbcxVfwbfoFFFEL9fmlz
GKS/KlSCrXqHoZ+L1I7gyH4bIur7wBvf+Thjr0A7b8NGBfqz7+I8dTf6neRzzNXxugHq4G7uRYYS
X+sWOrJdsxAbclZQ/QmobKdS5GaQl6e0rFIRVNUYJm+TNN56lS/vfhzshoCxpCz+ZRzxVjxKJZAP
OHF/6aUk+SqBGrH43v/Uye+vPm63dzo5J4MCQ5vLFSgFE7cOu7MNDHrWpd3O0aegzk9WPKP0MKIW
0y4vsMAGp7bbgaae0wUXx8XXVIMdYCpXfMR3vP3j91+9JUWHa7bq7m8vmFPxxm6P3SYc1h/uwids
0XFIDxxlZs2/Ak1VdOAlv0zMqFmbQ3MVnAthEXAb2w7ywuXuqkPkTnLI3xIYgW/eL29ppMT396c9
BY0PkwAaAmf+Ju/WsoX+uShrI702iSZCX6dAaPRX5RkZaCqsGbNQekgvDCYIgEXAY4yKxmrpdimB
F2PXJcFWR4LXeSibbosuV++EUm5xTtxpXU7/YMdQGkRKQAMOW4OMlfJJFvU316HIKB9PDRJsfu3B
oeDaICdgzDwV1S+5KsRVfPKUpQLPmiTRINGIdf2LDZWtH6Bz0G9zbRxdiFJk/dhmoB/G2ASBBQAQ
T6WbBc00KJKXVITyYNA3JlPkhT1yKwKxq5zqzDZIpFqCXQOjhULFBcllx8MvoeqQFpCq8NVaJqa0
UaFIpgyPP1ZKTcISqOBa07nMCz6ifVugqzHFXmd0vLQbsQ/VfohIwzYKpJo8KiibXpfOVbEs1v01
9L7LGMZ6hoN6PHQQYgdZaV9AigSWrbX65YFp7LaA5Kji70bFF+PCXxt92Di+Ebjz49Mw6s22iu6s
Y+LKzBvxjdHXQTPQuAeYg86anr6Llt8vRZO6IYha4ujYNvd5CichVjRZc0dntWfiojbyhF88Llsl
+wV5KLBFN1/KeimEtET/Z1hjuv70DnHqM7caW5LxrDMnCDsl4fzZ1PPukmO3WRETEmCFs5Nw+0n6
r9ElG3lIKn49d04o4Pq6vcsUEgeCBM4ZCkNxDBAgNJ5f47aRa7Gk03/Bv9unBQPlNoxF/CZ+qDX8
IiytwmE1+eJwAg+LcUFQ3xr6udzdpA7PriLqu/4UTCHsqB6qddOGeDqBV7jmFUHMdS3w5YEDxv9G
GY4HyAcdTnbOUtVMpWDySJXoIKIEUtzR2W4AQv4LVOOBJkgqBK0poWPsxzDcX6Y313YXqsZ2+5HI
oi6FPv3DLXd85grmxlq4yynkPBd+WSbKCM1g5WHSE1GHMTRXxilc5YfuKlVV6ayQMmqErgMoINq5
T6WSee+GcfWXJg/vIKAwo2I5SaOMTPs5nKM9aL9Bsid/rRPgX0IMId1f1qszJAYw0FD0MMBrJTdE
QKK6UikoD86lKTvOdIidy9ggWDvpVbk4bfGIUhHy7JpMa5Z4WWxtJpr8gwU3IJ2Xzt9XPuvYuB3r
3o6AiAqsignkK9DoBfIwu9hEiVmLfknHTcxD+ohnF4YmKHB22iYcqu+9mB1ypBeZ/k5K/fy9Dntc
fDkHvDKYksa8YTVFl8jPJUoOQLuMNlJiqA1aphgfTqsxpkaRDw5xN4Wy+2YSSNeL11XN8rbEWAVK
3F3iQQpWp2R9hhL/CnAocjQlYOK6/Z9vELlEJqjq/68fwawHHeaB8K8v2ztewtceUzCg9+mgxWbn
hoZVUINZXQiwFzkkgdU7fCQDq7rfVTlnpXv4IJoiX6FN+0V6gFFuyp+h9RejaGYFHCdhUI9ls7Cs
lAxdJjuuIs/zUj4JsiknnrAyDm02phnRcGL3p5imiOgdQ/gXtFzXgFghsF4El8eir6NJu680XRz4
kzNo5ejr2iVWI2MzxVPh8voDgX7yY32unpTeY/pDVso77Uaew7JGFad2zoVeMqRa+YkZDVDErtSV
bY5JAskHLx/BhxdjaroGcy0YExpQeu7R37CGAUosRIik/0cOVR6AvgX14c+t4fDggT6WLZRrTeEb
ooUmtHJPiEoAHXvlDDxyy9jd35s0XmYYLmXp0cdTs7Aa2UR0iKE9cYvn8ryQ0+VqZspFqwglLQro
8L+tNxtKmV9AKWWYR+vO/34FhQ/zYTe708jypMSqNOCrj8WvXPxrAMsYa1Xc94iEpAwoksw7onRI
C7ISZ/0DlPYu6ebsaY62MA7SjmQsJ6Ma8KZ9pdc/UiptVmzKvReDx2zk+m/WjqmR+ymdFDvPBDCF
bvW5dWDQTie6709ih1NJXc+yfkuL2Fim++ujEyJHLcUvbob+QDfCZzgIJtWZZfD71YPVH4/6ICLM
EW8bwiQeG+FY9acRoGAuo7FWM3pQ9+qRW2lFV5t07hYSfxzgxkBMRxnnEAvzZlshuoComWoSWkxO
ckeG6i/YIbTEsiBWSu0VAG41MV4aoE6Tsiu7TGcBdAFHoNPs4YtiAOVasylzJ7pRjpopzUX5mFT5
a5r3WiVRELf7WfESuUKymOc0Su65wMfh0c2LNr+/wAw+cC4ipQfBc/NGBo4tL1Nc7TYE/VLavMoz
ARRvDuMH4d2C1T40RaVgHPawrW6w5FTlc3UcaR2QUoz89ryMpsYVhbLaLxR7BI+pYDQEshcFKKKN
j3Lk67oQvWY+uNFWX2TAiMXFIi+k97cwrjVim3fAim7jHBV6DjqP4/HVcwpMvlf4ed4m9y867w0w
fihKDBGRrdESkuDskZCDNMhh+G4dsbcTB/bfmk/SrDvrhpxApFhW4P0dNF3J+Tnu6vbNeoOFlcmI
6KQlAuVmLjwe6a/5R63dWleDFMmRaT9EpFIdq7cwDOxsfU4YZqtrqPkiZkcws2WyhUo1Tyh/tjSJ
gaZ4rsz93eSPZhcZHnc3zgoPXqSwwYjnHfrgoq3rfvOn3dFwItwI3iJr7b2KiPfAb5J0lBHrKFrH
iN7tUobfcxPsooM//90UyxR6KW7tArko1ZZHPD/LmzQakxnnOvL+ExqhP551nWGCJt7dvKDDxuiV
136aGjjpl/QLN4GO6J+d5kmmqxOFdSWOFLM7YyQB/UNDK4IFjChckCadXSdp50DZ98ccxO1pFv5M
VHmsH5psjveH3E4aLwsefssQCJV+5iaTXZkqSJJiaJhEHSPaSxEbCXIeol8sPXLKEDaLjnY7SshQ
tG2cSpZ6NJoIwfQee8VESAzWal55z3zmSvO4b1bn9/BZk2YEOWrHRTLAxsncJ2cNAPwQUlNzyanO
ITiUVsxZXCuP34QH0dq/dtJ/S9et7U+XkMyEDI/XON0U4PYtkl8Ufjz/cA9bk9NqAe8E5WB2T/+I
aUlTVzNu37xeUe+pNGXNWM2vZCN4WpPFEtpPsv3th1Ki7WSjl1YBdmQVELt9yCbPHvl387aPinTv
yoc4Ku0IX7s6LSLoH0l9P7Ll4sCwV6m/oAG29HEJUZrNHKLnwSYmdhrXFNjSyxAGHDnGVXbfsPmj
lo73vaYoeqrRz/UabxuKJf/f3ub6ww+ne0+4CDDCC8CgaSw4LewYJYAQW254BZM7ZJpuSQXBeVGS
uFyMX662JTRtgBTQeyFaJ2DcQ0Qzfh/htiDQ5HebMqMUXjS/7lyYJYCBL9a4B0PH2NT8B6HKcV+0
50fYZawWaU2eLDzBbVnrBFjqJ5wr0tOmiR2YP3VS7ygrNG9aJ8stD7fsKAeVdzkkMl6DiNo5j1/r
Cxs5nv1JuIsVgunsqXkddGNEJpFoX9jBG9uW/AvdpEY7AA9NoTsvSwhPK7qEfePUyAPvrFsjjW48
aTfiJjJcCviPpSRbgdWTZ2AouKOnf7SNAiUT8dcG/asydHi/RHH6pBtMpAuVECdTvWaUwEIjMhT6
CFfM/SphN6cTqnTHQvVQ6vmpXpefhPgGpl0hR1HjHsCcr1vf9AgDnD6GWHxHlL6XzD/6pK09rute
OhfjnTufa+ngbdlPdEw86itP3asUX98R7lz0EHQp/ze4cP/EZPNWS9xpNS/i28GhN5Hswr1uI9Bu
zi9rWNrGiNPzWRpumBance7JL9tYEzBNrC162U8lNvJK8ADsYOH1r3MN5PyGDIyhQYfqaRURDk8n
c3rrB/8/1TbISWZvkcsI/oQBS17HZQLKRArjKT4+pt15wZDdIbNDiNc2VIdkbOQ/UKpo0vrAq7TB
iNUJLxmPsj9HG/qWZMLOnYUEPBmctQ7TrjKBUFGI1MDJoh+KQdhNcn43CGAzl/yLUYv+dpgsVapX
8FaGhMK/bRAOw77kYl4pnuRVYg81P+u7Ct+an803qhWSLrqVkCW+g0nWe8j2uDZtwIANNV0GpVgq
fPrLfgfhK25AGUmV6z7TU8Q5Nu7RRgm5C0N3hR9sB4AnQhtBJmrFFrTh6q2DC4ff5S3P2w2CaucK
WHUdC1w5MN1Q55TfRxErpr38t7q+n1AxyPUqRB8y6+tiuCQ1nO8WXhNGd8dghwPDNU0BzpJmQapa
94zsnIUk0I8TbRFO6WAwwrX2mHFKlBbGZx81uQftM6xxvRhd1NpWZ8GjZftecFi1Zr0E3tp57Cwm
TnffQbRnuuOrc6uKYM0193iew0NG2oHzoxaLjieAlsr6G35nPqaafuxZXcngt3w58LCAmxpErUky
C+F++19K9BqB2sakf3+EmBOKC9Oj7Vgpl/hA7oN/ljuBgzvoXUMAzvLuI5Y6i72K0AyfPWQryLIT
nhXls+9f08FYC/xEJmtjr9RpeFHYSChzsAmEX1L8xd5lEkBD9ZuzMTQ9pKIAOygV8Wmm2IFjYUZ+
uQqJZYRtPzr3NQW6MTbRONwvqQq91XqwGzPzLdttmmkir5kxnhe2fhbaJzWiiEs2l1TEjrF3rh6Z
DNytvyCkZR+isU08t+sj3aO5MmqtlGAGLMUz8CgHxnGjYFDZW8YwROyl23BYjEVifQn7VkLdEfGB
ZDK/mIGF9dUDFXCbLllpZ3gjFjHXbYeWdsTsLRo8ie3dbxXy22rpwpxP16iyz6Sr2H0Lr1ty3Gd6
p9KRr6qfQNVxEySIDnVx43vocDxfLj9MMR75ZF2fyjq+djwndi0MwkqM5fIlW8+4MQf8Y/UAh4OR
NW3DYjjjYfHHnJQiUQs99C9SFBcVPnEKKRHUh7R+iB4FwRF2E+w55PZPcDSsTUySceopV0CyfgQ2
4dBGkSjgiZMtDuapblBNWWChG/4A8Yqx9R3qGi4PbDYz75jiIsOzlI487vQJ4BrgW1tpw3pbOM68
DXYuocCYrzp6aa0+LHXv84a9MDGmE6In3G0Gxe4SMCdNFXSq3ri90Xw1+Zk6Cbu8LKH6uQLqzUzl
3uKFG0OPHPz7XgQGPMf4ROKh05WvdS/4hDbDC5+ByQXgm9W7puFivf2dhUHM0dAxJCA4hl57KCQc
6IpndBKui9jsRx9TFT+G4qTtpdtvFVzNlq/WubscyEVeIHsMPKcVIvPmzpnw8ECZlOBklt23AnoO
GBWFVdWOVOFJyC9HB35VyvCNd4aJvdO922n5cZC6eK1Or0BrjLFZ4/SM396Dy+9PW2qpuENocWmY
B+etr3218b4YxhWmJSdQHxoVYIU6R17agfyj9xBsB+KzUDIMMEVB9OI1L7rHYbQd7XMzSXoliG7E
808Xk0mWzXKYnLpbPyvBMV2KqAH7j7hKWy9sV8TLx/DRf8UzOkRa3501Ldtb21Zr/Vg0cpyKSJEl
Af+QZ/8PL7mZV9fo0sUCUU8SSG/aro5vgyrA3FK/Lto+iUnlMjHhiWmBYFolL85YFbJ/m59vMtN1
N7pkRJDckdG5JFZx5RxsCVpT8UikxdogRUDG2NI3teG6iVkKr3JoRkTrwjBnqfPkpjOMj51/yz7i
nVaWIgG/zCYfJZOuynwd6Avd/iFqFHyUxgKW7EUyjKH9sijY6v6qQ6c4g23HVuJwuRo0YNu/pPXs
rFL7+6wepzQc72X6aWQebxG5U8uEC0n2Iy5fyGkWQXoNNwlVTKqnPf3KkVWLBFWdeOZy/VP3e4zF
MS+0uL4+iKEJx5/ODPMBhNinuFa5ZDmkG6dggjerhLJqMQifF+JkDtR1XZ464LhxFn/hw7VoDCxP
ED6Re4TjqidY8B0v9MeCJGEPqlmAOM3C3/O6ihFZCuV2s+lc/D27M0PlpC4zmdnrj48B+ZeEBQ3p
N/SmaifJYnaFC9MV+7MSS+ngwmMcIDN7VjX5nAGEt4Y85fWzrG3U27tFqP/TalObUMoNKRqVQP0y
VZ49KBMONFKJCzjcrZlkM96IQ328RTM92yqYWV+fyvU83My29f116LKhwrE83ChnTMqxDIkMwYkl
x7fyFT+RW8TRH7OhAoBbWO3CH70Nn8AX29FhyA4LlKATBrUJOU5EuuJHEbTUS0Z5ulyAdRsP1kZf
ZFOGTuQ2GUOd5VHAp+B2d0yNzOf+qWZzTl5wO2/yJP9p0G+YR25GUUJc0tUE6/o8HFmIPqLOZwE5
7GKOVASYnnq+B7TE6sOcbbaTo4Y3yGbmx2ZNXXzj54uFzJb04hBmHlmdoO+xfD4dI9Bplv+8/FY6
0KK+eCpBH8bxgPrzMTgbEMwyQjwUI6KeTQ9k3WQGwf0M9Vdukq0/rCooe7jq/kjlyMPdDVLXxs6P
qMR7CU+3JA3hANwIw+YRw/tykcSeeEVDyULWo0/CwRiFaHb3hhqpoZEdyIAXKpdHU6sObxUj4h/l
Opn93GlGX3CH31gwq8tP6Qo5Plt9YLXiYxO+5ylTwCpkkw5Q+PmUJz+K9VRCd6eZ6Ntk5bgPUUW9
DF3hpwgj630XPB8Tw/AL4AyTkXewjGhAXqlZnJP6baQY7SseFrJraoI9fIcJNg5jNQ2VruBnQbF2
d4FLsGY/5H+EnviodD4yLs+vP8hmlrFMiIyorlZW39qIN4/kul40EtickeMroJUVQuPHZUzWsPj6
D5ohmGFaiOc+sRbnsfP4fDeX14DSKKuwAY+jjRmz0tnPaL8xL1OssDfAVFy3TPWHhfuIyxgRCUcv
1hy5wwIkPVORf8UXooKd+vK8EHroQT/XQm9aAvFgtHNqoGy2Ntx96JV/DzgynsZK2ctXIMUTHXx5
UNln6spNU9WApX4fgxEyKpaCzwfyvMQFlAFSX2KIW7nOIhgikbJqcWtuUDh1IQkxJtdF4PY1GWzO
WtO7EFa9T0/x0C7UU0q74UFOb9l0z8fPYXK/M0R9ALRFvga2wnY5VQUYtTMN3TqXsXJ5ubzEbmhL
9PLQvKKkrohpkF0CS9SvBSMldlTQGYJJSKUO6+cxke4p0Yz35l0bXAVlNvH99D0DGNNVtDpEx8Bb
KKS3/OLKHl3nOUD3xLk3QFltENzXQxXPh06SNDN+ZHpniJ4YOsarZTmxDTnQkQT7xEHv3G3MdqE2
fZ4GB8nKezuod9qxVh8jTNw1ah6+xOdOuhAdm7MHcWoJVIOK6lAvDUPplIycxNrIvNJL8XgZ0Fxs
up1wgGBqf+YP44n5eQKDtIed8GD/RuZ3DQZAH+kqqLiGb5y1UZsViEirOrS8kRcVD0eorWFY5RBU
wixVXe6bOR2UNiR+c2dh/uieP+4M7x0J1JWE9JUnjecKdutAz+h13jy1CDJAx0B1tKVp+MIWIOgS
OnepWT4MCLoIyT5t8L7a1hS/2JsgahguuEfjuZHOmexqpTF3Rl6Uc92KXdeDzQqbVqnuMcYmHXpg
mnwycM3zqLlhmK2R0RkWRxelQnyP6wfCg/iz51rNliea8m4zLtxoC63jNW8+QRwunB6Qh1xj3CeU
xSMZ0dpkYXpL3PeTM2oiKSY6Lcu9wveJEhVJc2Tz0XmRwIsD3WgR2fWpp7Dj2yzGXFHKGCP6rWq/
DZ9VYMdtqBkw+DRlwmfJALeSYiTr57V/qWupCrQNme0xUdssqePNBckSMBpPQygtqQ8eZPSkUY2O
q7VzTya83sX0S4R7Rvvzzt/oeTKG3uPhwGQIDkq2Qyf+u7S0Su1djsuOK+Zqs3jUz+ECCW6sRwGa
1OLHqMD5kGg+3T8x+TidYWveyi88aBqOefUfwWUkdqGsvwo6v+TiyD4ijfOtoWmd2Ro/IOsnBrAr
fpsv+xS4Zv8+vkT03MEIiqvXRAde9B5yq8atyl25niSS5+4rxmETq8ZtNMFqAUucRMiopZkWYVce
t3vngtQSt589Do80Bdozx+eiJfr6iXEZFEuBu1MG7UP6Uls6P0SjIf3G/ITKASpqKng2EhOTv0+x
zfVAO01kDv2wF/v3ygm1xISWvP34NeXMCNBlGEl9w+I6LNQBuyzzmLu9jkPdogTmRTZlBicE+qsr
KgWNVq7x1KBPUjeYQxOPkru66HnTKLStJzkaNwodO4fym6E+kuwNOcLpJiqWDMN+nQ3PL6CJbNXL
FIsgVr16mtwqTx2G9TqQaOlz28cK1RJbyKBHY5A9Ys5gLxhTSOY4kTJaHRe86/3IZMAK1/RAt1Jo
/hq45+NReBjyQ2/YWb61+/FUKM/KODsU5ov3MN4iSw2A532Dl1nJ1ye0BJ4qHlOjHRkL6OhMf97P
lsBhxTCvhWckiIhM5XgeZwoXG/9RtpHhKUvn9LEjBT3MQ8UKoKGzy/g0KFGwYWUB1SDDqTfPNZc+
3OLwy2LAXYmCmvD+4vQz3vGBdxkdjv7wJKsEgtoNtRBMqFMemt6smgL5wA4hqcr+GWBbvK/aqi8V
isLlDRpgz1GiLr4dr6xUzEo+IMhgrZk0O2rRMP4mdroDG6fUr4idmLPW81zHTkmakUCjK2xYeie0
B8QmFwVYuBubu4TD9QFQcQBXtz2odpZn+x+1b1SwagISt1BBVB1K/7G/kwmTYyjwkAuZDIhlQHv4
T30l8oDCJx5+55dqE7MF70vOVNrx8WsA8efNCmk9eFRh4RGWqsxcFQq6+Oe9NZaF5xFz3GSsEkR4
vOni3UC0x6LjEZD1A287dFFl2oSVwiMcuAyc0EupZ3VZENHytKOT5CCJLBYp4iVYewNEcq6/4cWQ
n+CZ7qt9YdYODeia4wktHbkA/R5Y+ovwmFoIuobsbEDVZ0Q+z2dFDql5AcSmfUDbhhQ2c0SczRuX
hATduhJaIIdUjJvGKCy00PuFIp5VC8B5GGXnaaQaEAG+iGyeqnn1EwUa6W+mb6BurCQz9fN//CGb
5/O0Tk2Bc0/cWP/mKRfUcnSd+x3pI4KbxTORiHpqy9JxlaQ0gImKZojpdgZa7iDLNsRlIIdQZ4Ds
CPPRGl+08A41u41OOAmmUkZIUea+qMLFjcqQkbFkS6h8qe7gM4i93fbBbJncDAcRLmEEcIWLN+kT
od6/I6CNuZVkHbGfJyUnclDjV3gMrzzut5qwnYKX/iemourRHWly5+PyCHz2rcwu4yaJy64Cm1xu
YXn/vISuQX7owb4SlUrQa9ARfQf3UMUVQ29LHiMbHpvOdnsaQzLN3QryLzU3bNsTP6QxNnKUEuOA
PGHUIiV57VOifEd9N2LLoL7hMgr3xj+RRXa6KoAXb+yPS3I1Lb8A7jY5kpvnL9ZEEYgkVQFX7539
b+g69GdFucREHK0dXvpm9gGw8Cbp/Gq3gVup0u+zEATP3nLC+CUSkyGUUCg0IYbhLTVJvt4LgmYo
K6UvpQ/+D83wr72GAJnh5bZBdJf5NmiCscUzQrTuAOER5sYilGCYqG7mXzhUatQz2bGt/yXeP0T9
H9pDl6hNBMnms1ypWvPQwASrMkH+DFYMRbyJQRjwye7loJfEs7Ge+PiioXEefBdU/ZCtqvW8aYSM
q0493xFs7FFizREZAPnitFHXc27TH+0sbVdwldGgD2t2Y/GhVHeahcbcgQG1DqKeCMePetVghOxO
mCiS/f7Kue3a2Jfo/+ir0UQrpcQDs7Bh+pJrfXI33ZwI1fX8T207uFlBn1UNU2BUC+tN9s6lTly4
3p/QeDbxrqHE1+7JdkGaeB6mRRSOMx2h365v8CsyGJ+m6lT8nRgkWJbr2cuFtkYkWFU9SHlgaXTq
eAGD1lQd6Btf2rqdyEHkU5r90z1ov2PH+DpbiVd9I0q2f40+1Yrygzxmu2Io8hk9652EVslBWVfa
C+WDo5U+3hOQvUe+kxyJWfKmIk/KcEqpcpTV0uu7adfFPvC77RkMWLwCUDj1sjtjgq4kA61FXm8s
V0ADAPjOaCkgWf+pAck+tyVjK+jr8o9tPo442VSTsOLowh4qwab3cTtT/h3EqJU5VOLpG2KhKBAE
bkpIakxYt9527Y4xSyL2rkWhjOKQ0C9uHFXO35x7923A1IBa3yNobSPIfqbErn8wA2oMO22fpngN
OPFmhfvfApLLueLSMNmp9xFPfkPurhKgWQsFtu4gD2h5LJSm+B9FuxIaasP79KJlz0bPI7CnaoR6
+3OV/WfhdOU+oqEuMXYU9Xaqp1jwO+yDaSVYIex3um7xAS9+Hi2X+aYPt4r+XVTOfaotG4nN04Tf
SxEt5DJq9LR6z4qDXFfQ+fanu1xeiW8YA5iXGtdPzPYCjTT3UBGFNXV6vHza3tP5y9krRu0dqCpI
ZDZADyYYS9AfRHok71qgBd2LWB0UO/pHVvVhsjnYJ6/JJErdnTcpK59M/ZKka1jCMVBTkHO9jiRO
odCtieXUs5vc4p3CH0CAsAPF799r8rk5HFapKIww9BQ/zXRwvu9khcioP1GqM672lyHoHniR8Sm8
tMmMR+J/Whe6giWyQr6owaOUyGQmjXDLG/a5RZr5mw1WSkhM2wrbu7cPS2USr3sshxlvZG/o13Jo
etWKMt6min9EYFHOvDHtZXj3Rc7vEmE5k3+gDzUCEhvvMd1Mli7SaqM+cvYvzv6P9i2+Zob50Z8K
F/nsF3HR+N9NcDf5FseibD7AAnxK6rxB8oLo/rtIG0RbP113q+K3/wH0Cozl1D/6bcnLksXvVJXn
FWnfz6etQiJIZ1eOutfvmTHn0VRltHJKV2wwg5beDIalNzPLH4LHBrmHaLk3cc8wV0yXRie2hyM7
bYS2tfqeqa1ZBsv+If9WK1ukC1ZzO0kUkMOF40rMhM7XyL9OcXFwvyLyeq0BUZIoYqLl7wqpKEe4
NiEazdNiDsN4ZdurCLuazQOqTMsDuuNJKetrgUdPC7UorqQ071VL+VrqD+vfmHY788Jfj1lFf2oH
mKKG3ipS/AQpcdh0fhOhJJAcqFQe9H9PLh7KNZycswxaILpSTprk9hEoIbdhu4QFFlSoI2cwMVbY
fTNg9rlEI65hJWu3+2RrjNp6Wl4ZiZVuIWdlkaXo2iiFKIBF4OyOtscvIeSNyqdgqnyQoE4UOQuX
iA4L+ScJNUpmDY2LeAgBZSlAkmr5G9sK1qaX5bdbB6ZcuFIDxEjxN+A1Dlpo6VrQzLFEElzNQj+S
tUTBGkamFJ2B6JyJDC2DYsAJQhlWLCEg9xiL0C/eNhjJ7HNkfYPOyQ6reOZwuTqBSUMr1b2LLkaQ
kJruuy8q+TaxZKJDERB562IEP1R1JxY2JjxmpLGt98QgBxYZGqCHeR71nzlW9BdbHb6dWry31Bi/
OLo5hZQdB1TdikVRYP7eOqGn7zqj2ivGs/53Y/0lkI2Fr3nv+aAlgWwm+rb956Ma/vyEKeL6cZCQ
EZaIpXIWAmghx+K5XdupQQfGm5gsf9PfTzNt62rA0wHRRGs1+RLgIvvmPLBJ8adq5KDibnQPu5EL
yGfGTcNEdwwvSat9knoF8v1mv1+sTB0Bze/p6YlZvGEGFAe9ncjyuUZSMv30tJJM3QNX8TFi6jwP
166Ii2LZFPS2IbYV0v63APj5TKSrCqPpWiMYNyNfpEEpSu3GOoW0IXMjWqIIMu58xmcMuF4Y+06g
Kqkug4I1GN+Ov3N4BlRne+gBM5UgURX9np8LmPkOwtVw/LICc2QKsS2mVc60HLfKUBp0d3tMC8t+
/Pa/JgSh4o7iAbza+G0NiSsObz+HYJKLsqEcTOh9CXby9nAczpv/M9GZOTvoTBGeBOevaN2mZ/48
rTqCkUhXo9Mhn/POmI8f3r1rjtcAHQZLQMQhYgyIQvwLiXknZVQMnUJ3pP5U7ulLrVZMs8MFfmSG
BHoUw2VZHa24XtYNKbE1FX1tH+MCDY6ONtaRvKgKcqJI37H3LY+qW3gtTYw/eFKQeB+5z/WR/mfz
vqxAd4AouoYjVMFkHda59twA6O0EyKntXf0PQBuNRYf3F4v2nmJyrOzuDZpseVr6fGNuKh3Xapd3
52QTitLsGR6cw5D78TlcuZQwtSzsSETC4iqqa2N/ISicgLmdbrOEvVVEC5jZL1dwKM3M4e1JY4u9
qEqnUeYBQ+CnifjJE3qp6s3kjyD0393BDOCCKegBpJ8QPZdj3QLZSLFs3tLAt7dufgWs0a9F89a1
lolVfu08ohz0FK5rxy7U2QDJf4czOtYGNdzgcpEzetklbAujFqjaG2ocV9q/M1JbYyrVsXKtVAOq
/w1sUvDEHbhWpIZxKoBj6lB40AjoN5ESUnHSRG4a80ZxNhtYz4BC35uGIndGaSezr2ZJ88zQUmoj
frLeBUedKMJdzR46NsOUX0l1NM7iBt09GzkrguZFl3ze0Uy/MU0e3hXgVuOYmXKcXeZjRpfwvFbt
vEgmlXBT5o99ngf94tP+170rdo7+HpW6eNbf8dpzhstYF/LEu2ttGEsA0EJXWiRLgRnzIJbY1fjj
XBgU8+OIMJptkrZN0konyNZEvn+p5QdYzwAU3HUNkz2FcfXGl5Sps0LtMbkltEWyTfsMPOQ9Q+o5
o1gBgpYXtnVkgPf9n5Lh4tRu2DmfNOqN1ipF7M6joTrRv1q+mYPlHnhH8zQeZC9rdizFplb9z1x+
dYQTG3aq5a9rJBlIMrCpBQFvzfym2PV2lU8VZ45TEi/cJU3YtcwziUHLofNGN/NeFzA7fUI4m19w
XuWOnZOZ+ykg5lpw5Az+FR7nsbr/zcE1m8rtgzrSFipHx+X5JB/IiQyhT5W5hv60n/Wquqo8X6tT
El0EX4VhrjkC2NtpGxf8gdZRtHTnxwXV0FxezchV5IiAhFG7V2zBopkQNXJoBSUeFTUj/kMLE6Gt
TWEOglxOyuKRqwGp9sxUjtyrdWz955DuxyCKmNu8mS0TZjAcFN7QIhj+/WSquWCsbrg1H1LBRImP
Daxgkt7mDGXttjdvdIc4oKmTi9m7F3l/T+KTohB2Hu8VWFC3INKESTcmL1/zhF4sRQ/Aomn9/nzO
EGR4VimVvAJJ9Iq4a32LReb2isPt0NJhU3qWRDKQumBlUzjf0D0jQp9NP7lALibRiDJSvb3muurk
IYzxfLANt4Scb6dKzYb+6oEWKT8wD4JkhaHBhNaJ/6wqbSZo9iTWFXEVJtwkI5D4nr2w/LfXs6JW
9lqi3aliyDmdTBSyj5YkhgxD97ZcloGgTSHQ3T7fQlsXacb3/JhB8meQdQG3XaEvJw+sKbgiflB7
jQG69pBX82L/1CrmiuEq46Xbk2hPMS9wrUjnGBRwagrEImV7scyepU5U9vU/T8EfyPn22cYCC2R0
pNULHJshvg7TN8oVPpSntZyftxoC9rGj3QZEZbLrznxDPtkUt1MLJyzM5pXMm6SbeTegD/JVKE16
nmaPIi7EfyXnjLy+C6/A5kEQBNVgU1bAuAEcoZES2WqDp7fZ1HGUfN00WNhBB0j5WmqhqWamILWh
EfSzRB4mz3DPuKoGAuqxhnwja9VhiMvBzZ2dVLv1t0JOodiIuiWGSeuSWNR8PnUwOhN+rMWW6AGI
gObb64yM428+cUYb1zIScP9QU1TqP9q/pNrKrj/sdSZscoBzfc1ltuHQjsZb2GDq/cJhTmcVSyD4
E1C2oBdZ3TtJEdeG9bWA5yabtbSDDy+LtKj2yKtiK6hvjxWE2kK9u5fEHlNaa7/H/EsNPPO6N2RI
d8BEPvr259lx7oe+gmAeT14KHmOR6pRDY9XMuqYTPP7Sx3Gtlf3ng4soDWABa4p2E6aEH8nWoY+m
OtrzCuX9vFp/0CwQFfjLOcv9KiTWjO4q/x27Ml2i+bP2hxXzfK6s6/CTSFAhMSvms3wGGvvpddgr
ZdPHus0MGF5nvFjRuzdFhsrm0twHmt/4VHNhSPpciw7vTDA0tWL7Wc+TVqNm0rDkfW4+L+I+lWpA
uM2NRli8Uik75nERqcFZUB1PqwqZ7T54B0VA6JECkverl0xUwGhZowwImBVfAuBp1Qgm3cLKKeJh
bOu139rl3WRqtC5SrO0qEvu96BOUzdzTBFaszugx0EFwj6VXcadTxJWpE3I3zJRBIyaVgQrBwEUV
N9tfaZrsFxy6DgfX2kkb66OfdTjMZVp1FfPKZ3dMgwvSM0qSG807CPmvrdinfEnSw1gJnjB8kLo1
lSzeTxN5C/J5PJP+Nf2G6h5KTFrfPvEy5UpGZwV/YAuGSoLxwLFMNaGtxRJ03Jty8CVAUuNsSjuU
BtL5tAvLDPhoasHXHmXkqjY9KPltPCrZM3VW+jA6Y2WozEFBdzc6aQVuDgdypc6393lfPy9lxmve
KdjIQrUcAQfQwpbGq8dXnT5Svd1Criucw3/WNCEfeMKeAuhIsb4qvYdGA2U26ooTKi7bSA0F9gw3
vNPzDcL3FoClEV2Ib9G/ztgdCFgtxo/wNSmDC3DdUxSgjghSKnrHljKKWfxj5oLw0M1yEDOGTRoh
KoYGy7fjUzNq4GM+SEBNEztYQYt/01RqpJj1YLI+/2OIQKAji/tGORSMjr5qXOAxpGcFJplt8CDC
ZhikyjxXLRaQjkxrAO69vEem8iOjbCcyPXxIfB3MllHtfEOdZk+mTR87tBFBnsUKdfr0r7yJX96d
9mJvEvpsGgJcJeBjG0bGIgXpnVDyESUzxVMqIoALSVqLbQ1ZrPNViLCVdKMJMyR+W+0EzI43QD/a
4nzGz8zNWVuHUIBE7t6l4i4o09y65JX3ZeZANi7WaGTTf2T+OHJZDJralCOG3uL9pBAmG8v09RRN
JI9Jdft+nHk+z+6tgIFBFMrGVzPbrxvGHSwE90eArX4cDo7ce8G8dok4JiB4yiyAG0+eKL5Q6m+k
aYW0lg76DIR7xXPPuCkCsUnYA7FiCl0s7qWmjKqjtYeUdsZAngxw5MTuvYJ4T+G0zmLpMjHoJ04O
268xNyg/tZG08tUNEaLJOSrfyoEw4LQtO8XoOja52znJ55OqE/QYdYi+tC5MGvwnwjXHZJEv/bwe
SZjSORcjQcTVuvK6zEWFDxrPDetgK/uGGKBZlWmKkXiGoITw5WETHTkcuXGmxCApQOSOsOgX92+q
zGp8jrLEU65QKzcw05Un02Mf+51j4Tjb5769pO9Bs3DcULTEnhETfjBOoSN2yZ9WdZVH23E9Ej2b
WXYSjxOmHCsaYTbDfzx+nHL6rvGpmTCZ0Z5c8Uvasl9UurcY90DT55fUfvIsmgxvWF086NJZ1luX
lmGuyvuLUXn+N2e3jujpIfpOPKUlx0JLEM4MHn8B/PRTBNNYkfp6ciIwHQ+XVfLMF/gK7+Iffnca
dkSO6l2gc62ENABUWX6rRrEv5OFyCOSiPwS62KimLFagsVsctMdnWR74UrPE9kMFj2o5vkRAh9Ta
8nmTTepZJ1wN7e3M0EsS+ox1cnLap6pXcyp8ewCPGHGX3H//52i7QNKgpqBNrA8et9hhNRPshjXr
mL++oJOdTpIjnxS8+dJd08xJdSpD0efSFsDRTmhgbCde85/S2SZXYzPwO4IvEJIdJHxOqfypurSj
oP3/B4cFnqG5KxTynCqugEr4CmME2H8ksWwO+5ZtSkRAMJr9CbQ8ScMl0X8YzzrRrDHo7BoEYruj
n9kS+VdS+o16YJgUGSGpOHCPf82bTs9zHPDfMyirlY9tngYO0mzhL8GkXvjnc5ZkolRNx3HEpBqf
oaloyFJ9qZdNy1nm49K8MtqkUcSsEnZGTNQ4NPRj09cdXsEqwa0+WlWSa13BMzaI63Z36BfG4dVF
DVGvXdOlyvJf3y/YIYQThC5vyvAMB8xkRkWeHCLyNas3LmRrRgG96e8sLSPYT/pxyVrOa9uzY+q2
PwKYtNRyw2jxnqSSbzcAq8e0aaD9oRdSkADTWdALh7fhzGk17o+WmhZzBlJTGw9JlOtmejTk8Owe
rNNzLh9GiwPJWGamxPBBr/UlL5IjCRz63Ptv3qTYNT0N0wBGDlF3ky7qpkw6refqErb4oS1U5F8W
ZYaGUndiv7BjWUIje5HKvp9DZofiH7BdaSV85CnDN28x5pVn3nC6BwA6o6MmZIK6HOV8z15Vvw/N
iR/mBq9NxnmNon9wYcFs76QR23JJz1J86PGzTjkTOO3POeRbqq+f2xZSCy/uVPG2kOQRJ/iIFukg
50LOMVrYXnoO2ZUMgW6iJkOrjXhke18wrXjGiJ0igD6I6gkrMaD9r9z0GswrUgq+/dspgqRJWft/
70+y7Vfra3xEECOktJWlYqQKdwwG5/dcsLkf0Wc7Pr+MdWsRaSMa+O97tYNwZAHK3TJv3+f0RLmT
U/wD5Gfum5YmzNem3Um+9XLKScqWIySBvv1+8n1e4584uCNipksqdfON56FT0O/eAP/2UYZAr0FJ
LV5Ve9ZJh+NyLvg39PHQfphpTMBJ67HBjdUMZAPzTcqTTxjiFFAOVKGqmt1cY7ujdHtXWmfBbeya
UiEfVHySG2vw3jetzHLytHuSMJQrVQV83dBoUFwbo8G8uBdR8JfeLKt7BO6NmaFes9mOzOgk59OL
YoWCOHnn8TuHIQt5TeEB++9dDpm2mGenJejeJ9jXlyODHeOBqi7insXe+aFlLjnmkrOfHPFVFbS6
i01ii3sBBmdNNzkkm4dWvhclkL8Se9i0LGeH3JqG0kFOvr4tinnwMxQUO4l5Sqv86GZGuvlmT6ct
ixqQkZGxzcvwSJn0d5J5kvgslnXhA5vAsDkzQEN0KOqSyUNxKKEt8UbGHuCJkVd5Xx4UU+paQfeR
P983DuGE5VfsDsnJ7pmRoCBthvFobEN1VHW+r24EJHHVqauSfIk2rvbk1GPywjgPeo7LyoXkV18S
zYEvozTjpAsCkhmwCjmA1HVm7E60wf+hnTt7nDCqTbwV9u2kYDPvVf+tAUKxoi1P08sKgayXt4R2
Bpykl+fYMjVhG84jzQmz7onQ9JdhEb/cU/UR5WuwDxmG/zyrAG2hkWytRkEix1aGF9wCfEp+Pa67
oGsScErf3zW0jV78QixT7u2h4uCA/nOxGr1vGi399thKO93z3joYJIBfXnrFq4RqhQHLeqPf5uaR
7dVNbqRxxhzaulY1JUs9kiji67+Vi+hUxwlpmfivWSKNu9tVhilI0Gbn6NJQt6/4fVAHIy+bbKHh
tOm+ouWIJKxuH0oM+wL3GSXGr0wYU6HvVTfSHfJ9Bw6YdTpX1AuO1YtYt/BBhNvOagU/+MKq1+GH
IC5nBnnqK8Ct+3h41HUE1KK67gTJeDspmYGL1ueIa3C/UYfGIfneoNnObHDAqxpV49/9Z8J9OfBT
ye/WHvnqWAdIhQgw2NkZK+C2Azan8RMedq7M0rEg11x9trIoA63rp0uaqXIPm9f3hHinl/DIS4f9
LxRe29AQg9y5gw1Nf93kt7y19ENMARGLGT5n7FhaQyLKDpapc6TD3aiExV8cnVldN4TKpXx0G6oC
o8Fz3qaqjKqF5RMoicHzIrPHluwxzZJESDT1FI52PAqEpaxWxBfrFKOCnkeWh7TPJFOLPgK9p+HU
GvA6voqreaMx+SoxOiadv4gF1VG6ZMFPn/21+PE06RwxVv93N8Ib6sBQbXl7DnVoT54Kt7Atuauv
NGbPxrXGEKQZ7kGQGk53pbftil7a9vLoQMuaRxQ9k0ijOOY2Pv9B6orCYTu3dsML0F6MP3nQ+Jeh
Vc9BLvvFT1smEfHP+sctvaU5d3IL6w2cnYVc1PjPmP5JxhmyinpnmLP15imB73H07tta62A6s9aK
8u48SS1zsloiEZeEJZ6PxQjshbqAumWLiC4DYH67cZBAtKtGS/XJhha2Y39z5iDMsKxNbdypr80F
vHR93MfuEfP9G8N5opwPmITY1Qz8KPrpM6TAA24biovQta68ZAWQDQxepe1/XG1HzLKCx+NW57UF
Bz9IvM6j+YEJGkURWB6Tsa/8IaSuLFAaunlA6P1wkiigprnS34gt2gypzkLB36LYDR/B2ljq5d7g
+73aoVJbCb6vHL1F5l4ZzGu5FSyopYfVWzkzQGf71hMElLz8WyD66K4r89X85RkXalXrbZhIuosc
dsFNMt3rDKUOsOBh9h4b6UBzNTUCdb6wSQ6CEPiD33a2P3JcM7vChUF8CngBsjSruZKZRwe7ipK/
DDVRMyL4bUdV3kSFYjPQGHQl1bdRvY1lWen7qBGhHDIxuD5OdhM21A9xHdsYP+pu33zxFD2TeAI9
SOzPFo55rPINBmv0ECpnoTCOKQI8ZscCwheJabK1RqTDqy04fmYhpsxqvQRsuyHzoUOGuj6FByH/
7EOFkVQ6QkXjgAx5ZGD5L+MopRhGisDO7hMlPI1nkfsB80TIjqluD7SCfXw+YIKaTiDBeM8Sb7q5
jde2oTMADgXdtXBVLjkzTrZuBwHp8LJVwOcnekE7Sqw8c3zyopxJ68Bza+GLphob9m5A9uxnE/Xc
xPUjC5ulv10EfXriOIZo8dAMlBvRQy0icq6r7SOjMQiYVYYjnfb0yMWAM5RbGssBO3IaC7FHGBkX
0MwNfrEtr0CugFDQmi8Be/U2cJjJR3JfbfZuV71qIOZe4VUlEhNy3BqTsClKuila6cmRTaSqPKh9
P8YRIG1ALEAPJGhJx5QeA/Ul4OKlnajna8qhFGtlqJlOJqrH9MviOqXCbsCn4lucGDzOAE9Y3tDX
GvRRAzFs67DisP5weXz9tbwTCXp6YGRTHML0l1+i7GvkyS6PIzZiqV3iPReMdWQvYf/cphbyQV3B
EjdPVkr4h5kXQD4gdQwK6FNrLOVmbqzoycuaAsb4E2lmKQwT8wyWbVU0z79ZuG7b3O+fGKW9KqWs
OdYwzzFZZEyWBAeK/Ci0mVKBaRRQl06BGBrIfnPej1vmpzs6JSicr1FotLwoH0YX2NhrMb/aIVyk
oyzn3Vwtm8JCZ/a3Yx086MsbSUsptm1Xy108MdfxUjId0aaPAAETNGCCOOp1L6UgdA528HWLT9Mi
2rlS0rV5mJVGdq8qnuLJbAMAfDoZJ0YfnUs/2rOwOGFqnprF5FMOgpU9NaEotiZ+uB1E9KEnGdFo
RMTwLWXt4XqM+1nvdu9ZbOxR7fYShc/8gH0TP9m6b9F4ZOm1nyDlBjOkqAFIG36dpChfREDzBALL
brtWQuibfqWJ1/uPYoSLEe5rtp0E9q52Pj/gP46AJagczpAeQohKAda4FRfcn5u3BZB0bTX8of8C
sLuKAGhpbHGIAAdd2lgkQoV3JMgHG04lejcRCMj83hQsuKZyvzvlvdCp5jiTXhylRdEwP6VoTUdJ
XxsKpSRCzZHTIehpj3FFtP1EPb9NgXCbLz5OgGNlDxTPJodN1qflAYNmXIwIO1dQ2D8HTf2jaMcD
Tr0jGRC7S8X1jJNQGBI3plLTwMiHaJt4aTiIZBPdx5L4zzdc2V9y3CgatlJDXzp2JVBCQFtWTB4Y
AdjSEpOj+S7lsCV+KmxxiPK3+NEiyVo3GAvmtMoJlcEquWmKSD+NWlZZck/5JUPrBWTCsych/IY4
rEr6GTzccPELakKWdBnXx+LjGRXkf1JUKKNSiBlpr1Rgj3iI04s+cY5I7Dl0alJcKG1+UvKIS7Ac
dXO3u7c+/lGSNWaO/1vV7z6zrOKJnxyaL7Cgl0SjXWd/MHqygJjAXAdJWVa/tTt4gRmQbq7tOTtw
/BebkKO4rOsKh62xKM/4uVA7KtblaBD4qeLvEwgh0hVdqaWDUmwfmje+1h32TMhfm+i2zWQquYCH
0uldQfuGiV2PZYzEKx10i2Oy6KKowsNw1iZp6ANivk+xxOmzUZ/QRVzJHLjPADp3bpujaV2k89bQ
BzZ+OiGsCnYygAxphbCuyfyweIS7IDYNItR+vjL9GpJuabgBt+bJsA5oXahrE2W0ecrsZEWcojrq
5djkpCOoa/dx48hcfv/qo6MPskfmxRyTiZP8YsJvk47hXkAMD+C0GbEOVzjKCmhBeYjSLQcmOiBv
t41QyKeViCBYnhoC6RokeI/QPwqfbRoH3yg8Cxn1AQob6RmN+us8fn/Uji8G/pRVyo+/OZ79BFN+
igCxLFWgmYtCuiBfyet+6P1A23XJtg4IbXauqbD+94K+nj0ejyLHUbT29AisKvbDf3dFcGSniEFh
p7ym2ZHkrfzPnGfWx3A4z7QDO26uOTDqyeeIFOvLhBtNNk019WOhYNEFHIsm0cWeb99gY9eFbNph
/ScbY874gYJ7XSwIFkx343VRl5OhJzijMHbnhBhmfV34cI0m43X5OQAzdfOVyKdo8fMckIyYLp3C
1aG/XA/0uDFr405eLW1j9AcUvTTUILN3iKW7IAkhiPekZe2hkA9HTDM4GQkmBPUK3U3ayF9xrlQf
a8ZsI1RnBYCJ+MjRvrHFQhQuAZkUfsxIi9PiHuU1qq5OwNwM0U/4CNEN9OpsW/mh+wLFQSYQTHVk
bUCuZQwRdBQy6VP6TDDg6lHccC8n61e2OqtSPGLUD/QrOTfCKPourQizB83qVj3xhLC6SGd8dTJ4
7azqVU7smFjO/ulrtVVFPWLA2Om/nPHmYkwg9kEOBuSx50ZrToOe2/x58OysZVgQG4rYBTWY4yV+
xxSnhRmogNZd0TznwRJiKLM84Xi7brl1P0+45HlU8hTZlQ/3v0uI1AwSdye9f3QfAPKtSNROmY0e
LW6WhOlAg5fRF0FaD/lvCxVGRxXL4NJm/TGXmEUBHD+uaoWBpqp2MX3Jmqwc+VY/x1qymeOcBz7R
itw0cy5arxJgJUbC3O4MrIj/W4s04PPhO2de4UCj9+CEiErwZp5+RW7ScaInbWtFkKQ3lnZJqPdY
WvKb4AlX/swMa5sHJ4rbwwV2PkCpjnSmNPPYyMrDCEpRC6jmpWRdfEt/QZTfLvPFaEoHhmIUrPAq
E7Q7OtCtb70SwKsACf9jPMUeydW5xSg9+fancL7wUyV3zpIIbnLYQ8ewSercQr1YLeV3sSnBz2QC
scaw1bpJqEjxrafxjQTaKxrI3kiosa4N/zOPmXy8Fi5OcGG6SFAsjA6e3SPTvG4tX6MFM9zGirh4
YzPXJNBmisPD9Zwu3UKxYltzyKxxbiGYvfef0XXajetbVrvu0xDfGGLPnf3AoRvF9QXrsfYlIvUZ
Elh2BYiIN/TJzCkSUfK1AvxEpiCx0vmq8/NFpNCGbXPqiE+NfulQqUuogHhVbPymD2M7i5RvBGaU
0dJ7o0ztOCYY5Lc1QUcxR7yc0sYxyxmrwBm8OHm9XnW0AVMlwE6TUeOEG3UQ9tHQWf/LQaXXAtua
e5z47HkjzXz7hbp3UBddnAPSPucOByE5SigacwOWL8ajizTNmfzPf9Cf5IY2hSLXvEt5OzHXuu7W
zvQrYgYnNlm7KN4NlJKe5kLtC1clx+x0eycATivAu7eJBNJ7xd8MvvKVQfwjXdjP3vWr/fJPSZ4L
BwP+MLc/SkuuWgDJJ71s01ucWZdTzkdNHP/cCaOHKZ+JqLuNdZDYHROI+wYS358v3/M1poSPgZXE
w26XFr+mB9MIu6/NxReChrNHtUo0/1SXP36d5wIDrByCf3NY69LWhSqXirpnpENPOmn9m5JZM3ZJ
ejKBb/dx7c+8BxPeBDKZA+IsAjJPbmEUFUPK/lyCpDuYbpkszIvBEpuNQGeiGq0wQvszm4oEk45l
dNbRPuRYVMUxZc094MhfYJ7uy1loA75LtENsnKjgvnXTsa2aYd334O0T0MQzh0rfIOwcd4wXlg4t
3EIy9xBkLtCyBBqh8AQ3Zg+/Hm1cPZ3VmWDn5wDN0PkBYvwhXKGwZbkF1BDYl8GqXMWtFRIa2V0M
VaeV69YSscUBIq0prXqJ2MWLSVcr/bHJOXNNHzW4DO4S4stbW6NwVcDVSCeaS1jlDb62yclLRDXs
NeTBzDZs9MO2h+0v0PjuDuc64VQ6WziwkG4Mxcok4lrmPaTs/xPjZV9u9TNxH+YZGPVSQ5LoWIfV
HlcRSe9yuOE1ybMvKnERDdrxGweTig8OtAcWhKtlvYvv1l4h1XQsWNay4MMX3N2BQT1t/u8aZRmx
7XlVq00wvh7qYpsOTwpHHZK2yn02y3O8/57xyhDMWGTPswXRqvMhqxin1FoKe/UwnIhtzLlrFaY/
0xgx8Cpm0VXCc2PDsBNE88kgtzWvZXKJG/eeEtJszDhZTC8naGE6pot5wGmpzU4YgzG1Pt/zp8ti
OpJqvoUvzVG3cI5iBEme3v0nenh+0BQsmd5LPHgA8/F++wCvsz3TSHLrg2YXlofMqD++4miNnXif
XwhficnzvgJ+ANDVncVNJ0wvc3hBbz+nUVFbyvC3fzHLyDvN7PeSqSzp+bGDBxWXSDJs32ScBq9a
I1vFEeypNy3N6uOB3slk7oRjm8bzirREH0gU4taBLAzNRL2tUtNLE1ukO4BNwGNNnoZLZYk6bfi1
x1J9qkrQgYcd0nEu/rkgCbzZm8hpa2/vRZOrnVE3104cJoF0hNxlj0FZrKmV77Kqq9aE/9Ht0Q1l
kGseD2omLJs5NuvXJFwNl/kFHBv2L+2ifWtZCm+wMpVdDCNCRHgnFPUoEOQqFGwNNn42R6hCmd6u
PYqGdVCw5u02wIgchLEGeiU0BX/7wTNmfKbsghAQEt928uQ0hNRhCWktlkYjHprytEtVJUEF+zOQ
lL0WT0ZtPL4piozxfhj2m6B8U14HrdLm3fBef0v4GKbT8UzETS36WQNu5YyqgbUSfgpimdbTiOVt
TeaRM1DG3KzF/YewK/msscZgiZjIhkl+u5Q4kUmRHta8d/fGMHqxL7+CC/YimPqIdW5o3qiC32gs
+O7v8Nekb14p/wzohYrXjHE2qxGSVYc4FtlNSmjZGN1rgC2i3qpgsnX/NlzwXkQur27awG6OeVmM
3nCfygt+tEg4rYsa01zE8+GWgUrATEZA5p0p5eTk6UOeExqD8WPf+uAceCpm2rgqpA+GvrOYsO+q
MAY9xXgD7vevXn0Wq1qvSH3UfDYNPLM1+LuHssLIg66fYdowJhBXkAxBvvWwi1j+3aflXhb9BsEU
KqSy5r+odG6tYrb9fyOM4Cgm45+2VeZWxVF48e4VkCoHnB2bj35CGUfthd6K1MxTLTLdeCktNg8O
Ib1ObTOKH1230DhuSvSsauqCTPDZAkRwtznzIfe/Ozt4/sI49vPsc0WGaAXwyCCrCKwxz7xhvFrg
QXp4CwuhlrVrQun8dgq0tWVYFwlu9we7sk1FtQHMIb63mPBsTeqdyBDWZjgqJx+aHJ3vXSUfPcAB
37FMWcxWQuY/GaH2XP5o68+kgBzM1xyRiX/TFEPolSdFwY0Fh8f86zoMRWpfSdQk6OHRuYkqkw5g
N2tbJk7GiT4WHImyOCleZjCy1vdDO0vDNwVBLlDAr7hGtF/um4XsLVW38zMlOkyAHAXIJ04fhZkq
2GKuh+ZtyqI97aTP7k+77rIFm4SX3Xil/UC34dduyYn5U1OFcz3J+7xT1yMVd6k1EfzRHwBXPwPC
Urr7vIbvbQUY2U4zoZ6WdMUx6nCNcGP+NIpMFuFfEVdGgty5XPmWIVXlO7oB1C4RsFPGoIqJtEgN
Uwd3GlMnGZ+dm+BW7+DUEmm5WNrfCheDZdJV8A2f0gQsPYtmEgoIgtpts34Tx/3NqcvBpGKBhl10
R9Ogsnk2Oupn8erU6pzhMTKn30o9j6DRQ0yu6BAsDEcDFjJRFf5FguqCATVaQ0GVAsQCCtC3meXS
7o4yANpJkVVETGf5g8QyA9Zg8JQSk9qjSdVYyLrfr47tJcw+4Cdty8OK/EsIbvINxARc40bVV7GP
BQWXd5+UOtjpgeWRcrYE9AbAPZloZGgnuw3xcAq0FPJN18Bh7MQdUdX6dbGMsUNokCSLzP//Nlpu
hEbTBWubAX+dk8ZzqXtbTaZgMgxiaJVupixRF0geJUjHKDeR9nefGNgx+d57u5A0qaIGdc90HhDc
nzKcoaudN6G/3nnja/svEgbdyh+AauoNtITblE1yeGN7wIkgNQD/S7PGOut1BqyUWvAm0MtFAByo
uumz5qgyWhcL8rPLBzWxojuRskTKxzRBA5MZBva7Y4aQ/TlmqqovOTaj70ETTgfr9nrOsXV6tgBf
AKW6Y/bgpP6PoMIvIqTmA4Xgfu8jBVubQD0JM3Zo9czNP4lISZK/80Lhi/8X2r3PYbhrp+LzW+20
pPe2+3jF4FTGkxwf6HM/CZTq9+3rLpfwL3EgdtTErs0nRWMHQCe+vANuCQZRlkeJjJYB2e0A6Zmp
DDmXF+dAqJrQGjCzWHHaHBh13FlDCoh+acpzoWCncF3kG0bDp8unuZEmkvQDX3v1Asu9dSxQEGT1
Vz7/HKHkiuRfm6iYStzh0gtu2JJKk4DvjxKJlDlF67e0KPZQYqDAbDwxP+cPdS/Sej0on/XUSPlz
BGzOFHPLeZ6kf/S1pnitLzr3wCsAYxd19VY82GJFrXuBO9dlHH7XLRTLgRA5dtXQLK6g8RHkm1t9
7DlJ9jf7iGMVJEw4f+3wskddfoVvRtJwMVOAQGwEG3VLJcYOKjIAvyS3vJBIBoN1ZcmVb32oCLG6
f5tOSOYXcIVPCpS5QaCrFg7eJ+ZsPN0n4XiNZ8DRJX0UyQet70vPQP0Vx77d2iXwtV7aEY0n1GwI
T7HApvAL8uhH037Qh7X6MzaIzMGg/W4cE1WlhdM2UVhLLdJyH0Corq+/aV8vzACqdf9YgB7aYagH
Et+BxwLwo8kx7Hk8f+QdHdGnZkRuFqsdJlPxTtGLXTMjUi08Ihu85UrsgbaVTt0tOX9hrxY3kIO3
0DV5jffZlcZB2/ZDdvP1eeQoS6Kcs0Ut+8zIt/niZYS1y7C5zXjlqEFjxUrmxWzYcTSw/z0kxgdX
PWcUW+hsqtcEWxjzUneu1335wwktEV2xJh9vOsMIXqtPCM/6H0q7cGRVvsRmh6DI8GOX6X685sBY
8EN0tvlGgmgETTxloMnc5GQj6gw0YvK5JMJ2Dl+Cq/TlfSnOfKt/OfucUavKWbDIXB4o8JuxhG7h
v/4LAK95+cU3BQk06KNKbYoDpGZo27r+ECoxNm0FP+/kCY7pnFF7SWx0drQX5LmANSl123up7hcw
CVkeE757/c33mJcEy9sj0qflCgtlWElqm7eNqz3pZFiGhNaFdR4bcPt1bS8ANRQcp0y8lwmhpvRL
ecsGVEUKuG6nRDfvgyKwA7oTCLTUTSSUYAtZZ2jLm7BDavWHjMCDzQsIevE3dXlfCZAr/w7VySjK
oHJEkPFPB4/+pREInYK3bQMEHTWt8Caz/va413eXUv1W8PQdZ1YaSMh3R81NM6oi+C4lOdc7R567
ioFZHgC+U6LTE0o8cHozEdlJNhqjVGj2kSfH+T3hBrlTJ9MtNRvrsoXm036OAz82N007Ep3srnRs
1JHUcIeZh5Z4tMHMIQU3YQf8FUKo9ypKT+EmbH7UmiJRxKhAQDTJ0A10jXohkvP3NBuTPTMmhp6J
a/oxnCKkgwS8gGq2vbgnap6inaTxkRb6deJxV8NQXI8Tu1l/5oPOXBqAREJBlkkL8olTABtvsxIL
nsZj45eNs4GugR73TKwRaBoUzZupSQiZETxLgHk16elbOHWwkkfI4MPLLpo0vhcs8nPx8yJ8jssY
A54mAnE1Q5Sy8LWijJ3sOWbB2Vgb8BBOU+po/5gAD+4mWJ93/zAPa/0qF+AN5Gnj6oVjDY8x2MUZ
j1HoUqCh0JyfTh0pxyjwDUbgPzZ+vd6irX+ntj2R1qiF/ZHesQwoeuwYwsAaGscJNnWlG63JvLJH
IdZGczCug0Q7v7iu/d0dBvkVfbm2ziXMumB8s6hBOAYV6Pk/qa3xJiIVjtS5cNqoc80SSn6H9cO4
xj6HtgaU4of5PtA+xvXl6yJe40IajtD3Eg1/vQ4kSTlbtpfJxJXoBor0q0BuhMYpuJjzJRu0E8R5
gRg4UG8oxAJbvmKotoE0OAT6BzAnma+xpJNorjLiD5k4KXz/qC6+mjEEzGQkcOwDCQR+Qk+Jl+RQ
VBR+v6z6vAYpypyjsOlOVOLnRHtche9hjx2nrGjgO0DgH75vgKafVZ0UphyKDfzBJmWjnc4ACb9c
beY31MeQiKVuGQGga4HrXa9AlVrXhmp8AFFsDAg/DO0jDTahV1VZ7mQ6bze+Sn7WMT1I+Denjz2O
MQ1dVt7kCbEY27krKW1A3YjOzvq7VI2N3iZIVKYKNVRn/5g6Qdcp7giydWG2BuyrWnNkGVMzBg9E
4gcy4rZILGy+x55vaWmS4Rpv0LcwNKYEIjwreBKSEznqskZVuhCsKU4QXFt/P2xhRe2rKgdCUCvV
QLWFoZM9PcMe8+RaCO7b7+gzPJ/QGYwdCmg+s2FIRiHyy3q3hq4zvgu9dalrdMwL0O4VhWHXaFhb
co9JKaBonyhRB/YhPvJNDRAW2a3DB5RL65PErz++kXMBx1/hCbBLaK3D0/6yvnSq60vc4PCzhB4R
FYJjf0rP8adJCX82wym92EXvpDUGtm4ds83SQqMvMlThEVQG61kxQ3P2+FIRmo6FrCOSl0Oh48iw
zK24Ug4Z9j5hzCs2GEjn2HMB3SflIEVTFD9AmmrTe6IYZXKH8blG2tLZs0GnzDaGXMaZEsFtDk3h
Sf5I27MabUpqlELZbPDbpsfLZ5t/+znJ3o29Gm8+cU1M2OC2RrEnWUYYA+0Za4wLyzxGT7ypB7Xk
khYI4iquaHGFJQd7I2zCenxhVpFpL9hRz8ZNPpzNGup0LVBlvgJUtOSw8Fq99GNYJeRfkX9CQJmp
uwSkMjlWTtOT8R6hsifimp0Zy3A/6DyMqjt6jAfFUzyR+pto1/Ps+RkZbKaXieKDwrp7/uCNgM4c
QGBcEN9utuGXGtmeoy2Zd7Box92N/NXACiUYM9QtlzAmPgwXoCvXKV2836k0VwDosuRrBJGT0oT1
tlCb7MsYEM9psvjCRXlxs3LsjOfue9obA15V2TA2LcND/0p7A6mpPLD0Fh0ytBsBI34B6HAJmMH9
Y842lKMnAb4pQGbKQaGqnRewBDvpu9d+OpIkw8WAChTzWhlv5LjblUFvouPrI6xUcRlOFz5IMdlp
H30xq0yLspOWXyelnx7Ofll5jAJcYIaY9HvfcNMSuAlaUmzIoc2moThuXDSt0/9vYo6FyVoH5x0U
Puwq36eAXIh+55JhynpFsfwliAkryY339OQcotMbxn7241YljLxscWfpF9zLCi0xR31sjmDX5nqf
mlrJE/Fb2Jmibn4euRenyBX9vzHMISXe015jC/DFb5dAnuAR8RixREmiP7emXoS/o2F/0lJyFgnm
Tid2w6ZWsm8YFLOvRmdgCbMXBxMjx9Ee2VF53fFZMTT50baRF7gZLGKt4PqSKaFNYtK2rrjtSnk5
YWxUzJoFwG8M5JhzPBQ05jfjigSBVoG1DAKIjuQ/rGk90GNLEY9s6AmN/7/7gd0nCtv7BM3q3vR/
6af0mQgRrMYxIN1KiQwhwQI0Q0SGFtilmGaAANLEb3LcfQpG+hhPHbzsH+9BI1eHM+p5RXsxR+zY
m/UVQdYbimGcuVRRuhbpuhdODHE+Zy3aWMu9VJwKVPlSJ4UB04aNQ+QnsHpgkSL8HbwXERuLIFvd
YDCIa/WKygnBFt0PCw7jRRn9Ywtbts+QfyeqYUNtlm5eEbbJ8oyv1EnNSsFJMI2tCK9tBdEDheVx
JDyMgqHRs5C+fFSfg+L0zpU8cuzBqEEzVhRGBhdrkw2CFKIFxtdf2t/L/arttCltDUSm+nk35ICQ
YweqIJPusjZdDJjXI5p5EIdypxKNhWqGc5TL78QC/O0fDXkX2C93DYVnqkfUY7kHdPlEz87k+vZL
K1uIFahYxE23QSiOaQJ9ynnSVMmItdVyYOnJV9Ne7GXirgLW+1zPV2EkcHQCtrx6lOyD9WCrOpbM
zFMLW6prfY2uBa/uInJOTOcynl/Uq0p+YqMKTQmFRnJXZDHOpBwKeRlFewKwfjfSFWqWzwlMdlUt
uXRkV33ioXw0Lk3wcs9h2R6mRXuO7q2hURyiixz/1yottwQYqOOcjB38NBkiOQ5f4frSBanx3XC1
kOFVOc8aIKIsSf1MzKqT6jaAS+D5ogB2xM8UzSZvGfY9HNLV3Xgxp2ScrVj85FTUhBWVAsoCfnHH
Rgf/6uu3Ze+yPinfosK/UgQKeuWQ6EYtUBEXeVWGyNg0umKdRv5dgCxbdIxl9+lvvSr0a1ngH1+4
oYzkQbQvS6so9Tan7fPZdHbeAHwc4GZeBkBSKQ1hhXuAGrdalXxfoDHt7PiZdI5o59FrFiX+EUVk
x8IazdnjpGoxh2TzcbDB21ABLkjMHq2vkviW+R47fut5oMKFLUJIfLWyhhPqVbqptZZyCtHpBrOQ
CHB8GMpk2PPgTHHbwgcyB3VA1GDSfUc8t0pDj21daWt4udHFo7f4IAtRhnjBY0vOHMC+A9b5B3et
QpedwnOfGogl+jdBJrtgWcNogrV6CSzlqF6wfGk22+M7VxCr40iZyY3ZtWe/dRNgjB3GtwOWqOJJ
kJxnhcCuWA12qNDE6LKhWv3mz4X22DO9bOkE8VTK9aGDzT1yNXmmm3kwvtnEhAe8Q7FZtAbNLOmn
TFxkNtIO+AaZ+2f6OTaiYlxCAs2BdkXQBy/1XGo/xtkmzAomnQvBF1T5rcmA9+j9a5+kHEhjf0iu
9k12sdkUt1jb/u6j4Q/xFJGh85HLlMNTTqSR+4dXgIK+EVrz+nGD8qtClFYcQ8EKC1SIHNbYIk8h
zA6MmjAHzo2j4Ju4dHPpSTExJQ4TnUJTUA1pbiHx+vot8uIdMjYP6B+RpsI4R+i/B8VGlz5hk4da
JIssK0G1XRdGQghKKLrE49qFRmFr81YovxMUu9CrkgmABYbxs7QB2NUtdDypoFDBeXVoK/f9JH5y
TPWU8rNfTiqTn9ECRxQHivws7X8OcTqkc4ZHQ4bJZlfa8/toJIvpRot8F0nXAGZpB0455aVsj0ME
iD0nR8NW+O7DihNOl7w9FNq9oREPFgbxHP0rBpkfYMQRaGM43a6bUlz0oPoQ7UH27JxODP6jveKE
6MSxzmSIsxJHd3wGrFsMSQYwCe9vlWqTu2ce9/IzYxM6rtpZMnbP13nUYp7KYMrp3m1as9KtAhE5
V8Lnl2zHg5u5G40RiSokCalkNmHC3PvxaWI80S3AVBfpoz7WfusmhwAIU8c1zAV9VqtJ7FCSWQsV
u1jyOHMksqu+MU9dhHScufrpTAfYuEKawJ00vugDMpmIymcc+uwcU9AoYlo1+I57pxMd+Tb/BNbo
kXavWj9ckd7y6XDDvUOhwu0AwxYyOm3Omo3oAfno+TS/21WI0zVZlJr7eryHDTqXfQsr79Z7WTdD
XVCSPaEHUdbwNAqP8aolejhBlcwZsSBPF6KTOnIUxQhBL10+HqSRiokl7z45YdlrAooKWe4YPY18
Q1piNAnG6CQUb7jGZciBsep90Xe2AzCmNRl2zNrwCICoQoCTkn13M4ZHJ3wI+qohhkv40jE8YmNK
uv37q28/U0x7ZFFRj4rCXvGsuFYMBEfecOxgtln3KeqGIokiJ084X0vBO4NRnlhPiCnhlG3FJQxR
4kztACITBgr31CQL4fZtzVkOmSg+/ci3EymnBYwwK0i8F7JKXhMIku4uNp/sFBjvVKyarEuTH5HV
j0+bZJDS5pKCHBvmOlIrpO4M7ZhTyOp0QyJzqCQLNcanc8BJZll34EPm7X2/nfpmDDqPiZnzyY5V
ER5GDYUIGDckcGRV2o8/S4pen0SwioyuGHQx3eS5wwL6Fr8b+jlpZv9ZdXMfRok9oUNJdQIqpCgW
xmTE+/owaSSF4adT00JnBLio7rc3Q7VqjJODgXrraI8SEjuA53Vb+1FNFYmRJlBIEMemIRnAGHXu
95y2MMN/cg5X4IhkHz+i50wRkBtWLXhr5fouSuAA9vS0ED2izKDIKj5dB/dSOm3PFpSQGk2uDrVr
Z7yKlkMKl3IqgHNiCSwIq7Ug+r9F+R5axONxTxRU+LflGKL6cRYhkESIeoDmbm8VMzqMVbRinADI
AoaMhWIjCIiSqVwKLhDKBX0zURQqqsOWUqxvI9Q3yknSYF/Ofij4AQA0/RY8nwXvn2KGNdaMw5/f
77biUv9uqpVlOK3UuFhBqM74exyzcneYybpFLf48H5o1aJxEZeRNg+GY8zhbrsEx8XiQTfIKx6cH
7dHqAObgAXKd+VMFJAHrcCXiFCxF0GaJN4fOLZcyxs/rJXxvC2hKq9dNqncu37SREJU1bUPSpnEE
7uRk9TBaSumLk7bBVwSrc3EcTTbgDv2+nKfjg+HhUaWaMs09FfWmmQGWdvAN1zCX5L8ntBZ/C7GL
+2U5PMWve7Ay9xoF8To2F1PRItsrUsxt6VuthrNX9RYziaqnVMeOdV8GvpD/MES+c8AAp8r8/XSs
cNxpNAiTyShFoRNqqMrnihbdyBeJ34w2URw2O/oX35dpWwN2r+0Z7GamrIUlpDeziy0YepQrV+7l
s4nwK3yIxeEoTPV2v8Vfk3sZIvu8D56XBAl7R4bpCrhUHnmSYqBFdzZoEBhnLqpCMv1M/UsonYmg
gCsZeX4aAOB6iqjAUVfhy4u1Ew63WL5Ywm87DYlK5xT/SbM0lyoQtTVLAqllf7pw4BEX0pljpint
vMKL98FjzcCrR0ivFXYbHTa8FXJIbiA0VG2LSDqgVJ30kMsT4GGFs8gh84YjDYXkUAOyZR+Zw8CN
op8Y92aLsR7cHwG9SR+KS5qjY9T1YY2ntHE4K+hY+9JQxycI/vze0t1kTfU1FJPyTYGX9hHUgBsM
V2nY33inV82ppZA8ngDWm4qagTzjlbnbZqXkp67T8VA4XK4exVpmXhmXJ2jbROkaZ/t8eZGbdSiX
HcL1SZ9WxwMGbTlmfpQSkVw3N2dES0oNt23No43Fkzy4dV+5xXyvzBl5dIf/Oe9SF7DbMHhBTx9I
qX9w0Mis6dpl1t0l+cF/jBT+f2rUTZjJ3E+vLTHQqzYk8ZLSRBmx4DGM3ltPV5HGxQKZycXKLp+o
jQx+LMYSjTH+U+/JSGKFpagSC2v78+MBS89dZFgX2MwVuyq3lXQovG1Q9cALnXF6D3MqNsOEwR4m
3J4G6No29Zyz7tRliF7BAxiNZbs3ypvVJXVlkPjemlbX0J7WsEGjQzBy0z3a+CaIYujr7iUP6bme
l/8GRR7v2u/iGyIgIsl8VzSRY7LezRFLEJc6M72vxWlxT3Rw0LEYWe3UHSVVm1fhQGRz25YW6jLY
ij16nceXU5yzoRtYz0zuWKJXfo24FiWxxVYcOGoZdzN+ctYHr2JFdAcIdTyvsEEVIPwNcDFBCfjO
Z30cP9QlxvGNn2gigkRiN86xgW5iJeRBXlad6UFQzqx0oKviB+aWur4xkDeYaXnbEcAAKiYq3sGU
8XxJJnuEzg2JP/foJ51gtKAoWz6afXQ1mHazJTz3e04/GpUMQZ+S6vEXoh/Y0zz/rVKwlDbI5j1N
qOl4kLhqRXONYdSsMBmtMqA2LxWlJKDJteHQzYauIphDQr5mk3kYCEiJeMjLE/OjqTp27sn5RqQj
+Jiify+notpsOdWOMxIxAf0FvkzQWxUTGAYlZu2zXhncTjndc4d5dkS6CtTu7qcsPX7p0Bn2o2li
0AwbccCg7fujZUEZkL0na1rcR7d9LwqLW/34+rhy73PFYPOaEx/YjE0R9s2Mb0Nx3wrgWKUq4xnN
1RfKq3NAd+2JV+oX455AC3icfaDn/LRWyL8mj8vqe53XOFdFYRrziAM2MVnhazZEErIbR3/lK0Rm
0mE/zA0Sa7MaVnjNFS4Cae45WyiV92I8i6H+WGsRbPLCsPTsxOoAiOy2o+4RnPnLpyBFqXkq33QT
LlO/qkDvEWT19G03vOvvKj0qUle2yxkIBTdjKna0UgNC4ZTvPyYR1ADGzntiWETCLe9PS2f6gb73
mtvPxgqvXcdq4FSKj0BfBP1JvENsbe8Iped2dMxARbHlv8EWKb3F0ReXgdaBugVA3n6eZCVA6VEG
30Ibu51nTCqLPAKqk2g6FRWW5Auga5LZILy+gaaRDCsjZoiNBfFtb+EhCzOU2i/Jc24QR584CEHX
hQqyPr+CKhIY8SPD9UCGazVPRt4QS/WxTXZM3TpoIZYSPKx3Ym/4Xg8HPc7p0H4ABU7CB+tni8WH
COCfyeT9oFc/kmY/iS2OamhnHnUTPlifE+bikjPDwcf7/v4KhMHSs6jCxFU1kaT3/AYnVbVVUlol
jAYSdQ+gJOWVazI/qB6oH60aAg/bOWdjCEWHLUV8/BMAaliTD/NJTni2KbsbiZvRSvzr3ZKzHKlr
gbxPFb5LSaBZ4xZ6wfKl/EIcJEkD+lvG1CDn9dkG8yHzw/3OvPGM32qyNTOP5NDg7xHb6ikO/jj3
8EyrpeLD/aPQ30z2i2obQgSfw8fx6Sp65weva5rjba08vdHK3KwV4G++YUwa657kLmxqaJq0Gr+Q
3gualRtFn+akBO0h5FTkY8OHOlysHVQoGugGj1q6QDZBxfLvotDakYQ3AEtUcKxAc52tpGLIIehX
so5KbkR8WdnWaJ84Wz8Kfl3dK+785QKLDA4d2++EecglJUU1Ej865Retgjoi8LXkuJIuHr29MK2I
3jSWc5gQ41XDYk6MyfuF6U965cJGIdxzo9dVHa4Zs17LJ3eeLlOmVMmv/lxHm6TyOyo5jQJdiZSP
d5XcC+fRYyuKFPRuxZoL/4QqyiYCXUs8nkQvBB/V54N6QWyyW+ncYYHy7Wbq9Be+GfvQrNL8IXZ1
311dD1LWt7NLskYUp7hywMVuqM9O3yQJBvk3V9czBsbbvUfhaNxjjesiPrZC+ZCULIm9IwbHyQ0o
cI/uEsVLiU4uvPGbb8KxDbfGhTdJjJB00dP+E9qz/C4dv//TmbJHKosBP4skO3pOBZUyA7fQeKY8
jSb7YnEjZknDw8J9YJ0cWYJobf9qTdXM6Xs1obciViUYxhAEGHRaTpw1DJqa2nm5qC6hoph/ngC/
GmJU0mhkcqXhFA35iYKaGWgsqlN7KzSW8W69pTle+m2+1+3FB/6dTzP9PGQpIWcYrI3yYXeRaziz
3UckmoB9ugO/yVdjSX2zkPdSAxnMmlckRNCme7Fnw8EC773FFioMMRtCvjZls2DrlwEub5g/y41Y
GsL8Xhrj+POJq4sxc1L5sJ4RM7D2MfvlOZ/Vva/h6A9IaKYm5R+AlDlxV7ItZ2pQ4eLfUwD9G/Om
9XOCSbX/Jg45EglZEwUNSRsSxa+6nESpXrDsGHtTSQbZZKZ/WdU1WkdGkb3LFkHY2ppUAWOmV3Nr
hFZ7E0Wi77k/Dek7+pp6oUcmmU4fQ5egc8+HgidAkftvI9vhLQ3n82mCXiJNkMBKOX8CZwvMrHk/
x2gm8fh4I28NTApyIxbITSYrcTfPgIEyHwj/yFhd5JTY5c7XJD3moAqiryl98d6152uE0kTFhGMQ
D53S6R3/CmaIx36XJVwVcCVHXoZyXYvurVZx2oI9PaQoPZrTH0aFbkARb6KF2G1K9jt7OD6O7jjx
pv5Kc8IXRpT6OqydFI5qox/F4A+/sV3nNcjY0sBtKga2z4ssUhNdhDP48UGsrIHAiblEZWeUyPa/
74hr8fdY2Jb+DmaKiAt1lvEH6P6FW48+sz4c6m2kAvZyGf1JUv+q42LSLJB5UPQ9ds1zNZWvG+HP
2VOW/s7UGNEB0KgtxD+uFihKWoSPbaX8N228M7yF1YAmbjUh/nbfRuIGmXG89ytjVpFkqG/QmOVY
Ij9fjwljwxbXgQLk803eiV2wzT8Sknn2A4XZ3vZfORhZEWtdPMcpB4o9wmoc9Kb5w6gBXGWNBNMy
0hkOaeDd92/4YsQgF5dI/QcK9jrcbnGAPQ1ZvGpbqfepDPl0/IquEGHjjwXlKcAdIvLGBbAyjjMj
WlEZ0oJkJHtnRHXB5aq3pNJwKjSxbIWpSM4yuDrbJSOOsr52hqoZaW7PhKaeQtF0p5SuqX//zdZM
wQ0nKtKyE78id9+xzV0MjUAFM6J7xdTsMtBQQaHd8D1AeKKx2vtvF7/7DeTRm+vH1AJCRwI4V9mG
TU2nDNyWxlZnz9cNrRaKzWs+KMnuiOfjHPFAzEIhs7eLgEBTvaYU1KNSyjg3SiI9x/Rh2JHiynwH
u40H3biExrODsnh1DbtAJCGshTd2YaD2D6bi5w2thm9AQ7MjGn32TpG3OF8yxBOadjcYJyV7oySK
X0cng8wSmrzjIlT+uljtAr63rYcvWeLvj/4tmLw2R1kAQw7MKXHYepUM1yjzmm4KJqvRZJzbZXOO
w2WH84x+yTfD5IZmzqq30d/49skVeb2aj+dBgS/YUuFElNF1P8VMAR4+bmer9QAgC9ztveipv9pN
1U4CryyZgEoYGfpTZcd341SFpYNhMZ1XZrc0aoQLwS10mI1lfSy62dvxP6SHmb5/0UP5gigxNt/1
byxk41/9jJZi5uRECC69msmyN6etsNRjPKh8yuwJZ9pEgVW65Vf1c4DEdVHmUg/XOizc8mZ8GSC3
B+qrS7xFdsP25vuultP9frQ6477dtX5+ThpmG2b44nuJOJLw1dvZN0wxjt2XQtoU7yisOgTqrxqg
cUImvqY+H2JOmn5nfB3MG7m4GIDpqMS+A/EX2LVbGbfP0PJIs1J4NKQ2jc2Nr1bljrsLMPVG6LMz
35u5DCoMtUrgeQsxvwXUFUU27wGtu/6yLe0C/I6gaGqTkYGCOEkVvENJhY4db+L7SMGOquCDakoy
FQobqqmjsjJmRjaNd82jKZbvn2mZoOlw/0Jt68GTuDoAl8YzJJcxPz1tEUqP5pR7jY4dMcHyNJRO
MwQpo0Z9+WEprBIEusNlkWtnQaA4ZGPaTp1XNNnrREeCFkCNCpoZbjZxoSoXjg1xCDINmNMnUckv
KjF6IcjPn+zXWIIsg6FtZVP3L0V6e9sZK/o/EIgFdSyTN9Irotm4TPjeASlvtR6SM9Eh2T5EDVPo
oiIPfFWLQ4ipJkQDewDVa+kUfyp/R2CVCG9Veiv/ExwJ3zZ1czKphaaMV5j5XPK050bQzlom7jIu
KvmvBQ8fj8RYeSPeCgvJ0B5Gou+ayIgwIw+QaadEM3N1dKKbmOGVOSRwTzCwsfWa+Nld85a9OUws
nCmfc95LjMG1pESoJtOT+fX+et/g7uBejFqAHtV/SpQA3LcaO4wuC1Youb08bipo37Rnt9/iOwCB
vA+5B0cYKqpCwAMsW5hdNQLxRKavd+YzBlHdMCWRTrsotNmNxzu+WCSgYdQhasRY7qpc3LzFTDCb
NS2gEf+e1GLbRs9k521mT3YF98uLLdsdR4OjxpzAUUY++zuEmbs2OBV7+hDVhnS1MxA/p8xi3l0C
bqDZynNIhs7vo5chbS8NCHO7vFcDT4jzroK1Z1JJ2g//e+W1OSMB6njVBRi/CfAPX4ezWFfkW+24
JVayd3wXKmw1HRD78MFaBU52RDe5+EVSJYSo4Vxcwn25UDJvxcRX02O95DH6hYMwPdyDFngc4xdy
GMOlimlCpFpmj8n97EtxyulgPxVLVjpscTBjoPWeVsG2/iLZcYCAV24aDKeQgB2TZ37OjyHqdQ9r
+zsw9sPZfla7FPjC6hWc6DsHIYiXPN78y3D31EB49p1G6D6+0aejMocd1vnI4lHeEpPqsFyy6PXT
V3S2XhGi4L0kTFf4q3meUQ0P6iXnWV1iPCEcbFXwt59nzdotIv/CJvwQqY5uBucJSIYzlzCjo6s7
fq8vTE7EINNzu+4ihYtYamHlRHDZZhlXQni6S0C2PNFEYqUPhFRZlAaToFufx8KLHR5xMn9Vl5UD
ctWEQq8BKfgXv3z9tpq+/sJeHpU1o+0su/gpTz/Du9vQl5TBQiMFPUefuRBBpzN3VqDvRWnGGLtB
tVuqKOG6K0i2Z3bnnLTv7tH3CITFrjDlR4xUr2iN/4rxvF06X4G0ITaBlOE6sylKezHVV3ler83m
m/Z83pzCP1h/9FgI7KDR8sXsHozyezfROIcsAfS/qP2ahP5xp+HP/BcSPtb4/b6rTQE8d85S2lq2
nZd0AzOzOV/IG/Xlr0jSGWlScNdmXQDetQwl2/z3TNv2xZ/E06BlZKgZz0zRGHvT98D3RUJ0dRLS
T/cE7HxE9DQPJEUd5BvQy4DWWikG+tdMXytOVSLC8Gyua6UcBZ3DdquThliQHxIMELYmD8L5FTvP
ZQA28WXn9do1vXbG5uY+56FY8WWheJVXFVombytl3PR6HvG5Y7WnmC1cUyBOmm7vW9floo6w1CCT
Lh1S/PqafE9lWWHkuioYFeEecj/D2gB6WGyobjp5oRa1IGIGUbomcgN78d6rfEF3ID5Pb1jFK0ns
d5gb//J9cTPOVQl7eb00ATuXzNjGptqwyLPQts4WQJI/8AK72hyK9DT3ykVtaE/eQTYnVG6+MidO
eFCMwDe7fWRvdClDNOSMIPfLU+NJ6t+xosIMwb44Mfh7n6AW7co85USrVqC8IxXepYpNePFNqnaU
a+5wSCZZR8ls7pZPV1EV1vzik1Ubud8zOYElr2X/cYlAvc4YXbn/rUWXf2yPOOPhpS3KvQbltbgn
lo172gxVelfJrBclNNQ1PF78TCKv8tMzhmebwIDYLA0hVdnCJ82utlW+aDKLb0/1aSg7KvUY6ynr
ckY9fTMVuTH4HYcyXzitGMc3MWzRL41ngnmCjXO7cpvPH7ZWA7IpZc4SPy/lsbC47LZjvfLOnRWv
z2icLSu3UoimCDUByAeFDIc1E8UQxHynHq3J9587VysvsbI2CBW8AVsTBaEiyxmXJowyT8dyDrEf
Y4ohnCfzVKkNyIx1Ot4ms6F14WhLKwVUcJVaQWDJDkW85hAoNURj6d9UBMkqghlTIzBfiFYwlbLy
RU9sF5jTqBcXVyoMYFT++N01q93mNcY6DR1koZManvnM2J0SHIslZqtHZgL7v1FEyPKKIlGruuoq
AVKzVJSGTnVTkFloDRMrNfEc6jzWj+i0xiIvNLzuj8rRMVmGcRf2trB7tQfKfc51NFd0ir9oB0d6
HzKPDUijvc9tJLBTUPfmWUkJjJAr1B5axfOaYFkPYBwakPqhUSnk/vu4+yX9HTy4MjyAxbUgfEom
C4p3ZZBdpWhLCIXvkeyfBsckBpGN2lRP4DKW6NBxEA0gehoNKcFO8hqO1nPziVmAFoA9uKgXtLBX
Wcutz45qXJx68TZHzHqn0G9GCk8VQYbgx6BNzwruyeSETsj+rVoOWf1Iq0jGi2yvuUGdpPBpPn+g
O55WBaZGPA8BDSRC+VvVgaZy8V1LeD//rihEAxFmsE4+b0NwTUrztKnKfgntT2hQXjQ2u53hkMWU
G3btmlhZiHYD+sNbAAHr/m6YzSJOu+4KkoeugEcl1ancPW6mHuMMNLcwWwxniYbxpclzcTCtvdNo
D8hw7mmFMrozkRKnsgg78iuQCXAmTa5IJVASgtdu7PHb7omP2GvubHcRwTxQk3K1eKirYSl+BXI2
1McYPWV5n/IK1UCvcVL4HzkFF5upalSrfDrlwiQgbPW/CjLDJ5ivzfB3cLEdT0Vm5DIGnmIPEMBR
F/ygycIVrsfJ1fi4n2SQw4tR91CK9rFg4Z1IvHAPZRazZI4dWn3wM0VYwq9nZsxcBSqPmN0p18bQ
yNu0gjaX3rb8za7h/voessn2lRfI5PZCIBuSdoz728SR58zBXhMLzt1B/ZrpL0O/9HJOw59x30CG
tyKVWrTvKLzn1P8+gPY+vtCYolUSMz0lM60QZ6uWgnLSq8Ze8GE3ChwS13PSi3cNmaeEIgzZ9vi2
yqyJZn7Ji7faQNQM0Mp59Dq9ziwfJFU8qrDgRK+FL4+57ZD0BNTtCH9LABNGc2iHYML9ODY4+Zjz
LUw7U3ovcC6AGPL57RTdRjv1c78+7KPaSRyHsJdxi7+xZbBiwh9azDqGZYVHE/aKeVxdE9u/mcrj
hTrqxxFNf5elF5X/qfmNrv8XtZufQga1WUa8sM+iA6OU5ICAXLSCXol8A0hjyBkI+EUDEdZJgVrI
/Atsw5FccYtM32XjqWS1NHmOKT6K0uTZ+mvT5gY83MxapgccPqtlYBV+Yyrp4MOGo9OK6H7HA390
rBmuTNfGDVfyP3BSS2KktrrlIuRxPkaGs8desDBfRIt7kv0LQz/un1/vF12aqV2keo75z5PPDFC5
fyE3zG7kkunGJ1+6oH266SfbDUGMhnTZBd8eAn9GtQa+9Eyr0r2Q03sJKo7vytZbbDcS6z/+H1fI
1OIwUSlJeP0O4zmWuwWnnDwAoWSJe2lv59PN2T8ynVynfZcApAZB8tob7/dncLmZv7eWRmjdDezH
rGqHA/DGBV9hWGVYNtzTbnuPZ1KRR/x/lf/GnMxgfoTWYX135Ap0KkmSHWLn2ZhW8fZpdkTP/B7p
u26sMCRxYldXkZMRb2c8SJS6EvEMrN1khPimGMiIfCh8XqvZTteV1jP2cq/nzd7fwZU5SyzeSbQX
+Es7cSvjk9d9TJ4c1c6l/EITOvQayZEpqmNl4nI/QifFAiEdGyEG4254+GV86UA5alDqYabLboN3
ZNReJNDHSQCsFL816wGvmkoWasHHN+Ss/JV55OZqGllvMqX3YNJpuRmyuikhCzXlWQr3DiV0+eRE
hgHhHbmaslx5itTwFmWsVWb10RnqCmqNW+f2Cu0PPplLcGhxznadlddq/AIZV3ML4i7OUrH6BmAR
AMxBqjIuG+++Tzvxme8lFFScuXGRnH4XGXqdDvYqjj2CzuGzjBS1trRZwfnDeOgKwa8XRf5fD0y6
rjjFxAZohEIbLqArwQyOAl/NPxcvI2LJ2EiEZtF9oMmBMwzm/X3+gxnjJJXtVPqvbL2A4KmfVV5v
Mm+1QSaoI8G5Icv6aE7ZiO5ePKLJ0UaYyUcP8dPBQIGHDY4jA8eduSNxs+VRBKZjdyTYKDW/ltri
+RlAhkiR1Djafflv2LAupqr5pHjlk5lB35tXWTHihLVHuJWCxADwBXQDHqslZUKykXP/uZh7M8sP
8kt8U9GhtVIglDU15LOub9QC7xa3Ubw7xD+TxoqDD3TUf/LaqF7zdLNvtyoA35swP4rk73I2R2pf
tW3kYtIUQRNHVeFdpW8tyV3X+BLdGh+hjT03XIwaptrC5AQ00htYTib0VAV/s77ky2gkv2DeFa+j
tyd1R9oEefkY7Ib8kLVEKD3vS7A2g4EjyqKga7gGfmkEIbvEkG0Y+Z2zMVpYwSfH2VdyMZarEC70
AOXRH8D2tpC/NK+AHn0djcw3HJK0H+GpRfu+LuRLICourYUNxGbAVu66/ekwvfbrPoHLVV5DiePc
h1aA9FJzrWYIkVOy+ONtKFRgS0lP4/Ki4aaXOUH0EQb3ijcP4L89hZjNJRuBE9P01PPGAAWlDDWp
RJY63Vh2pnWCDKId/tFqY03A1WyJJMOqvMn2ZiRCM8l44k+Wc+hoZO+8vk+YAvokY/KI8aUfiK71
u1P9AWalvTnhq/aoLY+V7SshnM4WuNCt3bFoCL5YuhVHd+MiRRt62G2huK6y086ErmHyY1oQ/NqZ
MVibky1IfEMsHK2E6VsjwcFBqLRd71NZzx6HArzgDK1cqTRsr2FpAycRdiuvBMxeZpNuKW9qykzK
afez002B7VjxLD5rt6PHC5VOWyuxJKSXzfm7Rfmwsj4N2t5ynAJlNLJT7qEDCikCLhKEoR6lTl3B
se6MAsdP/bDQ7X3A7TPbBIUyKrDKA/14PWtkxSIrCOcYxRzr/pxbkF8+cNRrIZ6HZGRVpuGfmPU3
sTHPn9a5PXRlTSk6V6Xct/iyphrKENq0DGoijMKOT2oAm1k0eClonwoUiFu0ls6HukJ4qBrqJOkK
OeNsKaJsjLwEqhucma4guFs0v/3kcWYhE19v8NYHonvCYl0jHrPXAppKbTzeXzFKBCE5KE4PaF5t
ZroDKW2H9iZUSujCAfnY2jZj35wP9uAf6gSBWjaaVAVVjUX46IqHYyCEooO4QeMWZ/kwb0Whf+aQ
gazqh3R1kPM1AG1g3tKMqraeOkaoV1cjWrmBBvZgDcE226LrmubcRjJxUHU3Zmev+nb3DwkTl7OZ
mB9bh1yFr59SXr4fvgkpm1RIv805+zIduKY6Neobl/hDXkMURrgMUr/TdM0SgvSfIGcJ4IL0b/GN
6Z1w+IU/GdH94FXuKvkc6/W3TQR1dU/ZYrbC129aLbcgW3YIl7KQyTRFeCVswFWDuFupzPUN6su+
3Btr/qIecp6gH0a+5p+/DMRAOJBIc4BriXMVS7G21NI9ilt+WJP9kAZoodrAge1efGof1GHNlpaV
BpdR55nZ3iQsLuT5svqYPX0g6NGsvc39qC5JzL6j09W2siaBhB1YLO0TxQ0HtgFZf72aBy0KFELx
+iyRydPTKSRNDsDbFKHlMsxNH9MSTy6rcDLCez2AGT/78iALjzlxt5GFcEFk1Yv45e9qTnh9/mIz
HKGTJDVXYh16khA1XWRIFsn3EtRLfAwuqvEWInpAQqjKLuL5/tNGkG+p9mm7D5wN7A8+OkEKce93
HDYO0MO1RshHSQBktrH/5CfLP2sxnq2K0iTAJ01gdRS2gI36lChgCDnW+7NZt3+1mt5A8d4ZIBA7
EtLLDCRsGVKogjHIYVw9KjEAI4u7bNqT7+Mn/vL40IBf6BELgrfsGOZ+1JwwEIyzP+rhxf5mrZ+5
s+L3gXkDu9vfgaSG7jo5qjIXvAkXZZ0/56A3HMg5MqLfHVg1CINInyRMdNyQVgaZKwFNVAG87x+M
YdXvhKV87wedwmdL4SRUSI4DsD7weLFEbZ0s6ZPonuca9nDI35sYVlqTnWprNZFVK2t+9ZretqdA
PArhlDJl5CFw4zbXQOQ5TTy4meV78MnfCuHcPzNRqi+Zh9oZ3YOTJElJY9/cadgQNkIHhOMX+W5N
AuKu4EDtHBB/28nhC4U/Xho2vDWRKYZ7B/zUTHCUkCnplUINOVRVtj7q8/KkcsU0dOgXdOp76C24
NOXDk4xR4J4OcQPBYyIa4eTI1q9T7cEvGcW9ImAQmRDFMiXgws7jYfRIuRF8q+T39Wvc93+Aa3id
6NiKk/AorwqHnNFT4nE8ndlwCuPHV8RhYMMjo1Qr31HaMxARAxlAEVzcR6oL/vLMEBlfki4yLyV+
NRx6kITLEFnxJnBP+R3q7u1ymDdxVgWv2CR3OJfLul9I5B0sQOB4yv1wIi2BptV4N9RQGkddfUUM
7SALLaA8tfaVPzjRCLMDOvRySVz8tRojcRIUOG/sbgYv4jQcY68Mh7OmYCgGnUUYcZW3MSKKkMwc
zpJRXP0xKrBfXdQn6LpqZF8TSKUntdFib2oVUjNjDiMhpdECmh/+IiW0GKk6UCBMB55o7+LvzXge
oHkwHIhLtDVMU+h5tpPvJl8oxE4T3KDxsmd97wN4V+1viMNEEJPPhJxygKr/4kGfen451p/vI6ex
9iPk49njI3SbaogWEWqkWFNe5bfK8mwBoZmt/zFME5ZwVe55Hpp/Wde51THJT3ulK0ZCgHqrwWNj
EuJEFPrr5AGFAQuX5BFNc99owQrZtBDHPYW6QRtTCy0NElN1P6Y8c3QPJOVbtBBRk7BMkZPA7NJD
rte/mAua63GPnK1kWbbE0IcdSD4Uv27qBFcxvWlDCZcPFn5nDrnpiskRIYJnXyW7GFWK8q224FL4
wBp8amFWPQjH1KOkwoH/Pt9S0zzdeY/d0eLqY/WbOWdNE8xhqvp0274AAk0gVsW9Y2XCoJDROT/l
gHHzXwRjoglXB7ecV7xuotOtX8KFR2xPlssC4HgHWy88w8CS6dx0863JMCC+z77FfHr7LqvPpigx
obHpFNa2Nk+MmwDO6cmteZ718blQIsytLFs47VjXuDlB3oQR6g6IOBerUv6MR2sCg1MDx0j1x7H0
vBfA2dqXgA4hkXyZfGtI7lelQ2yK1dO1tTHmp16MYmCgFx2uVrDopU3mMGv8snjQYf4woUxYg03v
9CFQfyB0Ab8lJuh5I/4lgdDLDXJmOHzDmbUqrlS0ozPISBnuhrswNhDGfnTQyPtPOGd5Soh87Oy2
vEDi9fy9LUIBmwVOeZWenwkg9GOFZkbVTY+O6GIzCYFDCBB0MIvj0oQ14/WGUwtR2UxL/ycwxsdI
9fGvCRzwOrg9O/hWbQ/di1voIRc3IEpEb0dcgpT1gncgYYkS4x43o0g3dlDoc2ITWWGE9sbFtX2J
cUHUpqQ9u2zAFNKDskTGsE+rnHUI5jzRdeuTIioZgI2G+MBvbFn+Z9BmcKBFTgDctPbp1Jpssj2t
7dpodYEyD8ERGvQYdiQvgz1JJpv4hTvdXbA82tdZnYVGE9g0d+c7JeGwN9e5ZD7MgmZk7pqePMG3
ElRGa4yJrZ8Epnz5xzvvP5v4+gGI/fx4qUn+b3WEAtwRFIEJpbGs7EgEwkCMIQWF3DZwJyI8Wvgx
4rSBmzjmX0s5UuDQbjKMkuZ0vA0aUovVC3N/NvDqR3SFkGGjCCtc0dgclQKbrDV+f9zRjWc0TW2v
ScS04EUzDQE98Hh5MCWdV/pWSLK+eI/bMvDEmhRV2VE2OBGvXoL5u0px+Dj+h/jghO06qIaaUQvN
3yX6waCcUH2Ld5qlCXnPpqUcEHA6AfPX4C2EySyQl+k3KEKfiLvsbtJFY5GYbZof54ghyNxL6ltz
2RZta2Hcf2JCC9v43cHhpnAGbsnNrma9t93n2lVj/3yMoC12hQ7OXcKHcQtz0ALZMwy+yjVKkoQw
epC8putjZfH2PA/VvEhNG9ChM/D7BZhijEZ7IAd5IIoBY1ph88LAghlnLkuMvccWwDBoEwy4gd2x
AYaxygImLzcUTmEqSzD6Lymedt+yyWZHxaBqXwCAxu+zWpw4yRUGbnUdLJIzGY9v7o4q5f7/2hOt
O2MCxOsDbNmg3TtBG9kA0HKwsrWKsYeqvrYcxk6SO5KPsR8HeBx80+KSxqKePlhQbPAt8xcpo71G
OiZNqJpbyyDdf0I+Ikc8JqK31A4nvJpo2vzxBk4LxJHQP1uNJ+dgFm0XOC55D6VTfywh+BHfxDrM
vLtBuvq3+PpD2z0ue7GqHBYn/MZYwGdYmHEkvP4onbROp0raf1Y7KovjTvfzlN9WHeusXjTON1EJ
0I03E4WhiKJK7mMNryJHVrOCaJ16rOrSEdAKiqxoxEYR6j64r28cPQ11ciMdZfRKZMo4+qq3rSvZ
H+PBCnd5Re8ujfSHtbynHl1HG6Wlp1RM9cn1xF8DrHulsOY9MrNy7QzLm3VbiQ0HovhcvQmVLDNJ
8jiud29ZGwUUTQ0cRizfyFgtv+39KPrxpb4LvkKt7ISajQoAEOHYp6rj1IWgv06kziTILVFxZgW1
Bidr6ymA9ndrFN6RHV72LdP0YeRJrp7dbZWKos6E0yMU+NrNpu4bVgpySnRRlfFtdG3SAuPE9mgL
ftAcoXp00/FaTgJEm7r5QySjzUvgcEYIK2KMQcduGVBesUm61qKaWbOBK+P7ADahIruPtoU2oBo6
jO1fguXniaIe1EEiPNIcHXWsFbaKNXqDkH1c/mzCFfWhRr8OPJsc/p4zom1eTGc7e8FLEYBCW1Wb
s5+3YVICqrOgIG6tQDb7CThqcW9FG868/2Xl5LBkKsQLcyHVYIn6NmkNyuwcgHdugFydyY1hQRVT
43ndXuom/bWlF6NM0w5R8PIMqM+6XHe7STC20xR45/GyQ86myrkdY6A9LhPGMNcs16lL6LQEHqO0
+Y4JJ7W5Hux+tMlN0rmmbznRmJqDbEDxwwo6Ub/pnB4un6M4JK7LEBKnsbvzxRBWz7SaFuZ5B5B3
bIF7wZnnRG0DFm+pyMZFvHmaE8rb0ZTX1wslOrVWtATGwsS47oJtwTGgumASnjbut6jtBrROnFrN
bBO1aK9UyXGyu8csKZtD5QsWR+DXsWPAqRiiDnASTujO/PJCqqXwKtB5S6fkgNGmE5sgFbrmgs8+
Gua2N5M8JAkqUHDIL31yP4PcRTisr6YApMx8h+xhvbNWTt03b+4GMTWlklI201XsDgLplpUFpvvf
wGIhyraiwy6HKYjUVe3vSiZoId15RrO50r0NGdNh9ruqHmwW8YG1LjafnQbu4fncEP0nL4W8/Yix
nAy9uej5srqcixpBdBiqeGfNlbeUA+2rsVZ8TjjqTs93GSjmgJYJ7s8w1tu0P1OvSAbMZXzNkHD3
Cj41TQJNHIbyE/3pQsZELBGiOuqeabK5yZuPa89w595AA1Po3B9yMF6LvkPrU0//nbl3jsX8pQjH
6g04nTHpi40kjt8RF1/8G5ywHSouT6X+2Qz02jfkmkeKOBeHbvZzewUC7b5nSibzxcBXTR/nJxVa
a/aoYKMJvDxe9Qnv7w/A6Ltwlc9H7ak1kbo+xKFMxBXJ2UsL3ueqJ7z9DYbwJ4iK4Yi6LyxY36Ha
Hl5tv9gtEr1qsD0mVa8wqG3O7zG4GBLzc2uq3obAX9rZxm+TmgDGvg2UcXDmPzbMWg3i6TDoKrfy
OVsU3L70X4VuaLGpa0JMZD3bH9Dw6rdsZujlcsGt80jGY1N4Ek293B2HMTi6dJ+GTyxuiWKcYLp6
B+1iub0UIbJ4s/CSmoS61KEK1CA6UrfheO08o/+ic6zpkcpSJOh0Jtm69NaZvqNzcUBHi9z2UrZG
XSslMWyB9ZadURp0KUamQ8JbH3XNGlg4JnpoNOS/3wWwep4vKs6FprfMDwWw4BuFQ2rIod+2NP7m
7ZG3YGvCunSxywWzs/HCCUggbJjGQ9m0o9b5FE/GsC8eG64fzNSpQv+IS15OMdInz09dAfmE87HT
pjpTRGapyIWC8OiD/D7BMSj1jU4u9FBHDi+1TVfFq42snpC6rFCuqOhoJP1j0FPJFg4CzwujuLj0
ABMeJlz7IUW7/LDOToJUs9sh0aEVGGTyTOFKKvzOxIQMIjlNasjs+qbzWvBAoYK7rWRtLG2nAqXv
P5kAXAPkqz1z1HndiuQmQijCt1EM4c2yO6O/i5Z4GUq7NjaIejdZ3AX3WTEZqcPc88TR9f+KtngS
SQ/LnRBtbaA0VAibpIU2Q/GM0aqsQp/Mo2KnvvNZp+Czb/KIxjaQzRLGtTZY2eJYLTRWxkgDOJ/l
Vre3vxaiKoKGz0rZtfoXsJurOH46KIBCvdKZn7i3d8w748tqaTQMfWjRPcIkRfDop0ClF4onPEjW
pljh1cY825/A3wvoIfxVOhv6XOkeGTMty/BJxWA4teAtzM/XMiQMUDrtDnQPbH4Lmxg/wJ0o9ee3
Z5KdopLxR9f3o1Na//OBAnHEVsm9SQlO+y06p9iTc2Nt/kE9o84vOGop/wzqG8wPrwVwCoN2fDQn
qDfOs1hLmEwEYklDJMyJxmwj609BY6K2TYLKR8cK+40xI06prU0ymeJuycMHv5+yJ873kkJ+q10M
EwzZtYRhqgLvCZHKQ2KmDLJFTAHvLza+DpzPnuR5ZmcCdPrh8B1rF+T/2FfdThgrimEEpXCqpelV
jUpVXthyn2KmeQSVP3JKPLMMX6Vyytf2PE37A1D68iWGcSOXDYDt3A0fvDtEl2O2KVaZh831yCG+
NYuCv5bsPeJksWZjrASvkxBA76IaVJySivL6zn13mkYS6uQiSv4CSRlUgyAeroglIG9gx2SCvhQc
fAZb9lm8xS5zTAkx2rEDiAD0WnKas87u4QNR/xjoMq7n1txsak30jN6diHAudRu4iz4Mw+fsKFkv
yASZkDVhrSFPEl3uQbEzJW9oMlQqPaSYbSANXWGldSLgeGsLtzPa2Mk0fyIjLLfb8m34OAX8c2QQ
Zc8hvuCASUoNU7V004qOSDhNLwd7wFDa0U2UsNffpthucUxG72lKaB2tblG14X3FDA9PtFLk9x8r
rtt0/5xaio50TbSxjEuNh05oSTeCa4G6VNFOIOGywQZdmfNkwgonoe3fiCoAmXR8ZxoIuNHoequ/
ZtS4JU3ofquue3/T9ZAxqkeDUXj9afdP9bSy9MHW7wPqO4FOaqyu4B8qNO51dckPB5lWCOzQxWwu
k32bG5DiBQLcX7ULv8GhVJveii9+4iTqmvjvpQbGUKaKH5g/KvJSCJ9KhuYV3R9/CUDcjl9FyFRE
PZRyiWvt28bp3yPV1LK0jAe7hErYoqXsE5raki5RLw277UHmQUp0BY/EmzoZM7wrZT4hFRr08feQ
OuAuU09baYjfcZKYUHOEm97zXlPwhfdujGoSSHZZFpf8vMej6sypE4c8L9HZVJ5o61PsVrujGI2o
0j28P2SFe9XxpSmAqsDOnIBhqBG5vyd3PiDG3cy0iCpUk8FwKXQw6FDI8Uck2X4kujr9rOJOgT+w
2pfbI7dHtaB8qw0FRSTeQYzVN1i+lix8ID+vdU18eNttyO1S2MQtHK7NdxBtIBpEoWFI6QYc7SIA
VAM7jMBTkIlR57Kyy0RtNWmTP0oPOTdptgT4NbRbsXe7acZcSOqS7TR87i2+cHqXTLq6f4Y20rox
GSIXCS/+6VpTZ1kQKj9YH8rukZgb8TeEJQfuFO6m67lr/TETZqaRcGTqBUF4k6Q2mQM8eyy/0vQ6
svRv6kr+V6L0x2/v+U1rC4/OtLg79E8Tss/qNv/E2jmRkfacvIfRl6yCQCSE8DpSqIvAkQyNePtN
NOtKJmY2amctVEV4sTwvoYXymCFx9mLlckOGMAtltRi/U5igXz4MAHGtYtEC5kG+Sp9x8i3AaJba
2zKRmWFh1ia0zx3gS192cIaixAiSlxycXwmNZXa5LofbC0ryrjQsDMqoBDMuFg2XPIzv80oKuNcN
sY29vbjrh5EtMPjr+/q+YYRKKkYSEa2dfawhJA0hq3ivYB0l2eiXlhFuSSMcV5jdLp8E8jK4sbOb
w9f07ShlHX8jSyRMUNrxbQDfCsHoft4bHUCi2taoiNt6CdysNTHzC7AL/fmWuLLk25JT1aEuBi0G
iarQ/RTcJGjlJt6MIjqBVs40tnj8jfBWL2/yKRv85svGUzqAkru1dYPRCrfyC5+Lk9CQ5+0NDJya
k+yVV0lkUdVo+cTvHOcfttHU0rdIRCRivpid0vR0en1zFWuCofE93eEZapj5rpR76/hoNwqw+lFk
nQCAWYZTyP7Imhg8C/LUg9H+df68Ay5DPXNZHFxlZxBEOxiLbnGlV8or9zVH5M6er6m8dMm69tuQ
qGUUm+PCgUJ3PvScUxAJklJpJ9yZorTLzenKdA37gPgakGTfSS+y5DCxcwryUAvtIm1l5sFYNb1d
9G8wwyLpFLJrOaVaeCPfg5AI6xwVOlTrPNgx4hHS1xYryUmuJR52ubuPZay9gpGDhpct/hFOjBFj
2vo6XxoHLsUZ4FlF4nZTUQDd4gpiH2FGv2o8Qo9oz8hwO3brXeUt0opvz6r3WGHf4NqYPr3mD4HY
4OtQcfTUesNyPfOinj4v/P2oVlHZiH7UQ0xVmECn6EQAcq+DTEmRuEymusvKhmVqqQrr8KeQa/m2
zcUS145Hp/zke6HBRpF4mI5zOhEvKyDoTWgLAigXbBJoOfSwqKNaNLsBwcdUySRdj+Lppe7K8O7A
sJsbMQE/C/WQpQyy2nwrlTFUmkIt1SfGMA4EOIvWdxuMfMmhIZTP1dWNKBkWEXL6LsazwfiAH5hV
q4uMHbgVAnYzKVjRY/mf7xH9fxOm2BiuramP+M8Ig+f1JFxkfDvXIKZsooQpL21Yw/ovDp5oFRZj
52tkZLWzgiRaT2Oh8Exvh7D1XoTUXYRTRziite4ieDqYai6uuNKgf6h/pX1lqYvs3ETGBhzZngh/
NxNqbx1ighob5Hq6y4tZek+36nlOc50/1t8MzDBOwW2f/1B8hP3wDPSw4yBfYmgQCJnRu7RGZ2+k
k0scRvnv3tfhhOQ5zNGYr22ui2+9lcHQW5HM/633Pl0edyhRd3AP8zsjkiYqeaztJ2WB5ji3A/42
vUIQWsfOjCvpoFLIzFBS8PMfVRvWc1XpNvwn1UivtLvNSbU6CImY6UNjGjgQpaeLvGpLjLX25lv8
9X+XY9AkJHddj2Wc7XwLHQpgM5d62m+hlzQ/GLKWf/ipmtnMNHLhrDRHwKTlYhfKNDZXxrR3qPZ3
/ZReS+Y+plGHD3gIgGzdYjd24QAHyMkgeCVrhgt3rhDmxXIsXSS46wm/3BQYs9VDCfbhn++nXdVQ
/1Mk8NANJ1THP33+c7zyINSURe24ssZykdHdRYwAe34WkQPUm534UfX+zfWegO6SvwCI9VWJlclx
L5Xghr7JYuBckQ51ipLtt2/LxTI+IokJlnB6iuR3YKqAW60s0bNIibEGWdHH3UR1wgWKwuFEDUNQ
oaQfwUyDPZa9bqzzKZ1Qg938N7Axrv6HDCbTaF/eLuHkbLS4AZAf7NZMRAccCSS2UEbcyQt3+nBq
+yjoVG6JzQhtMU00/V9zSauLT+PPArHusvAKYsZlFN1XIMup3AHAQnrRMaUVPhe8O+EpnErs97eY
eKFbT+5Ri7KSufb8gDrTaWSHM9UXS6B7zNuFGOCoDmwGFU02gwEO6RFef7rKfiy7j8qkEp//NWzE
0YYcTJl5d4PIJKqR64r3wMCa/SczXHOJq7i1DtJcuqR/fBYl00VdRFgMDtGZhdDem4V8zU6NuqG5
OmgcpvjaKXqzw3+AkYl2DqoxSCEbgeI718aVLgzAy9/soksA2tyuQ8FQu1CjV2WD3LCQLedCnqfB
yaiQxr+T0cKc9dudqC4DozqlTdtTT8sKUdsf06TldjndHcHioHmZ76kk24ldTLMovfrQlx6o5Z2k
mWJnC3U3ow7wrs4fM9V+X52UrKY/GwNDVhpndtibU7lNpo3pzjdgp0uRNaL8SBSvBY99EmxSHmYt
XN7Y0H/yHwSmwzAOQN2ixrWtxcqLGjzHGndy+kWLU9BpVQ7YSvB5l8rpEV14OPdjT8qFRvhTgnIm
6oKzF0+yEHyKop5qdS+xZ9d4/j0mB1M+1LGK/NhzwF0WdRxB9q/v8vX7bVpwv7n6efbhrmo2CZwH
XlGxXoy9ZRdVaVNsHjqS6EB3QuXLqMZT9r1fFMh/aLERm/LLKjBLzjKXsm0J17etlBWylhqC/TYM
0c+dPtPWaJRfE93iFpH6SmcREuR/VnNzOIwUtlrfrYJQvR3K//zPLKNsvphWCgkXB/TfMHDBPWw9
tDmh1Hn/48VI6fm9USZIfSWuyr/DGcbD6FdmqKPaFbA/iVZUIcvp4Kh3tl11RiUvWVv9d26MwQmJ
qRHg5OMcjAs+ZUpClfpjRwvdGSZMvu6EdTGRq37P4XRjA0oPzGX5saoy8VrAykz5HuLTfG2uVacb
PTOqZyp/OOEvFK0yPP1tRrp+AHUoqCtlNLAQK8rVT78xxfvF42c6jhUwsg9ymNVSW7peROBf/I9G
4ESxvqACyXwjr4AS+t1JYo9irXtRo1/VfZ+/BNeRd48xdQQUKgrGfCLl/OQ5NacsyJuNcUJkFeiw
PhWlK/+yM6piRz2cI0U9o9jDg33wz2OZvTy9IPkPtQOwKqfaaL5EyQEKVs5uHsbrpO6nS7XahcNZ
nxwp5fY9FK8q5WStBuBCfTgXf/WgPSteKHjNbMXnV+5SZJzkNN2qhcPSTB0NhAqPmAkSzFHsviHH
5p5i44SuGQiwYJNhlXMUiZb3yzeotL5PDnlIiZjFGj3YQBC8wbMxyDaFqfcaVVdSoM9zE/PaNbsQ
Pw4zgymBvC9PJnFZSGsscsQ4QMggzBkhrxbYd5ChS+b/UIecDaGWjHRxx+HIklOAzODoo6rQ5kmb
7EJ8TKWBnUFWOZiPoYgJKUHf6Oy6+REj2eI7oe2hi95yr1ZLF1Rt2volGXoHXQwqwFv5W6VQ2+fX
vDP7/nYP4xYwgJKFeH0t0YLjhfZMPd+8xnYxdZSZ9K8iAJh5KWoHBlXcFAeUNKA27jkbl0kP8CKW
ykIu0skAGAltAXFa9+dH1pp4YSmFjKiubP89JFsr3XjLFmUCXINBdjFpaA+6oNvyoHYElh+UeNZI
XY0vg9sfHwvHfkNIMey9hq3QoCwgdR82yQXMthdTFCfiZtVYPo7uCNDbUSZy0t6p96tZRskuoett
3M0mxfnYcLF772UVMJLHDgAg4+bqJLNxsi7HKSkq8Y50806rAQqjSQCE5TepIBHhVqodrXNCWoJF
YUFSEzOFOikO+9le40oh+ITYAsAyqOPF8q8JiY7NUtxm71ovQZG/WA4Wx56ffPIw0dQMXHHwpylO
q/XSFvE5uH1V2tU8PZDbgjQi1lICqbRJEWjykpUR2vfACxHrhovEWLPdBvq/5eoM7mKw1wM43G/W
JO6vO6aT8yCH48XvZgrfi2BqKaoNRoRWyRpG0aTMeTzr/isCzldWq+oUQqhj6cVwSO8k43G2Hkzy
Qi7BCFY6EaKcziY8WD1iukOogBkM3SNWHEnZbNa633sfeLo887RYeCCOHUIoSdfrJ8uZ9vS7IpeJ
/iwPOnyxJHeHfhsyQnSINdf0Ar8W10GV+YY2yyRC/cvdO5VC6xi3y6XL9zUxzeE3rn6TsLh/2cnf
It0HSfw3ZwErshly/MZ6VeX57/mfZPgU1B79hcJXoUuuKG34hvJoY116nIz1J9ZQKoTHow8anf4o
SPNSNW/0uKwydzRti6CnanQEQqQs9xIphw1FTt5o81Wff2zxF8uPYBOejzVHyXRaQqzA+vaZnYNa
/Zq88y6S5J0h7wYKhtda8xIO7lpx0JRwY7TrGgyNacke8mg5Z5XmxUXiUsN5fLG4u8TfQFlWXjM1
EIsBR2ej1Hmwto+3ni39F+m0m2qzF+qDNKcjkbMw1xCMi8pSquCE5vOauFzYmX+q34NjF3Yc1gnm
atkYwVAOGmttitJjADy4T0rlYiBpKw7dfFjVF/o6SJgf9BJFvgSgjLm0kncFH+wW+WxdrmHD3Ewq
s0YIC11g5VBGydspr+8lTozvPZqtMkwKd3GsVVCl6/4pFCCgv2ky0t0aHP3gUbWNinj9O7kpRCSq
FejGB/ptVxBS2tyxYlUYb2gCaRzpHIVWcIGMEzBf73pwgRnI8NCM4k3s3ByNn/ani1ZA360U3JTs
0y7iWr4KeHfpR/63hkEoRj7FTI3rF2khn837JRLTD/WTAO5Z+CnD5ZwKZI7rGKbFtx8i4N2mjM2O
mELR5rYMkW/R5+QUepdr/WZwlJvdP3NH9gQAKjMmr5wSFdsr+w5Rd3PXzB8Z2eNG1zrzl6wyj0fX
mme4pIY8cqVmAPkyX/cgcOodWZf2L3jE4sFA9qoEjBq6hl5kVKHw7XdxeNHkKGIQQFAR/lQ8iM87
u8XIGuR+mJw+T8Z/LHIKYly7PDQDJZdPQJcN64X5LEVi0H1+JkF5hlH6UO/q/d3Mve6GeFfpqLW7
ZUrWlTBVRAp4MKOMv0d5Ocnsl2Lwfjkex1E8xl0RtA9Z7AVANBFjS6/aI7SZ5OtFYT9ADbYNF2HN
E9mzx5iI284Wj32cF5b4Nr2qVe9ks89eZBTrkIywB+7ImAkFWTLsaG9KA1NiAaei79wLBkEZZtFJ
UFPfL90OzuB8DEOJp/LUdzlC2uSUeNih5pcQF7P43NFh+KW6qN8UetRAEFo9zueacofZxs788v+F
wckgzCvBG5NbYJV8lkAGczVLc0OAq3vDJ4IRc74IKojf+rDcNsA9WDcaJwWi5hIG3WXMnYEYKDkE
+IjS3Mo1JNDSQycDMjhatYdx2dd5iI7ulrKRLPYphNrnY0fMyLwJCPBHxkgiDVvRHDnVqOKOp8eK
CDUO04EOkLAvZmoqZDhQTzG8l5M/i744TK1wF2xRM9vOSY6lTIqHVLqKFDNMXUXU8Lt0B/hXYjU5
AvIb8zEdPkuW5jaUFetx8VZoYbeWaA4MjpHSxEOTBJsv3q/CWSHZTxt0eVSzcNaBRaJ5Sd8R0gtN
1Ilih1YzZzDwl8uEz0WGxXahn5Uynfh1CL+mZiSn6j6N/Lx6MNS8PvLv/mVxpOpGuiOChhACGZ3e
46Hn5IQd4t2RO4JiNBSsZNjLWeygfwppEhGAIJrq+p3PayB4W9qyyLnrl3BrTxh9KesmwXFKrN3Z
rj8Prelc3JIHhQLKcbi7hVvGAYXUU4WiK2c687NhG1F3rdQK7jbIT3YDhtk9AnwHtEyqFts8Zdfl
lKBvSWRK2Vor53h3bBxdHWAr37YP0wE06Gob6f8Gd89FR757nslxkvZqSygNLqm2qorXr8o2x0NV
v9S1u28Aw85YgvKE5+RCgWjWP8WYkFGa2HnSimeszorwQ6zOsx0eTSn6nByI/1c9rx3vziyPiHCv
piKmfyFQzIskvNKWWB/vBXvAbSW+OLX0S3zEpLQpbyEAKsFr6IuFwy5t6JT7Mn6OVtwnPKegV+qm
Ebuif084sz1iAn5gNgRVIelmnoz24qTa6Za5Scuy+gIoxBi2HkEJX0P0CCvGcJiFC6a4L4OnBmuo
aZy+ZcVnysxV1Ix5ZeRNoo1bzToXgoBXczd2OGo7XmBPBE3gNqqKl/Y3xgowbdLeEYhnt7+Vw+CT
YrBzyc30JdaDW5oVZ05laErTvxwoCKslo9vnnx64suzZuCnup57O7BOpw6I1A5mkX6ciYzi8YShj
C6Alt4QEBPpgH05Ct3ihrnXmGPIV6lykxpGRBaKPxif84HhXLHspk35xFFMHng3YVHIYb6nXUEu8
UFzFzdbkt/8iW7ZE9PNKi9anZpiYLIDlyHkH9EJKn/Ly1mYLor0H6YPYPlfcFCgswzk/oTPaUfLc
FZIWg5ai1BZoYTdYIjocSXhza7Q1r7aWN0dTOOHqAGnJ7Z95ASGCAgXYvW5XZfv8NCnaTkmBpidB
mYK4hNOtwc3v0GmvT+wWDnp+gApDYyEB7uCjTzEFiZyDGJpU8n4426Keysh75uqTu9aPuB6RuheS
khvXrghSPpWcGi7CUQufSnTm39fThIoBx5nzjPg+AVs7VrUixpCfDHFgBjX77aLgUPHMnt9Oblrd
8kzsD04cBWQg+QLcO2OKKN5yETHYYWS0GLe8R4EbDI75WwO82Qii4VR0be0YStq9cdT+9197Zgxj
by3EpJKKHSwPJIenN1ohOJ8H+cEBYLI8qH+DiHXq/eI5ChejoLfdCBkNRCvkQaa0sftUICCyB5Nh
AOzvmHH1SwEufB5g7w8tf2nFGMynkAKA6++mB+63CoS/h3L7xUL66ez1k3NbqwD05DbL/D+cz8dw
rSUZauuvKV/Jdb5GDVkNWl9hayTMCheEFj/6O86VEg8LfWxSptO5vJ8uXvF+fk9WJAJAYmiOMYHD
6iUqrybo/OoJv6SUNwkU9798C9Gf7p2U65DP4nC+hZf23ZuZc6onCNCm/rz8FtGiPes6ItRa9u4U
r+w5597u0J2zPvv+3ya/AuR90J0lH8HeztsIvaSi7T/3hBQOZV18qWOCsijVpKFkRAjhJXgeWK0o
RqV+t10f95QQVRDg28DWn9yGtDijOPAKRIXSp80PSSyBvlU9MktShafiZSJn2r6y7FZTt/CPjX6+
uW8nOgOO6nbw6UVWRA/H00PasmpqGAGZrZe2Oat318MMabLGv1AR0B9bYCjp4QmrR156KrxcUHUk
Ekw5rcsbU95h6vsQLsaEpmc7kZ/LjGRPN5RnfztlFOghCih60N/UoqRJOT2OKbOQ7MYgJsasExBA
V7vI9Aj1LcLAjpY4t9KI93P/qTxInXATBOFxsTcRBUiut9uIe0iDFweIOaavh0ooZ1trJD7TNUjX
7Eeoc+xuxG5jVfSFYbbbt6Pv687vwWmdYPwIiFX/AVn9PLBY4JFQm4BFVTaoG+4su0YlGCaw6rnW
YgFKqZvW34lY+saSriDHUj6VjWTgeCu2yt6WMxih3+NMbPnBV1/E/ImGEZDCCGTyhOmgbHcyKjyV
f37MmUcg6RxXKAFyrWy3UbhBm175nsC2FpAkoPRBOVGJA6XrWQqdfYPn4fp3HLitCyF3RO3MuyyP
+a8ipv+nU0HIG+/L1Bw9SpG2mga4lDPXg1ie3/oL+Mu2/wM+OV+KzRRZbDYSGQEC9CwTgj6tCSB3
DmAiUzBGB2I4f4gESr5oJrnn9PnSUDvqV+ByfrOhXHizso53yFxjboAheS3TxJJELTVhjHMP2dO0
dIFLCbWLJzDT5lrr/XJuh+16oEvqLTn4FgJChOAtof4bibJtAa8qo1hJYunWlqW2gzW3ZygAxLxA
ELY7qa5mnkWPUvwlg5s9gFuRs0aHW6WjEjZmAA5SfgUnCKVAI1qz/t++xY0U/3Co/sNtmyIseXk/
m3uv68kspxHMRH8OWmpc52+1Z78ME09TZ7jvOJamM8985hyv+uDi0y3mD3mP64Z2I7r+jAMrP9+l
VCLQYh0mhcdJ5JQL0/2QGsI01YIZ+k4tE5YJ3WWK+1MHsfk7A46Yk+LlBbPmzDiM8N+bIiPbrErQ
ri2i5uWEmeGKKm2usiQs/KPqqi5HFv2baFFPKKfVFAoa6TpmQzha9q4z+FSZEzYOhOC0x/MlouIc
RP/CizFHWp2jXgpKT9uHop7cZKR0CMpqNEhOeg2sBwboj83Q6YZ/tCYqhp+ATK4fBLwvPKqIpRB2
BItbSGEUAkZI65SR3xWpvIjMPWda9ft/4HzjjCnfC6Bqp0XlyP8Ew90SieFhoGETyP0E+5ZdY7UP
XtKSYyrEX8S3L+s0W3uM1oYJftY0LFMUwKLGwD717Jrip2V+huxtHSUs1jdhq5oMntX/7Dzb0n82
Mjh+Yhp50X0qL+8iLt0BEHj7ORF/GaKuO3sa3oRMbVSE3lEcs4Zkc/fmQxeL8hFTwBcKvzLp65U4
DS2vb0uM63yuBTbY0H6vgmfYkvq2CoH6oZAam9FF72EyjjD8zsYonO2IwNnMgugGcabRuNajK+yu
OxpywsS63D+Y3s2SSOnZDSxwZgVLyztoHeuoU0rOjvLkXyWo92dBtLPN7U/wt42CLOJmNoQiw/xn
Od7haCP7k+8febkl/NsQKgYRofHgcfU2Vz7ryXsOe2VbnasybJx3gZAmnCCRWubImLAvAo9BGJfF
MtN9MNjPiR/u1R9gzNTiDGVaeLqi9jhPvvlstWaoL2pQpaSEHN26TCmiwanfHub9n8HAPk5nm/TN
b6BSltcImjSL3b/HOkEtz1WGMhYbd8hXj4uG+4ZjiYYfDZP27wnVQQ4NI7GYlAIjEDdBb+AudoMq
IqSfLJb5SOmRk7abBoCQg7gwYAZXTg7pSkyB7qeYjVAkJQayXoE5YznMQZO2U2Tnhre2idCazNmT
Cn2p3KolEBLCQ7Op4QLsEcuet/BvjTcsiNDpQUohzXNpvbnWnALmp4qESR9AeHEUjEykN/lF0xgJ
rfqJj6uKLz5qkyHEHb0EwejEYnpjZba45upy+bXbr03MrZFANXRCylhdn2uS5FgSFPkAmnmiiiuY
UyIE0XDraWy0hPpmm1OrI95si9XgdRD9p09bWV9YFS9e0MIAs5DcpkQoJQoXTdk3qGJiE0UMYjOZ
UBvsesdTnh1lCtKh5zutEvNnxRj1itlIM8authvOi5ac1hxYFdnq2n4/i/TZGeNeraN5V2gTddAO
ninaaw2SviV7ie5QE+jVrdLLInGrXtl1Wjxo7Yt/DPAynBUKCACrpnlVW/jN3jJAAOfurC78q/Wr
u0SbgwlMmT00Lui2ZAvo0/fEHK8wZjT5CsX4wbZV1IAjmO05zKjCN1s0EqtMxoFglvfOjzIJZiC0
lcx//mgRKDm24NBG+38McSahUvmF4MIBl1Mhc7u6BdMWSv6X/8cPYLg0jpCzkLRd3mlH5Kyp71Kv
Sx4XVuoK0oWsCim4LQsOt4QCpM646GqiiFTvmQm5mT4uGOuh5Lg4tYRQiot37oSlxC3gsNS/93LN
Hy1gnsJjHGQY2KZ2K/i6dJdLON8MAXkjhiv8e/ar2eW5Yu/Ycnc1uWqma8dU+Ex6bWRmStXP8Eg2
kugCeiBzWMkfY1Iza8ZHXl3NrBmH+ooiLhXPve9e7gF44+QVxDgg7s2PoSY6BNGevowoZFDWuSkI
tOigleE217lTkVCHvmmdjH3wLNpGu8NQo9nYzBHcvfjdKA3K0OWl16sc2C8Bi/kRExaP6pBJywe6
fnmeAGZTuqVu3mcvGmkzeopGtr2zWV0Kab9K5PH2ud4oGjfn6bsIwfxJEFkEZB6X19raJCQhpdKC
X4Lo96PpqGilW7Nt9YMOXk+kIfMR+bj2ju4jTlQ1H2DgoUSZlJaJaVKGI4i/q/Wt1kBzKuvEdTR1
ys4O3Haj7wZpE4z/Sftfk519HWVLFUcpEIIk4zbGFUz1LVu++xAG/K+2ivU680knMuQxnFUZubbN
XpJshcfESjoFDeoRmumw3ixk8an/j4OrpY5dSz+DfGq+d91jkK13jgcPcA7sKptHDcZ+GVoccU3Y
h0ojX6PduKK/l3C9+o7GcN1GFQn8jlMHxwwa6QCw6iuYsmb8/0V3LXTbD2aWQ4GXAjNFfxurXdmD
BsCMtJP8YXpwBgDSoO91SZ6bJMItDDGKSWvuoMmWuAQoCRavjw29BxK1b4UVdStcrJnRQ/H4ckhN
eDrxDJpFyJaj6DQOHdCuY36/jsKP5fLrIvFwjX2mlxGqerKRbslsOWUqM+1rXgdgSZ4nJizY35KG
kZFTpTW1QHM57rTcIzCarEvhYwhu9T9F2GnEZESPRpYhnwLp9mbmYvD6IgFnq+aFsZhUgag4hPSW
Ohkbix51C1kUPkfpcQ7Qlbnvinm+4Uj5xCM1cDZjjYwFdILv+mMOJAtelbZjJZV/9iTV+2B18av2
Kz9c3a5t5r4O0wgd3GGgIxl5fRg6bgUpj1srI3zGz7PK1hbruntHs49AfhDB4HVkRuzmTmiXnmYd
OqyPY2OG6oUkqrI8SHqZOlZIfJzdCJT+rw8Kr+LnBFXHcYGCyHbauh1pccxUeivpVK1J3vVnqDuT
67U0UPC/vj8/QcfOKgFTuleefcPWyHtPuq8L9Vc3YV/LtZYGx9nHm5R6Lrwty/OPCAM2a48sLH91
fMZ8x3JUtS5XaS3z9xDXQlaxUXG2rsFnPoa6ZklT2Q7iWG1djg+Fc6FmeojfVJ7JGD2ylx0Uo3Nh
mwmuPTq6AuG2ALktX27aO0q6DsZZfjBY0DiNxSLjaw2m/b5+kxuHHmX6US53XmM4vTl/ocxymXFb
FitubERPR0VTsUcbjWB82ib/oklkPmn2NETPjvXp3lWHijQfv/4s6q7Yx6BpfLLGsW5bpHuQY2ur
YJyG7ygZB8uc1eoXtVnt3S89T0YceO9yKrf6NIYu3pQ+PfzKRQE3Nfrb03XjlU895tkbWEwC1/Qi
OEFuuot7ikKE0ksJHNGlnIRt3GvzuH318bXvWkOasXSvihZlThsPwOPmrjwY8bVUtlgDVELxHKHx
J/gpen7hW57QCCLO0QRDcG8ZLkmwMxjYom6rYh47yfUj6qdM4sA20XTL3W5J1D++pD9BpIZuK2et
A15YmK7zTOd8utyhBDxULnG0W1zU0oDRx7FhHVsqPeTEk74WPYiBoI0Qpz8MCyghGzoLBE7o7VMp
dPspLIsApNRmr5VbYwuiKLEKWKytoaelCfshmzJIlYKllaTckYEobCX/1r0+MLPSpkqDD4mLLetH
VFX2dOHk0J7PrdMNW8TDWKgDsRN0vwxOBwGT1fTS8poHmRyunnmA/rjKTzJ+pzCNpLUzHV/yDmMh
qozVCP0M93mr0c04x7c3g6oGs1y/YHUSxwoTjwPF7+VwPbj0eFnhqubni0wz687aVpHHpxdPmaAd
/TqGjj1spV5zrgph7TRzUOQFh4lidr5yJs1q78NjKewiZbgVdJcXQp/WOoQ4Msz4/9z/k51pJjbs
S+cBpvN34MHALJAL/H/59wtyScmao3bQJln2rbFGkLK8mxfvZ7NhvoAuTps6kyF/wUBn+tu/ep17
m0rYago2PV2tzEtSyGBSq7HtGP+wLlL82VlTB+U7KhLz45qv4BdIcsS5aREzg6bontyn0qjjX7IT
iM10TXakoZeibYxE4XpDr4boLTosRQ8bMtrv7pGRop8/XjZRMrOGxAaCjrebn949UVOOlAtz1yis
QJL2ueeMPfFDrt60C9uepm1BVExhQCjOOfEgkCRYZGWuJedIb1b8R+DkRho0SnCmUGGGtG0WbCp7
YQy0SBclepfwBAg1OChLAPYJ1J0PkXZocBGhviDVGnP0hD+Za2/WXCFcc3X7iPubNREOtjzNwf7W
wfvyswNfXB+ErFpVrkd0u/yc1a2ZOOuU/TUMC4H8jaF3qgRu2HxcUVxeRvjWMPOYAdRNXT4WJfUD
EwOPePxZ0q1MBYEoHwoLYcYoIy66VU/mBQUbnAUMmGxEtlspfSn3qp1w9ahBWyk6KvkSxIt3Uede
XjrtH0UgvtGVWyBV0h5qKwlKbiIgqUFZenI9nh6KzIbvQjS4E1rg05OjOlJW20JzoCqAow95kEeL
6oY0ywm/dGjqOxGGm3QvimzOlJmapKmB4WhRCHcjvZrUovXkdljHys+Z/ormy/R9IyUo30LzFO3r
oq2OZvfPL9d8mOrm/WCMkaxdON97bDwvQ3AeOnKLEYp4VVqZPVpYx26yoFNa0hxR0pSi6UHvsWxO
yav/IKdGZBG+2U81vmzgsjkv2rSCwq/FcJ3PaBhEtRpGHtvgK+FwnU/ousqJscnrs618QMlXmiFy
jo1jYP12tY9GsusGxQXcQupgTrUvEGOoko5iUewayyIJBpyXgemjXOVNUtlLZGReoOIty1gv0DLl
pK5BQr9cBGXenF7cphv2DWv3rSuocY6lp4moYy8WcxABYggAerxrQy8A4u46Z8365RUyjSH00YI6
Kh3RxmLYhxdtyoWixKpp1jpw1FVpTBYyPEcCayXMgVxuGk/b4FEj9/zKbkvkgX2VqHWqhPxVx5XE
vZdUDJ7HOl8+uSdvJGykFweBGNCE9f7ANVcZVuDF9v/V7VAyVi8e55LN8iwwkITi5SvviP9tMZxw
D5CX1DwOGeKAvlpB6CrKD2wcTegHB/rKx9dd+gDHtpHutxNKOl5RhIvi179Ghmijdjj1+uyzkHgb
KSLA1yaj2+4G/SCYeUDxrnK3S9RPxZZO5AY9Vxi+olJhvXmhbaX3zlWynozKXrM6J8zs9HPNm9Ag
k2gM5Ku5qQRmcHD9O6TLl+8M/ikGX2BfNpMd0mdYCM1L/8GdJvjfjhPpubeD7r2C/kn57xz4KEYf
nhLcA6VTVBF3Tsg7LLSCtgkhccFg6Bop5M3wGJlL6Q8IpxPPNwUB8jogYiMPY+ENtoZe1m6o01YA
waYjUNPf5p+hdqV1JOKWFT0a1EHMLKIvcMpu/d0WZfTHDKOL3Jxwez9Pteq+n5bh83VizUkyR3y3
TZaiAXaUs33OVtKGwKs5MilYMEce0GqMgWUuiSTgF0aELn6C2sdrPZIfwesdo/vljDbQSTbsrlNQ
Vwamr32R5H2BtI2vluzkb20VN3FQ3BJb+g7qswo3+ejXnyXRIqJ+Tc/IO9SqrD8F0U5ouYWUioZs
JO4DBNF65u/BcNj7dqhP+ONKYf5f2nkfX7Zx0GH9LCiPv/mZwc/pO5EjCLe0YLT37/wS9xAgHTpC
EvcjEBZo1k8e/puKE3X8Zde+sFy3tqYHtxVmyDjVxA5q0s8AO6sto8yB/JwPxEUyyRQjs03DwVG1
njb8PkHked1AsnWbXn3gFlHp6tzsThl7ohIyFb6q18b2sGoXXTcuWXku/UZw+rgPa+O8kvVIvGFg
yiWWFT3Vs6If5+EKU8FTctt7tFGLrA+eJyLYUQiN3YLeGYYITz6TFZsqmEi1VxD54JXx4Bhsk6Xb
m75PbiRSov7p+0teFtbLHf3KxLZpLR1fQ/GNZVZum4gtlIjkuP77Olvw2CHvr+NvlZ0QKry1waRm
caSDrFX1SBUFEXQrq9sTH6nSrUU5Urhr3/1U+WqOWlxU0oPg2d3Cfv/TnwSS3I18IJuydtlcsSB9
TRAoC9ZcGJtvoD3lcDXQyPAmEnjecE07eiDfN1uerQFLIHIC2az21kdLYg3a3orNwLVmEmTdvkLq
8E18Am65OP40Ym21gRrcU8CkLpSzeDT58KhnVJa+Uf+d52yx4BdKSWqZEPCsxbn5ncJm44SZYHUE
PHtvWIQDS0EoGmlm+PPY8nMWwL4sajkJm8GwzMJIyk/gXYdz/fyFvPScHcwzszqxYToSOlFwmHM4
LGPTNQJWOkLpDiXXZU8FOZWVeXQdrGiGJs0bZ2ODXocxlEb7YDq/arBHU9zD+zjm4k37+Slf4EtD
bhxMWF/eJdPqFXyLMdVv4Yk6AmAh4ybsmFJnEFwm8MPHlwMpn9O4K57ruEk3onR9xpyFrMZ3KMjH
ImuK8DSfgrXPQoe5KKM84neKU/ECm5+pfvVYQWZpxDmBdyOGj0p3gCRy5ky06HMRhWtdqPETlcK7
d5TBUS4AG+NQRPjzG8j+CVzhzRSVg1mofFyEh4wrqCaEr7/xHnwP/pCzei2CEJ8vC9xY+QiWvlDW
dm6AGo4m/+lMTwmknmitiJxldXx7KFcwVz6Nym8cA6wHa1/n/O1jHs+qQ7YeLrwm0rdOcj0UpYUq
hN46ZeVisiy5I1kytu0XowVWUkV1g+LXHb/YjR/fkaieEPRCvoi4rrIQyMmZkWy01KSs4Jl3u8tC
hwN4CLtSMdg3jh9SyEpVvBHPg7z3vs0hYsfH7+QUTZRLJwgiKnTkuFEipqUWS3TGDDp+olmDcxfm
bjK2uJewH0D3DHdPdg9G9P4/3DHkWuHyCwD0Hc5eeGm4vzkxInqcORsjh5Ho0HZazktisE8ey6zX
p6NHI2gJAWUhlMKDCLi6R35pr4YxXNbCgAOWUgv7E8IOXmVbp4otKloYWI77Vx2tBLR0BJGj5f/8
etfEgxS0xuqu2kZSk4LDE/1dauJbax9FuWc4yQOJmZKogaPZpVRhs1tOeNKabxv/CAsFaVoqAcfq
zeLIzm4Dgc5Bu8BMkhq+sUPnRZYHEOV4P9eimwVzYUrhtnud34aUclkO6LbjDrmRN/JJ+3Wl3E2l
0TP1FW+px9294woOHmAhlYIWMBkDKSkLHaWfwV4Wuh3r1rYHJ7A+qflZgFfuNxqa24Mi4lRrAZhh
PjSNCwHUgJCIBiUi6V5z9YmRa3ufNFtx36vFJEtBMIB1Zb7cfjdZdTmccxYWFAtJtbxf58WQoQeZ
r80vQUHMOI4iZzDZ6fGVpnXJIuMfouFFvXMbdxRoXPQXrpjsuU4PRr05VQTlqpwO271AbyYzT3O+
I7K/DCstw9W5gCXsuD6Bx5XUX0OP49kfxnozdbXi4nxxHDr8vWiGbynalbtYuYQVJOo0yeKhVDln
WUnjdfG9i/J/LEW2gFeeLhPjFTXUjmUt4/B12YWZuL5XR+RdcHNVJs9hqLKKVtWEQhKIvD6kMh3S
PAcX67NewDr0uJWvv40fJmFrXjHH6fL4grSqQ0PF0rDtczn4Sv6/3+SBQNSF9tXvE20mtKsKy4nH
oklEuqPobv5nFV3jW49R2KHZK7JkHILfUPeIB1yUalWP3qSY5Zfd669nZsnehfmKR1ec8/2xLo3/
ZVShNiemZdszUKBVi6M2nEuXnBOwZxoqJl0ARePIeJWg+2anddRSsCtJ/j4vi5fA4QHban+aEDbD
TqQvDyYQQy3kF6c7G3jQTXCLHKK8Vta8gx2mpVrdLwGIn/uwkFFehWIygLr9zYbFKUn0h43D+cQO
2zK5ALXwpO/s75U2BGUQMdFh0F5+Zw/BXb2zPSzF5rRJqLkozoDtSlEE8Og4S7kl2+eYcnUKUDcD
R6GGeAmoI/tiri4VVFFHvWBc64X4yzQgmdkI7kQ9iTHLEXH6CqGN5uBrtDBwxNebcKfz3moOOTtD
L2cVaKrhZABz8iA0UxD2VIe2qz53sHsYjvctb/WiZEWjyoVXXs9fx0A1jvmaTPcfhI+ZlZ9mPu0K
2f3FKvLomX27IMUu8Xq2UzMUIFqlnTFzJZ5hGV1fmLBJ6JnvDYrmogaX87kHmeYCXOX/TOnS1LKe
z2roC1xyd/4bcO3TsqYpzIWdBNapF/nq82Pm1vs6OnI7UDkMXimeSoHsDAnqlQIu8IvfUjsm8KKb
SQjAzQOShZznZwyUrqHC4HzMyDq4Vojop3yHAnjfiIej04uEhJTWOuR0N0p2U/ByzM6sCzsyImWo
fccvQ4BdiBZ7qfTRPdZOmil+pOiLDS47xu6gTdXZJDqn0EIApLbX94FyOZZwD7F3E+YuVlDeP4N8
rKGfCVT3kyE8e7IFReIeG6qu5ReylLDWop5u4mTXk8vCZ2k8cBxchGSXz/1BV0O5qFZLJKSRxZu5
83A1k9J78FCXK4aGxj9t0Xftv7wiLaBtpUQj1kMB9uX96NpWrE2S62ZblPeuJjetsf/Gb//UKBbc
y7pWMM0LS7FtbAfOeXwzfpzTDWHZo3uOWUJWK8phnIFToBbBliJJ+l6v5I6lLL5SnjMH6wVVP/jC
YYwb9M91Ws/9ZDyzRzEflWcNsr6/n4pQet/zRkomb8yg8JY4R6/RDJhCy+9TKEjdpN6NI/gxpUgF
33n+ZDWq5qmB7Y8fI9TyiB2UMA+CevVwXaxJfU4kp3dSLHJu4DylHNFs2TpKqWsSX+ZV3YUXH+cJ
x3/eBkW72t6mkAd7WUl9AqtnXoqrvUZD8eAje2NnVMuza2xye6MmZSjeNMvlUxljqcXT9TomqU0H
6VCcP57JslaqVzktWpdg2ElC961hXsjpyy7NnA7JKCDW58O+mz5FERCVpQZ9HlvLLpE6d7AlOtR2
R6+dUWVexABKfq85Ne3b+/Tw5D9ANV0aFJ86ft1349TLdU15RVxWFxHY3LnkQFf6kJGiITNOy1W7
JJse595oeQ/Pev6UNFkQLywb5jU4xWgI3r4J8+6lpE7pMq90SBObKGHmDigOTJvpM7/o8VYCBgjU
vOtMdUJJpEDZbPO4PZSjVgQ7L+OaKJEUJw24WC7SU5Wgha1FJ4gDwrM8lAWENty8KDOWbzeTgPDy
LeqNikIO9LK99PAd/UVVfrv9LiXT8RmBMJdDw+lwlF8Y2eksQDMgN9/eX8fMojDryl//E20ujpK1
pY5i73avzbpVjGZ4nnVZzlK0FoBKWZiXq86wKD89CH5GPtQD2Xpnm6tIwuAyjcX7zwHIx5O5BbDk
hvMqurBO+9/k1pG5pZe9ZbT20mGF9IvUoOtIyvEWuPqrLKXVl5w+325N17ds/Xxg/xwwEpiGUAbn
rcvLTky+yK6H8W/3oGVgeibA6YJJCCFHGCm9LQVMprBCcFbQ0WbInOxu4AjRKv7Dya10PQY9cBtY
1sk07lO1/aJwBsxJmcj/WmUcebiZLDH2TSyWC/x7zwr0A3uxWUsn3ZjQsGh/jb3PXroahG5f9L0A
Tx4HYKRbJV3kpaW9tDWGS3o5gZnO1u/yqI5mpSAWcQGQO1XWKQ4Hstm9ZueCpHZFMpnUiyGTlA0B
QC/HDN/AF7SDHl+JlhJcqUV9WolS15pHthFzb7m7qGFOqS+tuM+/rA4udWKeU86PA7szUN5qZTXk
1da0HAHUSYFm6HOa3yf2IcL51yMT+WKPoZc/Y6HKZHU4W7CtgH7MrvIwu/QJjYOM9d98J7QTUdmv
xR63zxWQek2RraGuCjzpqH4ugUJZ7/Plkz9VlpmDncI905LRPqEO6LAaHOcDS8JtGqaFxRs4L2Kk
iNayHjvu8VuedM5B4CFcDYvIkxKoVqTCiU+Ed2i/EQHkq0Dd9xBX9CWbV7rAQSGs/MzxW/6Kq7Io
bfgEyPi7KcuZ+mjPfSbHlS1Q8Kn5cPph29dn3UB2cHizo4M1n5jUtQHTc5t0AKwbwhly4TOvyrZV
8wfpoZqF+ISGrgGPHvwPgBppfnAqZW9KiT1XXvHJJ5Wd1QuBcOsm6atrXYxF+OcfbXM0yObAh1dY
FxQOvXdzU7LKwzIL6WOUkR9Ig0N7irLp1nhaFNKgsjmk3x9VAFQ5w8mayDogaNKzns4asENlM4+A
VHizmKcNa1G23Hljxmu9wq6yvaGf6PvMEutdpJc/GaVg13QIG6L5Xw9uqzTrrRSOBYw1w6gy+GJ3
zXvs+iPwBSjSw5jqxKYoWyPeYDiG8aZpJkZcW3sMIL/FDjssGZhb49jQUJtBeyn3sLT0O6vFJAIi
3YIR+JccycuZc6zW6HZVMeNo2FFGYB/HpTYwIPZQnoX6RazgfVR6jMTZZIAQGVnXNewVg30qa/fb
ErBMWBGI+5J+rkQKa3bsTrpxemcgrpFmbXp5BjW7AowXVEarXva/guNrB2tqikTpdKenqmQ/ARPh
tL+FTFdH++b8EZ92HBz8bNzJJw2SqD2hSGvzwHygMoYSyGBgJvbq57vK4uUeYY1Sh6o6aSS2nZkK
4FmIzBR3Nd21K3bO/ujmug+d3ULO6n2DxT/RecVAlDnBJ38CswpFfywFYZwQX48hA9eRCw9QMWeq
gmIopHpj8KGu+ksxbdO+CFWHIVOLn1tzmlKcXLYCLwoQyWt1B1fXf/axjCeITcyMmq6KoZkkBcWr
k+A0mD+GGisPG2/Q22oib0yp1qntDZmEgzSuvl69KIaKpnevgmoon+R8M+DOZ1E7xS8Lc/L/xV75
LsmVP3GmIRmJre5sKvMo5/Tfhsq9nNMSkMi3SEXoF3AZcmDtV9vPDF1tb2rpTIMAUbs1vFN4eDkz
/vkqZYy/6L/uWAoxFKJAAVol1TiLU8q+W3M84/R2V9is5pIdAAj+TAnSJ3f0E02LfyAUnnmzHLlB
g+0H/gT8UPxznmuJqRjrTl9SWhbZw/I3Wxe/2mRnVuKSg/hzXoHuXk1krWOrNM/Tg9sTRCabtJhR
4QY0KYHenBWEluyO5JF/qNxdFsgDoenaHUsXT/ChRHrIxpSI0OmL80cS1upQnV8YwT/cQZSJR85X
KvoWbMGiM/zM0hLKNsiojyonkBAMoh2yr8NiGaAOcWmANDZ5mS93SxIdJOA3IQvow0cKd0NMyCzZ
4ZVXUaxTFcVVEYDJgqyUKvOz9+IP5zZ14uimNNHMIMF7TIo0PjQ2l0g9NMqKBUQgV1xYlDq6354n
lCaHDHwg7a+m8OPRbPqFIZ0weBc+wQy9IY5AR7oUhfU9AXDxA4B/i+UK7Qh8koz2q2DRZxKQ/hFc
jMvV/tfjGYfcbccsSAKoFxc1TRfJnTIpBvSX7IcB24uNJin9cEX1tC7L/xOYqYfaTAQGmOxxtkEi
2ODUqsTKNoVKwhEeJ34EloqkqQCWQZHr0TE4Q0wct7xkVHfmF6Um2tMjEuDdAKLghJO/tk2Nw36A
k0kPKqtLiwu7swnCEP4vRdS+bWh7hx3NkKfmqsHU+iRIuZsT+lrWLao8xqzB6oZLyJVeI9RADgdn
P3pmCcv2rv0RWMVTPSd98xrHFhZssNAajadX2ZXl8WF5xDjgd+dN0GPvGWSO10/XfuBzkSYCnIjs
CUdrgHzYrcHIRv5GZR+PJIGV8oAt9mGiyS/YRG2IzcOMQyytnBvs3xARsrK0IUX6dOtfQCTjGqSJ
ftO2PqzkeKD5NpDMu+St0zRiSwRsneToalq9uTyN0c8nnfm8RcJP9DnEGLJhLcd9v5qg9Yq9XzPR
PJll3nr+mOAmjf82ayXGHEBTdg0sh6MXK6Bcw/H08ruTEb/u8EhdLI7YJ1u4JSx4gC/vkD2mJckn
8H+L5SO2bjrmmiThwV4w3nOd4i4WcCLelGtiizj+ru2jixYdloEo1fcz0w0MVTBLm90n8mWxjs6x
MBv3n+fE7dXGQpEJ9dn9fA0BmTgHn+aC1h8QLpFb4Iug7gYzjAwgixQ2uqRkUss23ApjGB7bxLMj
WJEvuBvR9RazdkyNrdAhmSRpmcEKkFlt+j6zNK/98T2rKCr4tpJWMP+6BL9sEkJXhpNDm4hQrCF4
qxdllqMMGyUh4EAXRI63sBg0O1fI6rOd5BPFoC0zni3pyVZBUooUk3Lt27LYunXYTORnB18fUXKv
04naLysw3l+fRoFUcPCtkfGnXMi1z0p64a0LzxcUkQKq9AY8fljNel8Dy4EzkMNcGDYLJk512IV5
a6BYEDILkFUpl3Fgu63otHZDRy62cD5uBbs0GtMcO4ixydtkemFKSN0vkRFq+F4oKeriYia4NsUg
B/7Ei8zWvP/pUJ+Yow7/0IyJFWEugZ9wYhk3zVg28PtoqmTfCvyQdXVapCiEAEqm/SmBAQqS82Ai
bTtxCKR9B+IdUK3Ez5tXtWd0IuO8qR2kGXOduhiGFRx7yONS0vPIwPbdiMk6iGCMr40LCQ8QPDjv
2ljJdZfwChn4sJ1ePm+Fm2smlSyrfA9R3jtAM4d6d757EXwD6OfRu0beWySlpOUF6vPdObhoBRSH
rvfePxSHmVAqsYKXoT8hDGPcaZAcVy/MrHbTKI/510YiSNr3c5UWDIpyOLSgqUmFydSLUzrbr8mt
e6JpltreqmyooUVE0cyimKAdUEU61hD4LsvUTuaxAN18W++aehYxxDTYMx9KO/LOTpdsndOR81WF
mVzrPK41LUJeFZWaK4Zf22DbCPmIMOebrlq15bZZ6shA/1v7mwTecZyTxdCGhmLXbS8m9ikLScy8
v5DMsCvtt+SiJM/zLIFapz0Y0nAVOX4ddYqkya2LlGQTXCbYrNv6RA8Xpjb+lveUeee/Zcn0kOSX
/C16UxzMSEfN0YckaiJifP0Dn1xn8vr1N5hSVD5p8hKJ3D0fWPh36a3+eIsEZK23wn6VKFbbpzVy
76GLGAKk7HTS0/ZViq5sI0rI3s6+EPvNm4l9N+U+Tpp1e0wI+8NjC+NwA8eQ/QDoWiCMWQC9Y54m
54WxnmqyFeA0jAuMhRKPpCvCuf534DeV1ZnpktNf7+XYrnvUHQ0QK7rYYKqKdwXk63XuZof6Ulj5
Nao2iKArBWJl9QrMRxF7lfY3YZbemijQttsqInMGPgpNob3eDbRbzdgbkuc2iVCcBvdUAsM2v2iY
YDHgap9UTuw+/2pzfggrhEciGd4AWe+uJ8djQb8IcvaX4QWF5o0DzMiN8YkAerfB4PIy8mzVWIhF
brV3E1S17j8ZmkQsGywk8hhal+bxns8euMwkXi1mano+P0dta13gGu8a6IIr1yv3bT7SanpDOkrs
26NR8gmHEnDeNKeMQZXg7PR9yRdEdECrN4iRmGbef9fV7UnW/Ni4P3+sdGeKnFRa/uXmKQ6ph+UP
seRmizWVy+tab6C58NDOL35xL9wP7uizBKnbrbV5ctfz0xX8XLo4o3rk6uP5FOPFjLUg3mzLhNXP
MgOeb5p7DQpZcc/E+zvM0yLfIBx/N+Q59zLpOzjxm+8lRbNuWh/Qiy0se/lQJC3C37eAw3zAHfbD
3o0Jg+ww2/kmGxRPXpuP+++9hM31X4EmK755nafnG6d71vLr02hoy+ckc8HCtFX/SfccoOdnUwNQ
JluMAR2JyEN9Lxt5P3EBPVztyjUL6g0vwbwVRUBVF60trgCxo5+Q4qYCs8T5aMqRQnBfQeQAoqXN
kn5n8Ahs0YXZqulzClFuw8rDh9CHSq5YPF4LTyAl+cFxFUjVcuM7Dh7Vqd/W6yrV+/xlCQ6CwN2S
M2J/crBTFYKA8uRSnkNheA1IQj85bS++Bmc9n5gpxtdwGjNrWVap/GBwPYjXkevOikkqWTWPtUtD
hNhC6Tbvn9rL9pect7wJ/kZAZzYofYN4L98+JERElV5dx1T7YtB+NF14NjF1RNBmM7qjLlZGFdGQ
Avo159Im5eImpNTRmtQYTVOSZfjPa3CI36JQ1bwFPGH3gcLOqopLtTDVWGJ2sPuXMChZbw6MSYNB
ngIjY87DGDIx+47EHnxebfizoZngOwZsjH4BDQZLGFAG/Mpl9CJHUtfG+4dmFlCv0t04GO+Xg24g
O99YuREpFLEzbqrAsEeGqs//M02eU6Fhtddo/FQZjkVjQAbumluk21dO+yJWEzxIOlGT0euviXyX
6lggJpEqSUU2vT+MqpwZpHyggWS6w6YtIsTAp8GH6JavvuT0XFxkkOUDCWMcpffj6s47aKb3dwC7
P1mUlpC8QW54NO6lClD73X6wjAA4uWNJ4LkJQEuVidLi/gBVKc4zKZra9vYWQxPQxVLTO+4KninS
5osF4mf7QjhuduhH4q8Y7DlRyb63rjQfmpVyBf8+/9rllnHRvemgD93DSnUMHYRdIBEHwHbuDL/z
SrPr/ra4cIkOWW5KEfjxVVlgw3FBqY5mp0FViczPiQ2S+e4xsYGYAkgZU0lfSXN37YjFfblZV5ws
FZ02m6oV2bocCiG36wojtWwglFDCs3QSW2Zmi+RTaPEuO6NioM33j4QpWQ6sGRq+WFQQF3rXiI4Z
ClwwB/IrSyS2Dm01wCjolF8Za2V2G9S2Yjg1RShS/fbr93RAYaoDfTzqbyVph3qhPC+UKo/dKqBB
t50hXYQ8zlyoBM4r6zqhX7xo/qSHr/biaHHohc765vjb8Pl/QJqDnCZEFfKIaJl89fCdBEPsmGDv
hFU70aR9xkK3elZam4RnhMn3t3J4kD9eoAXk5jvsDxMGm4HyRh6WqwynZiqYka9eUwvAlmpAA3Ao
BytIRln+TuTwXEdCKSdi4HENfN3qBcfQxj2WIYZxxtg0caPyJJ4KVBsFrJ/E/bdg2p2blqPzvRRw
RcL0r5zQ8j4O83U7lsqhoPRrUg8HTd5Bnfc7bDuixVxX/+XcyVPXBqUyIUbSY+fWajg0GN5fWwPG
E/OQbA6bxnWLL/AKhbLTk06nDHq1TyQMSguXeJ3agV5OCCEmSKj3mcdb+ESFBdmGNY6qJeeG2Foa
0frwMLt4/kOGD1hFrAdnu5vEGlNYjxTamdySqplcnRO28S/6V68rLbFyZ5KgdDKFyKEBbx55CeuY
2H2DjyNsZz+BPj0NbXRdfyxVPnwCXg5166zqV2k2Wd/ZYBKV4HwMa/4q+xTsEn03BngYY1g5R/f3
iYMeZI3PUJ9tiDiB5RWUjK69Ocu9ylKh/sv8U9wC69q74gVlKniojRy+MQ2sstLkr4MIkGGebYU1
PMM4iL9ptfRk/hKsXum+12/gkwJcvUP1gv+YSoxewjj2LgZQmkbl+sjTSF6oE0A0XoSmEDW56F6T
zH0yOY68EzaEu+YZS7su452WdAgGuGxs8TnI87yTlHr9iC9g18eYwkGodtJ3r4x1D3/t1FrQoAfY
akvtjJFGKjK6zLDv5XjUS/2BO731piIgfbgBMRP9GoCrJHuWqZfzhtCfdpaz91OoWLU2IskQb/Pl
giY1b1cqYsZ2wkoQEbNwhLhNhYarzzJgt9TfngLH4SZUdWV0uw6iVXF4vjewQdLxOpuyw00KO9w8
TB4QL+Y+9qXXZpkXHVT44gX+LEEWZwTGIjrcaowWuNEnD21iRRQrDhMVYeHksab+mDk9wnNsadi2
jrmHuiYcD5DA++fNS9j1v4Rvqo73rxIeI6QC+Y30S40oAc5TVGWojZsb+lg/UA5qav6mV+AusM2w
hco6zBfdXLh5Wpc1h+mRnRyp55OJGfzjYOpJEQmbRN6qSBmFDtMFRVAoy62uigoAdxmRyo96Hy+g
cJ6hvdI7FCSx6erzLxo/aPZ8zKljcCrW0BPUI6tWMvmpRs/AECIS2jfKcO2sm73kM8gpuaY/BgOf
/J25CBNdHHQlFF+1lemuKaGK0WtGYq5TU7BZJmWkYzkSXKLqEU6/x6+B8oXMQUnEXMRmwnSfWLCL
gKIw1N66uh6kPJxGmyhgz+8kwXaUKKQRTIzoZPzjOzO4kvnFAmZ5RONR8LJ3yfLq3WiwlXB/wran
LtKHE70Vm315hbHUqG2AK6DY65wo8gxFpc4lsmzRVCDjyNBtNIn5oYM39LBesu0jQ+vunIV/KcV9
sn6HXE994GZfappCiSGciL+l6McIl56Vjyqeh5Rln6url0nhyWjxPcl1zF7JN44ECaYxOWi9bY1I
K/j4ViALo3Q5o5slCfYaDTYHM4+SaFTFCxEwQTIHFZQ9A60e/S5SMfNStD6Fp/s+i+7lqpFVHTQu
/7uR2QeBI4xaWtJgpFEII5zVqKysbhepyy4VRxODGVQleAcE3/Z9wtwuiWWFQepldcXQpaH2KmRp
Z/MXMy0Hhk9nQski+utY5pzwB4J9TtXrIH3BXVAo8t6p9Q8VEP7MJYhxOYTEloH8grbgAFqoSKOd
SnIfTmoR3FUfMV6ixXfyEA4mA3c88V6/ZGjKOI94UHKMhC7HY+vCG907leDZde1KYJVeLPndG53L
t35ucKkWawWr66aJj15TgK0fhjWvMWF6qcCsOnjNbyWYezuyK0h5D74SqrsKlBu6YRwP8yIuBsyB
GDHp3A4q0tRPjPQIMdMpPUuP6knytHccOeUyhXa3C5FBl3A70RkFkVDqYN67l/6BCLU+iyy6ARrG
WcwfxAZcRiWO1txxehHMYrc4WZ8sYE63Ot/5YvWviPQxofo3+21DNUHeM7+szveXapXDm+TgSktA
m3f+nOzH/kCDiZ/tDRGHEg74voYJxZtTfXYQqncDnJY1y5Qa8K274VH8krpCDYkSYgSzLG9wBSBa
t0lxWdaUdHlHvTSJJwF00WcnhkOIaRdOqYPbugiYKBpdFJi+g0W31A0WGsYTLVl0j7LyTSinzSFE
vyRDbj0wrbtj9yQLs0wa7wxga0+K6t/l12zZ3HcWfmYafhoTtg/+ltO+fNkVWU9uFT6sfsUo7yco
J3xKE1E1/hix4nwF3qQKd7Jf+e8R3kjlCVm1MsBJnu2eadzT8RzispViIPXg4n2lUgmxl2W/UijP
LRXgFBvxuax7bZvb2L5NeZDgM4o7MrMZMneiqO0dwSAi+2fD0CogU2zE+q6YXEZUy1HzKD/DfYzA
5iHv1C+pTKvUEcLWsLzuU5EMNOVL9/jWvliUQqqF7eiQlE00SEMLcN3RzK1+BwJDbvjW0AwUhjcS
zhL6bENPy7M+Lcf/3KeBRbze2Z5qZ+Z5ql+DxgAzlreP0ySSUal2BOxdGnWBDovNuIB3DXsm5R/g
HBdJdYn+jMP/9qNl/rZJ1HmlI7A4toODVA6w86nWYj0RyPwV2lXPJPIvyXUQRSUGqoC9az+NFemA
Ah7KUhnhl+QCZ6kztZ95blr3SrbnsatwnegBA6fsOomEvleF7gA2dUZVC5LG7Ab3iQn4l7C2BI1T
njW/WBh3kTRwqa9IinXT78jnT0AekwD3yqTBj7W+TDSOG6Pule6c8TyMyW/3QG0M4MVm17I9NjWW
nBFwwNnJI7f1W2No20A2shu0HCTiDSSR+OaFkcI7iOGIqO/SVGObBS22m1jtiyroTmKLOBnXBHce
sngeq1ZwRXTtMg+E/Es55IkWTdQW9W485pijA97O/1EW/W1FSOoEfhP8LCPzZ8n1ecgV70ETrmqd
keMobjZes+XjuL9hxP8Rw5a5T/MJRW6FGF8SbsmxWC4xyYDPsDu34YkP9p4eyZV6slGO5gVHcUhE
LhzY/DsBcuxHmAApf0yNwW2S9uJkUL5DpMnpIdzyabloUM+MsEp4stqAcOyzRU4/CJAr/EzYNk3D
cdp8T4Y/6Gt5aeZ4QG+6CidJ8q3dyWJ0aLPyZ3ADHA+2ZrFGN/Gu3hxL0RHRrjaAf3Q2zNhvgxSE
Jj634Y5isCBq6ler+dPFpmMrVYnSu/bPEozMPih8SBQGgIRjPvfL3rOvsn3nZFmGRB7ErKD6aA1N
MWkrXDEXsl0KZKoO0LCG8unDSk3jkoF/AGUz+aye9nFYz8uAWf9zVaQHLS4vlar8yp7keNfX1TuC
aF+76JfvpQiGepJc1MyjrcK2pvxVN0JOFhPcYUcni1/pQ3Ew5aEiyQfi0r0a+t3xmHOW7dG7YyWQ
i2dPj39gJSbfEESt7bslWVq6j60imBE1JA4ChT+oM+bar092mOm8cObSax/lnM55aHGfNFCa98Bz
20o1uiEpEXdngKTpqn/09JFEo/TfKVrTMwHQZx45nVmOP1quBDL5y7p3n/AYRcACg25GgIqRc0Pf
h34efDwj4QRqa2fI88V9ZaklE1pVu7CyIe2P1QbeMcBKGyTTuzURnIK83cDd0O9Qfq1a52qi/JjU
ydzs7ELYZphmjsRnnCkxdyKvxhklOAGviVjcF/PSYu0T2O8430AhB9xlr6HpuQh4413jZ4QBVMUW
9QQPGBZxoE0iAy/Cn8b9JLaE/Xkr3tIxUfBpIbPWVkTRJzpsnomSbnQwI031zKuRCVlS9C/szI+X
WFy2NKDlc5erh9JsnMKLKaE+FgKenXmXc9R27jFT7jExVaflH9eOSVorKcAH8pZJU5qYeGXP7A4w
ormAkDQhUvlJmSFdmoDPq6+8i2EJcBH/tOiIdqt/47/TgEaiOrD32qbjs4tPzABUZ27iup2u28C2
BZagFv/LCSitlENMkRhThhwEqok99pv7dJnBdSlyBQdff7SAQEdaeg+2aMom/yR4Z8pm2MP1KfkP
XsU4rle99xrRROeh6uWe4Iy/rIVaIiRd3zpEqm7wb3Y32hnRJZ02jZSrHecCsWEz8kn/eeVHKZ0o
hAPZYRSpUi9Vz7LikKzotdiK8R7NdGITHwB0lpqpkutULh9VRbYDBT9db8t95sqJJ6Et2RfPwVP/
PMV2+8rvblo3OQJ+fYQMK58Kd0qse6l5ImtCuZ8mIoHFysrT6rbLrWDRcwxry+UwvqHEWjynq9jP
sIltZe2fPChQRX62yoZ3M4FGdc0eoJlIoi8u1pryedU4cuFdQ6X1+nRcP28XG5Wa17HLyu4x/Rui
YBSirKui7P0ZAZnAKbxB+fR1FiMw4mgHFB1ySb1Gaqe3pwv3FRGLtzw6Yhu/yvvYSnYPObkxfzEp
FevdRQW7MzDBhxU1fOd5fP4rReS7dv2czo3lnlxcqx70F0t0QXRbY/nv1SCE1KSnCBkHHUDIbmgl
EgSLJUkdqJh8TqXXFholPTQ2+G0y2VPLPIZE7mPVYN1Ar9rp+dJwcf8Mi1zMqQ6+/8+gpbmfR2OS
86wY4PlWB4ucVbdr099dpeteG8d3HYGmjxk8jNhuVDpFp3Q27wJ+6ODevgCYlj8H8jniDrURlTZY
mIMwvSrYxVLgsFa4bqUKlMFnw0yNJH0t8RqwCztVXTBEoFf/feEyPvke6OPY85D0BbZ/9BZOc9c4
AA3chUq7rzC5px/LFMO5Q7hUTm2DBSDLCzij1dUucrCtxZHLwlpPvrOYDkkbNSOUboH7hC+pvp3V
ExqcuPXO4ZjoidXjd4+ALNeGoBsyhsUwgAw8oVLIzeONSLo11/MiBAq+l9LSZioGiRqzujxEFVkm
WwtBm7d/mWwqWUn8ZNeE8umeIfYwVIe6DBSO3JJtsOkXlCkZCipYRxuw9qreQ1fpdPnkppwCmVGJ
pWV12ts+uZdEkNfsGmYurirnJwYlcRt/tYGWG69UYgKGKfspXyGOMePrRqCdxr9ZOMCmHUANjObf
/aSsJNspmcAksv+NO2smxY92zvuJ56nPrqxhGniunZMvu1zTJNTi3TBC+L644x3tCDzTsDu0HON4
38Vv20loguR1CcocY9eu1lT+7rXlc+Fjh/NZYF77oMCtTrFBbJ+LAGG9QARxum2+4GkGeCNHtuJG
YUjXjeMhMpCL56vX+NBuIViLg0FONktovGZ9rqYQesAZ+plc9Vt+fztOzNKtyi/KXxsnL3W2gBC5
Be2Vm2XRveQoGWfYZh5Vi8DPUADApwp/Xjzrp3YPncTztKBe6Fw+SwV8BTkbGTNe8qavSvZd+VHe
1nQwmRwdBxhLg5E2+D+lJHClRcnh7oafZU3Tc4a801gNMH8e8dTCbqGVweBMBaPziwTXy0Y7JJqR
KfMuGytx4NSbardK7R/6kWO9H6N4bYpNQxnfosX0x1ZMiq6Wkch/MTTx6G5Tp1SuWCgtm25C/ZIA
GnB6E5I+oA3fdh9rNnYjVbeNSbzL/h0WqXT8fboEJgN/yV58if+fWmf9tqlYtJj4HZ11e7ybbzCu
h2M1bJEiDbh3jjB5EemGiMHxp8IDLYqfqROdNGyy5VyO5seE2xZuMVE1K3ObfZG7gBwX4jragRaO
nbKHyZ6wzK0L1w8AebpAETJgattB3VC1xzVUI5iwNmggefrCYDzh2b3xIos5tlBMp0jh80avm+/i
JzA8qZMiGzpR8xGjGe1RyGkHA12kHb5CUEQQX0ETpDh6KyIYHL3efgiRQ58va7qzxzbzCdB/hr4C
++F/YztvGBmEe78se8dfcOVDAJTphGeAwP3D/20gxoFGwo9YrYi7yBeApUaSosaNwo2kgU3iR+VQ
xbcN+WHplCYBUGCpEYnVzZeHhHRZrOt+JwaqEhD58SH08d5Pc/Q95AHLeOYU1RecX9Wu0y0sKS2I
dZEfubWpdO5VE18xpVLyP45rXlbOLpmSD62hl6itvUyA1wGNo+nyhobkTM9TC6kEe37xKS52IdID
pwxnlendLlJ96kDFnB4fi0xnfRtLvdKwdBVeVhpovf105GPRYS07GoGOkgQE1fHhw4K9mSX0zlzu
fERnPv5dQDc3Gk7E5fXfWAfZI5f0DytAyX+WjdxgE+j+cKdJOMxFZ+oVTTw0IcbG7v0j23mlmCis
Fhcgp/rfFSwZJ3rAJJ5zvbloBSy/mIp2IZDRdEWJDqH9KHBIBFdPNw+CvlgSTgYnvtK0xK4v/+7z
sl3me29FstRUz50qeBKQeeXSwbs8o69hXa2GTx3KqOuAZb/RDuOqDqGRCiFV8W3gXI4iAFoNYkFm
ISqtOTL2GU+1X/lcIsVJoiMWStlwUtHM18iIizJYrgaM83OuVLT3Px478EEKx7C3LKHzQDgV3Ufv
T/EzaRxUAwZa3ib4GHNU43Yt3Qd4Ii1DVitlhK1pXSOagh8bHi4Cs67nWWWAlu0yIpCKU67uLWGd
zMHtg/r9Xj5fvScDgZsBum6dQEZCDp0mJYpLVyfUlxUHRvuiPCehkGik2ZAmay9RLgguuVfsuPPi
8/VFfQbWbDtyM4zQqHYBGVi9TL//7mfv1ltF/IODfnxHAzZ5TPDzf95LqQql0rOqheu88QInk91Q
8nMtl8edkfm3YL5AETZyp/YIHZlg5UZbY6xC2DcRXD54ZPq/mqOgvEvSyob12vLDX0Oaya5Yt0j1
4BrLpS1xYelVnRF8C7XKe+i6pHisiqTDTkqqQ53r1dzwZE+mnBTRHV1jBEWXPX+nKKhYkAUh2NBI
Ebc7jPS4n1+woFs8BZ0YK/b43G9B0vSmRZj87Vfavx8XeV5MiSOzFGw10lc0kO+/aEmmL32C7AT7
syzOXT/yfUXSF70FLB2MKd4Eevp446i+pdPDMS+A6veM7COv/r0jBAqYjaQReB8J5wQH/wNLStMK
tgIZ76JbNSeffc7+lPj0woEfyzT1ZsACMteVE1aL+QwcwZ+nYZUAc7PJwxJjTY4JPnfTIE/uYFVW
olQdNNJFIJKAb+ZHMFw8DLTRBDChofJvgOX1tqvBmMlvu3P97hOvuMdm4AEtB7z5ugbFNEZnYZDx
wE0JnHQEqWEOc6gpsX1YJQ6HuSJIRhb0mwVq1Xe8ooqEIup276TwucIWN6ZGstmg6I1FEYGnzuvS
FXSuxNcB3ikKj+mQIM+zAN7w6vhQXfzffevstvnmudJlEzWxriDl6FA1vpTfxmnFUQWBc84WmYiY
vI+k4e3BRU7c+N+BXGPDo7SGJC6OSrc3THeesiHw2e9Aqbpb5KxwIkPbk5hpzZQ/qi3aODnTzKAY
mhGxdNoX6u21vqWSy3/tV9E9oEljsekUVtsuC50ETE+Er+XyKYlJ8vp2/0BMIBNa2Dw6WLowcPFo
opwtMUNd2j94oWM43+V9qTkWKFVrdvj+kJeaFVUNHAWo3gsdTVf7p6fkumzzsBApicWy9vbUQwK5
kZZgfQx65yqiD8qjZdfUMkT9mTfAVerWpAAOlNe+4LTtp1Cr8sLnVH0ccSEn7uOA3i+0z08JKAPf
Cnlb65bMtfj4QqbldgWsWvas8xNHm9CO7t8z6y5F5ersWaN+WCHZ9FAncuMAzD9UHZjMfPy/u630
jLA6kYrcD50KtfJGp1Zf0CNvxcX26anNOgRA5T92aNJM5nVlYvn1xwfHZWTlLe0oDr4JCEA9wtZM
drdqgyKTpaMbY5cFiL+jmYz6rNRb/RJ7dFQ2oPaauNEbwYvKrfQUPVoJKruR+Ovc9kQvrnalJap5
SrGIPZfGMn1rJ2zNvEy4ci0NpFBgI0mGxSqibcgq8dIaqvJ8V5lu6zD+J7gi6zoA+1JHo+7OqcOx
VaGZTB+NyoJtIYCb9i7phPKjYg7XXZjH3jIYpvTBtOGrnsf213M3f6ShLZ+PRdhLJ4mqcwVg+aMV
B1hSC29eddDoC6WRC5fpxTA3ine1AfhqSUo6D7XqOi/GJKguShS5AB/a7Rp00J7ZbZ1QA4Eeeh5u
VyH9xrrfAgzFhulAuvXLOs2fZ89qguohLTjIZVwYea+Ep0NT2tWwp01IR45NOolTSDGzSDbiHCSV
2Q5PmHNnvUuQj5SF1BPydMfOQShJ/r6qpAG6pS0+9q9HStIOrjRGB/LXUpl3Vdlv9pAaMU5tNot/
QddJOabfWAobHzzmJR713p9N4ufcqsPsUX2AsGhyGw4kEuAtrIC/lQlq7azAZDr89EDJhUi62DHx
1DF67fs6aXfIUVI2idxlPXbNth2QqYJQhfjjZo9nr8sT+iZwdCQsQOOYuKTec78edqaZsA3TY2IX
yrYQlFcDy3x4O3TT1jg3OQEN0QKTPdvq2R5X4eBFMXjzUUDvqDzUJkU2Mm8iRg+WTnmSLvugh5A/
5JslYzhdpc/g6ezhTwXJbK1Cu3XScpEvtvI839IoEB2I7G7LBiWJHu2W1O6fOMlfAqJOeUxy5Yf9
tt0H6207Sp25BrSgYp15y/hvJAS1KYMsaqiyA6RxCfZ/A5IN4VyPP5blPz/qv9ZeGRhrmWkAfsyb
xBOZ497t5ZknykwTgYJLf/afima40K4ZC+8miVgMWYuBLH643Yi8EE3vL0RqqsAxvMOytc/2X0M6
oAVOOswc54a/N/jshh7ynQqNwBTPOLg+Qoh9oehoWJ1oSSgXCCtO2bAQulnJeagXDtBYO5JdwnrW
pbkHBEcF5L2wY0+0DcyxoukVjPfZ8DkAqRIMrKH8jts0aueqqyry2j9CWg/vBSYqvAAb4kXwBHIO
lfknolTyOrn5D85zbcG//gmUBSqN0KCVX2kvFr7GSpvoz3BwLTrPtdcEThTaKMTMZUkNzTCANQTg
VM08vVi/Mq5lubjz3V0/ugR7vps9gYlj2dagxYF0XxjLUk/DL6ZslGdxi9qUAeOR+38Vg1SuZmZ+
0L5LL/la3KImSM6KN5b/0bp90DB2QuVYaZJWJVEUbSVT/yS/aHjcZO/ABOY3i1vgfHjQmUHKAskI
yHL75NOCgcqKmxrssPIuUdY+E81Laotgvm3Bxv920x2FCz53RHm0Frjlw5uiw/Ske4lCoMgGIeyK
n9KEDKJnxs6lAy1Jbfu6m9dSkBt4N0TKNA7sMCVH4r8utOxEC5mFgyNNX7lg8yvbpCIwNQFqYjMl
yErxQTy0wS5AQ5nsisrGKM+vMsRv7x3Mm90fA7WLmPpyNwahJEFTZmqzADBeUz+TU5p6VqDXrREZ
dTEugPt62nRR4RSOKuZ35xQW72Gr8gmVQdsoZS9vNhTyWs0aRZlTN12xMgiUUsbLQVx58jzTIrCM
O+B3G+d4wvwLdPo+nqFKagHGhdguPpshv9j97bflENt0DrLPhhwe7zbDvHTNGsZCXly04dh6G/u9
VIXh9Y+y/N1h1aJDXMhuCSe+Iq+Yb9ZeiGoliKIi9SB8ODWpMWIFsWGh52/MGLdS6xzqHb85mjFt
HB9QCVas8Qq5/mi5zGasbhKRTNi10aiORe+XYvqSteRWUDcFiCgBqGMm4F+gIrMczs+Q7alVbfEr
vcUx50I5qhZAUDxE6DjikdEBYOJxLOct/FhYF6STFkWZelRiq08709Ej7GYMe90KD/LE2hLqqNnP
klOekR13Gy8cLBCA/mr9hVhJUAMt55vIHJ+tDWeiYWxPihepGI1R/sWV3mA2slTopH57UnTgFZlO
2O/+ZwxSvrPMbeAlfq/CZVA8YUt4OF1zY5vYKnt3mAwzA8L1dPzTyx7iWEA5EvrhPZgDjwoGxLN3
gSS/GuwjmeBQAr/dH+znQ1IbpOD8ZaoQ4nDeUQzitmFpiQCNCxyt1m+ZEnVQtD/sE5Vp5/sKCl3o
+GhL5hOtN+qmN5z3xOysK/acEnCVGOwBq3Cj7NYue1fN++ezNrDZxzHLEvEMh/qcbzxpJnJrJK9G
7KESwwRDW30Mx4VSeAwmmfViXc2ApMoMRN8s8Fa4GhjAATsucIgTkqLU43KptP8KR43xSLnnyuwN
z/uLfwUFr+/1dn3/qcZqIQSTSmdDwWjmxHhqanMbG9u6SDX2kt+FpT6R5sX7YrJD2i9omh2SocfY
Nxh8L1lnVvPmtmF9M7jpB3+WWSrp4BudU/Oam7trfp7dqJ4F0XJRUR8tCIEEfRhsD1GSwD8a5jmg
7VeN2oJPpZXpBWp8mddcslwGQuZfYYnkyL9yIcpivrXGwJnt/aDYWUVrtPWA3I5s2MunpSl06Jwm
UYz7Fa+LVllqxUFqeChIueoysE9bEnV4D44R1zJvUXa9HCsq1xlb1N7lwXTR5rh7mPqG5ptdz6m+
8/hAt26hhbju0V6joTkBZqO6IcxGHPIVlH2GEo2KwxXmAE8gIkwu4vb+Y2S6uIVr8T90fAmAt7Ol
GvpnouiSyyrCVzxUENvdFXERtaXr6ezWXrUQyO/hQxi1R3j5RLojbY5RQ0wcXPiHnsHmYDLeo/YE
GOgozjZ2JJ7GAc/t9UdT3KBfpjy/Ef3qnD710nfzKbMeLNQO1rJbBB/fp+NLwei2wVaqXl6y+8Pj
U8EA7OeBh8GKAP0NmuGVFAeGiAOJMCBNAMv81AJEfdlqAwJzTLoFsXcJSMPaIcFLYhh58g/EDDFH
F0GxgF7k04h41ccB/Oy4dhjLiezF66HAVlSKa3JTxu4fH5tEziV2NUYOxmtVyWSPmuUqNVLpwsc7
xdNCfBQWa5IY5UGyfBS4rCL6F8D3F/be8WMP/8xGr+9jPxBfvvWTahtfZe6Y8k7M5TTB7Oj/92vJ
UR+ti5R6J0qWQLNIwp8tQukcg90MoESlsMFRmf0N4/czjTBqfmm8/GTa0xviCs/rgOqpfSvmdeS8
XG7YsSpmguVePZvTUQQCccjZejlF9nM9t/pYA2a3wOU8siKtTlZ1/6g2y1KLchJJY5YjpcpMf/S2
27I/tYN+UeJbw45oHn5+UkS2HqXl29dTApk2f/ULGvAlAMs+SQ3DStjqnEm4FRUUIE0DdeHls64P
N/gxQMZui2mWYKktxd/SkTbYcu5OL5STi9tPnG+SdE8vkdErvU0VGZF+n0o8fDk8TtYIIv1SgMIE
u522qv4YYxakxbrJrjQ98M6M4grqFZiszqmXFp1QUhNtim6LEymyQ/My1voLYoqsuBfHYZ1UEo9A
t4AMsbyEX7NV6UoLBJSwEibLgjWEsjIK6W8sTXWGrCLTc08479gWkxwutUbZGedDH5NnCK1Xbgwa
CpDJBFcl1dCeJgjGSExf1MSkkeBbAgMcBlygCendYpTsge9LBdmF+1unuzagI84K5KoUC+hCIszk
bvO8sxfdYhkbCL9/B29/JeSwVUK/6RiRYX6QLHSnnTUHG9bzcBmht5bSa826ItN7VyFAII5yLQZb
GkxWAvXrkfh7w3ioDTc1JJSBqogYrD3kNM9rfZs6GaEJN1tBXSySwS3VpbT8Iwzp54vOkMF6XyLV
+kk68KPq1H+GhPpivxwgQCJk16K+eBfKkIm/sJZeJFKTo06ATBnDbXEatnmcYXeGyh1+sYh/0ptM
wlQtguK4Zt6uD+238d4MjWdKWakdGPa6wo92nyx16sx3NWnqpP6zj3aoSPrujjsCCsY32Ogo6h5E
fY8jiP16I4QDgEnuK8KZVU99al9l0MX08jiAODZDA7M2JFrteLOPGgYc4ZWqzXSbTR54UcMSA9Av
d3DKRvVLZUuk1YWh+Iw/yRAeNkBdrZzVKm6xkOthfhgJi68V4Z5QUz4aDTf0nevzibWo9bbUO9nw
2hIYRPgXiznBGzgFtqG6512y66vgKg4sWRoYU53NCaVnmO2y2Kex68Skaz0jpdamXWooIcrT9SEV
CU1SaxY5v95AQaOTWO3uf+PEKLyPmvMGUgg8SDTO+Dqi9c5QyLuVhvbCKSxPr7ZXV5NPMs45J6W0
d4mbOLp4ug3MfIXvQMMIwuGozxBeZEp1tLSSsrkznm1at9A8WoiIAai8ZnZ1ghD3QF1usMX4hDkZ
0LkycfzdK9PncRqfhY9MlkbZXEVL0/gUY5dtTYs/SvuXRf3zxEwSex1otUyc7YawEBudoq69HHH3
ECMdOmfqF1Z4sBFgPk2xv2E86qkBS6yor/03a7cMfGM7KJBPWa9/iR/jQn8e5oEb0Px1nFcmCTgE
K+C1H8CB3ifZ0d4izxCikBhYBUiHyEAQA2R13r8N48thThO7XFvrFqZbxmZ9PJETUtY1cGiEPITo
2eA4+9JN4bjWy0+P+FV8dZXYM/+8gXXhvUomWchc30aV4pTMDb3dJw/6BG6BevrcWWSSn1rr8Edb
WQzwdODmAc5ZRUfqrqv+ltlzHOj7/FQjLwZfFO6iEe6NbMkZNcIiYz6XlgGO1/0ZxkGpN4D2pk1W
lXJCIrFhYc1JVmHDTims064JdYCmojZyb1PrscUYc2rpCzvuUbvv96eOwzrBlUO2TL6PtQBkRNPY
sC9ozNsS1r9GY07t3eCDWD663ndCARj+Kxf6EXBlKvnSoOV+jP6Yo2gW/1CjoL3OsJ6TaO2FOh3o
AagQpMuTjtc8F/L2I7Qcx+miHiFBhapPy/+rywZyx6fEGv8pX4gPPxSzrcbQ4IJr7nfiGip25+7S
SzFURXIU0RdMC/6fWTm615s3Mkh1yyPK4npFcIfCxbU7emKcUoNFn/Vw5UtRvjkInZhxzoeRS/Qw
lil+p/kG9eaWKgvrlq1vmAuKoerBxRUs6cKJhYXBb3j46vMNKMaVnx23dOG3377/7v1i5Fl+1QwZ
14i7jij0s0OnNg5pmMDSXSCzBkWm0aq6+9QtGEM6HoPe0BpEs+ZWIo6ej/gSIyg5VRB6VbWWGQSO
Nj3GSe/owAnKqNhFfxgiR2yoXs8VxxF4iCGS20b3lKjAjvX3dFs5fIe8pLDFkfvFRnNIsHPYMz29
uzek5YG1dCLrH4Ry/NCeUdk9E+0hc6//RKNshRkkpQ0QMsb9H4+1EUgvR5sxxntgeX3TzE4wIndT
grZsOwTEMUyvKLJySQ9+cG3uieFD84X55nKruQSeDYSljgfaCiwqtT6oRiMGEiaL7LBhLJXbQTyU
gtzfO4jQEQH9MMD43CLeZfhtU75ysi9DBz7QNq94+Az9LkzhqKon5+BNtHVjNeN4JRu6StJOs4LB
1IbRiReCjoWgly2AABhB2nlI9wHAgwY0/vrjZphgRceSF+0VRaE0si04PpzUI6VoR2HvSIXuUcxi
HobtcLBOtneX+dexSqor7LBeqt+VR/kpBZsmlMMcyAM4Y8FrxofFQhKn+OXofeimxZi+dnECSWKM
0aseRPWAT9nRPLxwCer82ueLCBa0wip/IkDF5PX1JWPU1Gtggj5cUkC4/7FFXbKqQoSRTQakbwgd
sHa5dpKDzOw2m6Jb/lTrg2FxaISyLXQQBbjgGAMEPlk5b07i4WNzzVcs7aN1cDRaeAls2q2rGwaU
oLGeMUx3/H77EZqT6DrWIdg8Zb9q8OQYMKH1gmiRph1/z5q0aQDzcXEK1HuZtFuT5ShZ+2kPS0Py
2HvP84UBQ1cs9UctYmG+4ClKomUKdzObDbGb0Ij9Y+26wBY1jb8pNcn4IV6Qvmwt7oFDQ5t6YEXD
Zn2uNPQFCi5C0Cg2/XuV/+AHihaSke0rQ6cAjuTXNQU7gPVqB1XDtsrhOYVPF9a/z9nBl1iqN9ov
enh3BTqy7ObjzdjzthHXyx+QNnIH7jgxx3dga/32dxCVm3YcR3Y8lZs4Nh9EXI6H3OzFoW0HvGo5
JFrZKLuNEX2oU8yScxSVhe6IxfJKNlr6PMcXJSE69HyF6ZZS0KehmGvgzaitcv7SzdTr4Kfczo/w
NSjAqqj+OK3XdN0+15NdIr1EGk9ahlUItmiogLb5lBmMWu/Rzpv2CCS2HepL9TULLKNpQEgmh+6v
YhFPKK25UW8SvY/MIJCKXc/Vg0RCewhOrInBFPjL9lyp4QPwXSQSg6b/VZUc1BRSr5VjZGS4h0xi
2sQKyLKXQ9ibztyU3IFusYehq1TLPnOxC3fwAxOMGJRvzBz6YkKtnP8CKB9fapA5s1ERXNHWcEEG
73Vym5XxIUG/KCzSCghB0YNuUPEO00W/Q6SKAeMCL2rx5meEdu1w1gfEITFJT99Dw7/kexJhO/pJ
yBXlwmo31zJoWG9V4HeVnrWvbLXjU5rYoRtQ4dtydaYLAHU7esWhysl3J95JXK29iWix70XS3Uvc
ql4GOC96VqyllM403y1WbQaSRNUBuQWK+kJSjSa5Db1iQqA8OW9uaKeB6HspKqpbRqMf/wFPU0XQ
fA68evTaTBO2uzhH3J0nqG7nlhQ4xemUte0yO6ucccZABkqGoykBlKCqkKuUG1iWAb5Vh72aC30+
TVZUeBNk/Z24tjcgjY/TPeN4duO6iAZQhVzosSvHwxas0XCFcryIuRMaxssT19fPlq/DpJHCNfE0
BMxN+qmB5n241gb5mwDf2l+7E5u1sFsHgomTADteAmG9xHgTYSA61A1oyn+LHQleFGXhK+X80s+d
CJFSK/dAWRmzElYhGfLaASGHfL3ECrM1Hj01QnIZCTmJTyWbBLplCi9K8TfvwniVg34CyARxSKJU
QIHPdICDYNVu4wcEyf8KDGnW8mFJMpldB9me2K0BHKBvj+dChIN4L5yx6y9ww8vgZLZOCDboExSR
2nfhKiNXcUoCjPxVYAMBYkZmwzq27UTZ08gIjtmWPRz/nnIcZpEzx/HbG/H3GvLuN64DWDAaWV47
HUt2eA/Ri9t6zJzXqA1J3tcfsicJp8EHEtnDKA1uVxEhrLmULdcSwHMbfrQ9tGommLDuzzLMZY2D
9Q2HKRet294+stia8DnlOw+XsJBLTONHlGNZcmeffx4YjAp+1Kp2LlR/EyUZiz48dpJbXghDG5ur
Z1xoizpdkgeCj+pYK4ASqd4ChruNoE/i9bO/D8geJGzjM70CFXeJZkluo5XEdneMiATryE7aIFdg
J65jnGFRkjod/S0NEw37GgkSun1EJKEwp/J01gGwmctMPWGlrRiCUKwteGGkQSoBsZaasQVBtcyJ
wfjGVfN5+SajvPF2Pcx4m964OF3npz8YwZh9kwyfTa+WWTxanvOJuWfOXgzW7hO8Wo39yBG1i++1
wLbQSJtdGFO8bfhTJk3uVptlZR9qQZPSsyI9Qdrqmiq05Kk903f5fFwbY7s3M0M1dpK0sUC1DNJC
+CmeUU/4njTkily/XBjkAYlVA4MWMyrRBAVNWTr5D1lzKRlUSinWgpWZ74ZdJc5wcFkxM8gjdUJl
ZBCyMbqch1VmJ+C/YjYMOInx9QRZNeNd9lEj47pMx/Ddcry5kH0D3ChzRMC2YqiuXlVaX1+l+G23
UkI/r49hJALYIASIeatAj5GVy1+mcJPy+XUCwjtoJTXRx49AFnl/D1IVE6tq4tGIXCCHmA3eYo2o
qcB1SnX81SIKRoidPG2WOivwoPOCA+7W6zoJd0yK+ugSLPl5z1cjCuKoJvQ0Ds82oYnXPRfhPxLO
2iCf9ziav4mK4OB0C9vgprRUHqSs1Z+VBdyKXFOUe7fDowhggN3ruc21FstlSQH+4pH1AEsDCn8z
3YPmU3Mpmsk3RrOUHuWZLXDdRlsPpB/Rz0fzBr29IaLIZVA01+R2NYyAZCpvYaIwG3qwsbuD/4KN
JS0EzaB6ku0+y/v+LJNSRLn9+Dacbw9psHXcQwI73t1nFWOVyf9yG8ofdp5TqEVil9jHKL+nPDhf
xnH3u0SZ+lNvGJsB24QBzCIfLpFyDnZrQQIvza6+A/dXSj/yEBRo3Xe44NxH78cKw9hOfv88QcN9
0ivRqkVOmyuK/5nInRWtWBG/YqUqYmunm4/4q6HQaHn/CBAsj6xSUFErOylTRyWMayAiJGUHY5Aj
NfZ4P/TNEKbhTQv9Dy270Iri5Swx7lfDkyN5OjPbvlb4Dn9hOIKjGbmZT3UdTxx1ywAuJawU3Cpu
V79A59jyHCInWbyXkrwOjwVsid8ZhY0FDxUraxO935Udiy8HdWGEssvytYSGysVpQfl77g3P72Gm
gB29hvziJNaqTREASNMqEkSExHxDHXbXY/ECMk2tf5Kn0IN7zQzeSLXB3IbJqioI7coXyQQE2Iw8
2JELux70elTzUA3zvBpOtS0Z6YahaNi7vzX4hNE/JvMtrrs3uLjGG4YB8cgzG7UgfFYeEIHd9eOu
fm0N4G5dJz/iaaD+iZDPfaMQ13VjrohRjo2wiqSl/GdE7oQ3r14wgO2duSgxVKoaNLeKATjR2Mnr
7UtiG7cdnKwF4N3xJs+q4zIEEiQHj3taIyFXzXcG0vVcKH0VpfytT9n4dvtgX74K1erIYiIbzbzg
JvJsplzRIt1j1cNRw55nzvIAL3QjZgpSZ0MyG2fL0FM0JEvs0aRewMR2yzYpo6snqVOouZTViYhf
+IDI876tuLDaXPZ3NOPGBYn+bRevap0LmkhD51WdLLz2JzNDHaYw5qgs7UD5NK6DyZKUhvLS5XT5
Uqn672efhww6NtI4z98BsxjL9FFPaUkBgVW+S8a6hQdJP8WVVEqjxJKCltwTbAdawAtdHt/J+YQx
ziwMHrc4YkTwMtUSBR65hXnVtn0K+xOXD8xSDgSoxsWCSpGGzlN+1cKB3VyLLEsHniso0sIkBeDF
Rg37WhvZrrfmAdaEfUai7WIC2qbvYj+85ltswcCz4Q6Zj5VP6ZRZ1PfTaXlxPbDa1b4/19mT/5qM
uQHNA2O4y1pjHOeDdXCJzJWt8hRNar7WDXUFI/c2BmHNfwFv4375TThb+CnPK35mv9PJo0utw5Hm
f3RrZvcuZlCztlL6HPWu8lZETTp0N1nQ9f8hF2v0nVLoZwKTtstNmjl2jaIkkd2eR0rIo2QmRVMC
zXycQ65DONuiEy12IQKB8nKHMESNy5sW7D0p8wxX5K9i+mvHrmOKMxRAdS0Sw0gHuNwaaCSiXjq9
QVrLdaP9LMSoKk3ymXRmOr7yoXkA0uOJynxvDPzjaZr1OyBLc48TbKFkthkjlnOXCOWzOLP43E1y
RfwmWdcP2k4Kj4tuNYhhNia5wVhBlJbMKLMF2ZwK9JMhETSwTWoGDS5ck0C2q9QA+u9iRTwLBfcF
RbC+ADJu4JuxDuDRmAwsneTRKEYhTMeGyHLsnuBB5tFmmC4YXyIyq28YOon0OGtGdEJiu/g8eafq
tAA9LVLyYZmgFo+rWXufifVrsurWoKQcwcm2JJdAOrTFm8/T8LnckNiY+rV9bW/I1FdH4YQ5p1+Y
qlKcLAtdIZoxi4wbZLV+g8pJNaRIpXel1dSDnAgWSkswflMA/hfXf2UGo57VZgX/c0IbX2fiYdcQ
sljEPS29V6YkyaX7HKyXixFc5/RwCvlLlQVftGubAPSczy4ZmZPSUR/ePdKvOl5hugiuc+15YbM1
c75uX/KUql9zD1gcAc5XeTkavOzex4s1OOY/eYkxn3QTW62hLcyYlRHjpSm9yLkBrjVcPrOQILqJ
T86C6/VNQIxzlFCdjUFwJE6dAJ60/J1xQJKFbk6w7+8c7c1S9aXGugiMKbddErmT4YX5LD4ErPun
PA0iqOQ7EDvz62xceGLGJvFMPbTp3pGNzq4cr/Ld/AAXWND8CGhOuXAORCK5h4/mHegTYmXImaEC
/Flk7cTNS8f14xSxcT5scVpuykTMqdVhs4kP+Y8rVEvqg1PVOflBfBenwLr5qbwv29JdOpOinD7j
4Ls4U6GwHUYYRNVjHXn/89iZt5Hsb9Zmzc3NnM2ZkmOJAixLs5IByBK2qS/IGM0v2x7gCZ7loKYU
+snAln8lH3eu0/dM7+ozfY9HoXYSZezN/Bc3azN6dgThiZ9AjvYnwiI4PIbfp7qblWK+0wKcLH/P
5X3IR7Ww2jDmY9Wwkb8Qu80J0cp51d9kuBMNShUNC2nR6RyG7CT+WfnCMAZZjWdnsmiTopKX5t5J
DlmRkkn97uZb1qnIjD0xuFAe7asYbcYrhhhRLjWrpoyaBHYamclmRun9O5+xHs9XzOJ5U9juA4rn
01VFavIDmvwXjaFKWZcEOjH3agsF9im9pkpfoLHJn2Iqw50duIrxrpFD7lOOkl1MdMWgkFytuMU6
BmPANsR41uhG2VH9yZNnePlfGMHINuhR8ZsdjLU8GUsELvHFQxtH5+Folfk/e0dAkqPCX83Ym/Fb
k9p0I2Fe3w68WH+gRdiOGV+Bv0pmNlzKkvXowy5uMDapyIDIf5g+z14Nnbj/zsuBkKPSYkDhf0er
KAhZtpaB/D/o7GMPVdE+UwPCsSfg4sA7pOnfL2q0JfWHbNkeHJtKirc41HmlZTaofFqxK1c/ybZ2
c0kaaITXBDZHQaARAH81M7NYHlP1Whyv6wP0vYGpabHk8fjJeqQW1vG8EovwnEcOdatrx9MVePVb
4LO0u0pJ7HStD/Rl/d6UD31bP3SvkuJPvfPWBHykgYR3WfvZVR3sor3rKyf939uqx9xIRFcJyEkT
mawiduh8yyK6KyhS1S2i296cf+nuSxRCXw2LFBjWiYcTw3FPOZd8Bj0SMjFErmyWKDg/5MQvETGe
IdV6csJCDOCP/cUQKKtMqN87JLFK9uiTRz/j/DA41SxNL+ZnP27sqxbNGUCi7icX0neRn7KnuddG
muf41zCN5YcKgGX/U0N++Z6SzslsFe1qHmrEtF+vux7DEZ1Mqjf+fOngwvC+zG6IBoHsuK6wPjvF
P/Ls7eNeprB5gmPkg3DL8OUpiVMtOmDVHglVSHTme6NtE/ytEij3RHovVgdOjPXktUEUKvIC6khJ
izfyhtv+jr29aiDj0PrNzCOnBG+HvkxMgPAvEcOrSlmKciEtxIcdS82JQlIKZvwElKUw1CTttrAY
saCYCzGHJjNG73EUaHBMBHWTcBb6kWPyR5ggaJgorUGuriYSOLRoIdnxmt6dMXcJ7fp1DNgojUS7
0mGdKmx2Dw6eg4HAJwH1gp5hl8glKhe5GEwWXKnWDFWviFUZwiAhpF4pY8qoPhQ/XbrgPGykBIrM
1QswMkra4KsZ4wLgfom5M6vZPP5LC0ohYnsFUzxEt1Zfes9Jqs9dyn62v/q0xalqVvO4PTAZF+AF
lO5eMivALUlP+A9EpHuvXnfN6y6lfcdwkhN8mmRJhfWAFuYastZDg4WWNUbbBoTSue2taFR6y7m3
mFmQL83zYh1vhjzvmRDqMp4t0a5kZdgdI/nT3k5Ita+ijnSO8RmLFBjP65Nja8VXxBRN1/FM3ZCo
KlMHsXROIksmAO5KBTNo5ftBuXacNIVN/sKlYlY9DJFFQUdv5opR5DMsyopiUHlpnN2x9h1duZcI
w23OMHpGoHt4Zm/t3+4zOlcNlz7LNFG8wPobiS2Fzmoyj/vLRhF052rh/o8l/+DLikJ0MZZrXmo5
3E44eZtL+SSNtUoDgEY1q3VseDivFjpw0pd00cDoCJ+swZ0OQUttN3T/hsjoXLcJvOhGGgyk8ZeZ
djf9q2PUzQ6w7Q9wA11LKrT+HZVNcgHxGyRm1yBuSh6+O3F49sDh7CWP2HaRlHrMmrConQlPCF5/
BZG29ifCMau7wrd53b8Orfd9hZkPC2qFPg1YALMQCyl+1fibJH0r9KDmC0wMmJQ2sdlWhtBSh1NE
Bgtbs445atGFoZXZ8x2HHESNGv/EFUJw3ggZX6/2O2aaiQy0hjGf5riJGprnCZ5ooJ6UtV3+5ghm
KH7NSP/PRpoWosx60qOBn1AaaAOdMAFtEfXqn+Ma6OCbx80VJKmEXZ1Mws7ctQek7Le/CCwHuuLJ
f/frQWPu2NsqNv3Y0SgcWeJ4yQ6Nm0qBpanGJ7U8qn0aCVljF3FsSvGytIcPvJbm/JFVMJoMRPWx
4A/akfhv1ORoTByHF5D5Yp2Ay4vN1iBQM3kRBRQHQ0zjYi7+BJedAD3Gm5fNFL5ThPlk8oeXf1h3
uSl8cpb3HChP0RMeSQb6EI82/1FB4VVmlk88DMI94fACEeH4a3FaPW+t8Uw5MLx8lfyAdQMZ004w
GjwVjp6JVG2/INTWMA/Fi0JG/5O0Anb8f/3tzSeKn0iyzDaEqWEcTHlAtS5e8Qm7//eXiS1erMe4
qi7eogaC1OcCwzIxMENihYfsx6YKXs38DP2c/QLRS3DvOyi+nShnZP8QyM5Bncr4jSX9vJrfknVr
YCIjTR7UAhKGxVFvIom+AmTfDAKc6e7HmhonyyC3HNR/Rw/l1q8zuVFn8EU4o6pJwIOi5c/L5ovA
tGJH7kh6uUZqsjhPXPiuRQRctp2RU0/ZkMvUjMGedQjehHGAIiF1aa6X8r4bMDX2r8HPzm7jqr1O
bX2vdf0i8tWnhA1E5zmlneeSH6qqcrVZiE6P5CjXz29MwahhDnUQ1Rb6Ok+j52aLsdFgxQIPugDq
LWIRhW4k2R9ulkYb0fGRewe6wzIPSp5MitgRA/mBrFAyfP2uapwVwn+GPWiBBiE+6V9oaJC9EwaG
RpD/HC37BN2eJvtX1ElZA42Vvog9z20IFUzpequQJGMtgJ0B3bjNaRzBW92RIkMSTgSdYts20Q8k
aupn8nZ3rwHed4z5N+IFncPS9dpTy0azZklmI22Yhj5D7yGgee9ihNpy46Dt6GapBnL67dZ3P1+4
ao0ixF8IhfJJbjgZKTdywQ+OLsEESLXxIXTxwJPYYt73ebpiVGZ+m3KoS7d53pnrm131uDh+Lw8o
tcofA9Z8UWsl1h41PN0SnHyC/Jk/Uqa9r+L+wdk/O6W3xdbAgZVEHSDik1tN0DUQzjmAdhDEMLej
yCHSnQ4Pgj+b83wvJB614M1Fe1JJFrVefXTSRApi6hM1bKbm4MOj3SXV/jwQBQrbjoRDYBHZJZ+S
ApjJImby+YiFHO6Cc2NX1kNxkYUpMHwBGocrD7tvFOdy5BqAIU2ZcD1zkD8px3Gvwkp2bw26Tfis
k1uq5POo6rZugLXXHGCwTU6L43VVfmYsrNZ90WOAWcYn6F7YdvbYw7WjXvSzx8J4mndCDJjQDu86
W1CTm2OHqXf2EXleFMEX2mBUTjqCYDj1QVCVfMSDMoXIZyIVvgdlFsYOKYQeQfWmWqt5qa40tyYA
j7pOJzini85t+IJAMgNALRivpBqrZ8nLtmxkz6Rze1jVBIiyQE74iVLuoaPpFS/XKNYecbeTQ9bH
kVbRoH+IUDtsGIdaxiqK90w/LzSKNAYCrdxJa38f1eiasM3lmdpm77Gc/gIgiYb4SrPz8kUz/apT
pJHsl7vLDe8CGcsOxWvHr3InOe8HZtjvoO1FKZdTVfd2FYOiEvq8mcpE6sfehJk2+YfKDNj+vLop
PEA12z08jnT5c4GR01WJ+wxmqtRhpPliKb43Gqc4unBXXJKuW3Nntze3l4EePSp8QycGN+XaCbWk
k0rcD2UiVujfd7Ku5Dlu1ZCmsZXDn4d9KIhY8O1I/Z2Ob0fvXV9nMbEB7FsslCbrEsd4jdB3Rj87
Rn3HWIexoHUQRy+mhQLLJIKvyboSWdFLCEid1v1ydxqR8V0qRBeR52eFVmCd6EEOTeQ11FhSwBOK
perZ8sPFp3FOPzmVlR7mGdyPUjHl4LuUKxPpccrWZZOFhvR/hsezfwv5LkgNTTWNGvRyhDgVhkgO
VS4wNN/lC1zHPzsziuO4jGYuo9IWgrxukM3r4I5i2bHLjtfaONRbnNCFjAZ2dcH2OrBkuiWmUY+I
6ChzB+Jr/lAFRFcI1CqCoipHyNsi/5ky0dpz71vPT2zmMDFGUS695fnoGUf3/stTKvXmb9U5gY/A
exErYViyyZZ6n6J7ODWq0yQhXJHv82mfn3cpTkH/vClcqMJii0SwfVoGZ1bqegQFHBn1hJFrpbXp
U04+ZLummOyztOS7oJsimxEf3gc6kZUYruNADZc3Xg3cTT3tnD5EVZ1ACZkef500lFPBFvooThn5
ONFjcJBEYfdIJ6hDbB80N1fIvkJxMPQldovnwnwo45AwXZyv+FoM5Lbvvx1BGhfNtKcOpq15vNJn
rCM0VOy/e7plFozFWHfLqd1NbxRWLQs9TpbgMaibw4JTA9KEhQFZYAMwSq9VzSVNFGVxkGyxIIlS
xjepI5hbv7yqJpY2AEnSi954sh4qEbTvgdYRicCeIH9oeeLkC4ZkqV+DbEbyIuoLRQ0JAkuFjmbv
Y+wrWWMK95MXLJ+J399sq8PQuCt6mXGt/ZxAnMGkU7SZMIe2J5Qd3mPKLCwRyI1WwuAbcX3CPR2M
sQgCBTZfFzBM0oeiq1pfFphuzqQobEnRIN2syzAqWoPWEOCYdma60sGgksaein0MZ8QSnm7Z6mdJ
BlbdaIyCSK8IV2pIS602fEhUDQnzM69TSInjKz/uDUb0CNJowTmUvOaNEcsxrvjIsyC4yJS+rAsA
1Ch8Uc5U/7QkqbHORdRjiwzAhIJ6O7FPO+oENTJkezuWl4sk8kfBYyFInKwsHMVAOGhowVk+ujfh
kjmP5uh1Xc3jEPwBeuLL7jL1att9EfrjxCbscdaz7dbwg5quROEsyrucnHd5TEllfkSyRPgkXTBH
mPF7jKYWoOorCiE7VVd1Ol99HKtMy8zS038TKWbABsW6skZSjyqh8yzxLEO1AYMmPJXKbmJmevso
cp+gEWY/OjLRzK02XQosy6NEfVFP7ZqoOJmAzb93GOYjO8TEWvA+AM/qULca1uP0jAEHqqruecpe
uVWgYj5PBl+OfwDxrbJ7tWzQh2iTcPv8l3iZgHZTU9Z4W1xS3UljgtDxBLuHGxyqRYEhIv6hW6cj
WcVPAeC4Euw9ZTNoqVRHH5WvPE10u6GI7WVqL3hiulzz0nz7GbwL1Tw9sQ9mBGaHB21pREBd8NDQ
M6C1jUNBoIIS9yy2Y9AoISeexDmU8G/5bTWdzu4vdE7iVVS/UEcI/xpd/henTbZcXb382hIFWrr6
+iebk4BSchF6Pc+3UzhMx/QvUKucz9iYftiTEJN5CvTO9UiMYhGp2x4WqfPprOeHq/zqPKKVYMO4
OVDI8snhsIpH8eqHNdSAFcu4nk6H26vm+WIqk4aAnFnOn0iPv/Vb6N0gWxjNPKiWCyUx2qCKGeR/
73lFkG4HX9Kfx/8YkJuS/1EW5mIn1WIk3sAIzfin53pNpfiRcH28LEoLlxzxmHqVuMWieRSL5JqV
Utjc763RbJnN620M8PXurOD8tTW1Z0iJYlU7K329w/I0fY2iXmqbP2UHfEB98LR2thLHiBhmjzWr
ZEjomdDXAdizG61nkFXIEXVK0jpIDX/pDVOgS+JOMLGyfDQZav4JWcwteqVqu09JPCxaV/DsuReu
qmtStVFT9jLbhMsb5iAiYhCwKp310JWFZIkRrawArtI3b+GnhmzjCgG6Yf9Xag5E1JSQ+I9avzFG
tCQrIUpdY2BYBMeWq1H8DJmDNV4wKSAO2gQiuLetNVlfEcRptQUDvSrPTL4AW6e1i2Jh0/DVK6fL
r2vMVana1TWMfVXxJZyINweXz7Tutr5wX/Z3ZNzgws+U3IIPDu0/m07lf214dj/HkJ/Lth6SZB2W
UHLWA8WGJGuMzy5xHPPIyeJCWkIFBz38dXmeHIzanlrT2YX8UuXdfaWmvw222KSm9oUTgBrsMWtO
fjAj+tfdppqx3koUm3x1tSRsBoy8woCIOdMsP18rTIXcmUDrZxu0HkNhsS9U9W+uv7ADVvP3FUDP
sKK1nFJFUdr2aewYse1pZsYwBRJf5vpVFh/mrYwGbk4R3t6Ujn1eSPlNBrfRoT7JrMcbc1IczWXw
09gkN8x7fYjXvSE4Z+LJdjlaeFgc5GeSAijM5CzKTYTuuEiwT23Y6Cb07a8WoVEP3VUQ9ZuAimeB
xIg0uPXLPr9GlS2feccqL5VqtfViNijltcbZUXX7PhrJGnu21/NbWikwPBqtxqKdlFctqBSIfCSO
uVeKIsTIQeyaV0+NSvBcsi8BXHL0ls21/x9lcQ2u3GKtBqhmZLOtNIYAQcYdgYdnGd2BVHhtRA0m
bA6lT5k1it9pOifo1Q0l474TiYetVOZ2Rb2E35ZSigmuyt2XwEZF4c8Kc9WrUzoLRHEaRx+iavtr
Gj9hW6TGZMx8nHPx28XSbPU+qt+VLx9En6CrIysd9aOcKNLMZlfLLEPdhKG3JS19jc3OqPEr7RKi
5R9AVkLyY1NxRNk0jpuF4Mr3qZkRPBdBsAAA/FCTr9ptKtrr9Jxa67gJjVhshTwGHqKKrqPJ6QYu
VO9SIB+3icQi4s57cjbfo1Yin+6oEGTEkMZrOWTkVFoxRD0lil8ArYwRpnhUB9lsZXvHBj6/2mbs
5D19NywviwXG1KE3gufuHPGrnnl4xY+Te9OerKtV1sc2KBWkatuBfd8AcuSvmGe+GaYkANgr0dJb
aWwmjEF0krsaL7hpaYbk72eBGK7mlfeSfVULRWRU7I+0ij0RdihM87SU4/UVC4X8iDcqSe/MmS9c
q5FJ6NqxOr7ClGZx+7NkUy+hxIB7LGwV06pXdT7jbWgffGzZcTYn7DemQj9VWWsoWgNw71vy1qor
6q3mtiFtWQhKj/HCfipk4Y40JtucVbtnpr41ONFpiBkuyE/W5DfLJkncSHBRrVUluYFHMMzj6z1Y
MgTQNLbvwhJXuVD4wwh4oNDc5OzB/AU4bEwxw8FeOg2+8tU4SRE/zKrg16f+Zf7uFCMiYbHrNeo3
3lS2WXMsIoH4xcKkDV/nnO1jwZGU3CcsQaJCvjWROyrXPzoB+L5CmnS8XEPZlu5Ao5bNJ3ZktNxj
6Oz5OIuaTvXtFf71VIiIdPNNJay5B5QTIyIjXfJ1lpxoYUVWBFlpZXXfEHOaPH6PMNv5XbZbPt9U
tjlJQ+xI8pPMH7WLRpdmEa4iPH/1N5oqTE/T6qh815cab5TgBHxp1WYhtQP+vL3ARp4D6HpltGbY
rZpSSuWHd27dfLJFD035J7b2cQVJnE8kAOHZSqe8j0hm63aUHe7z32DBgqjZld8tZR2EeM9g8PZv
V9xYCbf/JSJWFvydNwkup1ju341MmWXKqAJQv5ddEns92mW1Kj641bA/X0cxhw2UrNmNT5dGaELp
2RfTQvp1v6QBnpenMNBwW/puiqva1Z9/0bcSiVIbR5iET8NN/6I6C8OLtGDOI+QLoNLDcVr1t4HX
6hpsUCSuadd1lqxp5BRKoGQ5GMk/uecOQrz76LClSCdvkQEhPgrEaJbJTRcqtv0P9IHeZEjJl2T0
HRL8g345buvmwbj7F/krhSc6jO/xSzdYjlRVJXtrgCLtvgUDxtB+E4wRdDyvgpQ72s7MpqkWIF+2
Ab0a1+ncixxIBEqArTlEXvIzF1AsVO+72H76HGgk3F+WRU7kOf/jayfsmvswrn07KRngyUQcjl0J
sPb7skc54ELe/bXocvfTi7rIrRQYkweDS9JFXDHa6mZOZHZS595t22Zws7qDu9qwmt4W0jm/biDl
qG4skKzB7TCj+DRMLbBmy5WwoiCaf1NyevUtggVebjabImBM5joqJ+bEuyXooxkDvxJB55q3KQBz
lF5RaPUdSjSQsnKTdW3ZciYqkvNRWrroA24yb7YSxFg67NAVzzBAAakzJiqaFGJvGPSFPVJ6KRkZ
bOxTlh72MQ/Ebtou6wkgFkVN5m/t2Y3sGV2Tnp2KD4Pnutl5QaAEXKzqvBp4d0JR6S+eZ1CSu7IE
FRieNxCuPUxSb6xe23J4z/SOZVCKYL5g3IGsqPkZAx1I2NrF+an7HKXhfV3QKxDDDlHNHgrXiP8a
P6kffCPpNq54f4VWhzt92tkmVollGz/szUlSSa8rz8hpLzY/oYe55uW3FwgLHVF21It9avZe3nkL
QtdGAKca7H6KLFx6KauFUK5yeDiTt0dDIoj9er2lJUnP9KgZF8V+qnMve4du+9sbcNJoRnycQDCh
2ahLUqt0ZGgsJC70VhhiBL9q001aJYC3PjmfrS+XGs+ov98/Ywq8Q2EIITRJol/s3bB565yhayI4
pm2Vu3P1ynLW3GFVtSxm7hfgNig2qTCxryof3nVt9K+2j1jm2aHaM20Nw9doP3gviu1JdNCkfEpa
sCBBZYjwiO8kWsL5VPhY1zSkdjYBpMBdouQuvZEOTCIcFAsnbYXSDm2JWJ1LmFdWgXQbMLOsT1xh
35CH8/5vodj1PsYvv+l5hszV6+oWYAwetoOpnB07FlKckIx6EmnPbSEIDaFI9ePJOwWkMN49F/+n
fzJMgTC7c2TWmu8TNfDfeQKablxip9vvgVozWMOEa0IuLS4k66oPM+jdP4WKfGaPlTg65/uhu0Vv
9keb2DB56Ne3Llqg8owj0IrgZ2kRMtwe221OplO5BtdjDH7y6sqNvP4s28oJrmOHC4pxmNt0Mnnx
4dU593K1LgEdxNpIpiUms0D3lhLnE15PheCWBw5jrfo9oZWYPoLCku5l+MAFmpfsup2dxIwgCZOR
OHHQ7Nd7RPerL51k5E+jDz8LbvbSSmmcchjmfTKEK74m9zxpPej+jtLpT0eKixgs37SlphXPjAPl
0CC5DF8uj3ylo3yUnXXCZ2Vlg2z+pDIHax4kScQTIBw99s5dhU4bjoPvepsXvJOvzyCq8DYOxIse
S7WBTga/PGzzSd6LpfXanbO390NTvPTYysu2rYo9A5oaZWgH8A2B3Nc9AMWg9mzaWgcWSPvbkfCR
r40j2kkeSusLWITuoBgVLEHAQasM38CXU7JBX61e62SwoqoeQiA3IC8UTgX1T57Lm1mwl/4EukA3
qpHEf/2h8XBWCdN4pN0mFZNS7OBuYMO+Ybuo+qSoH1f7PdpBNOta7FSFJ30WZ16lxr9UykGfOIlA
ryBUkuA4f2Yhbd1lbSuQwDCA5MXKmXO9gRaTWRXjHjZmp6EmVtkqc0x/wRu7S1ICBKPjmIZDHg1t
yoCafAzvZz5cZ4BJ+00ZbPcvxkUberkk1A4zo1nrYQkWF9xSsajcefKbf3cHk0GCmzqDEvQCgsF1
LIt8lrQ8S/u8gfovpt6KKWO6skvZYFkjq0U9Kw+UBn3yvNwPkMFZqG+u71acdXVSGDtHIJMf5rzj
R/3crz4AVO4GroOcF0iZ7jRe8uQikRLlyEaib8aNyXdIUWm8wrOhcyvSbk8hNcxhaNujs1iko/c8
RhQ0k0H3yiGNoBmypzPDAMA7uxfEflZJREtxVjdHWhVAWIPolAfOmWeTWu0ei8x7pDTrMU7FmFSH
HnNRwfoatdpQs4y536WVRcLQ3C0QCxXkFd/gCRgcyoKMlSNx5W4ZYIBlIDp+L++rFEXZXGpjqWh0
hO6NErSIefg3F+cu8AkpUT1upDlD7lp/q0jTvShhXiBk5Q8MHCYSl8MTFYv8s4x5eKuglI7BSpiv
U0VxajU8R/HAeTPYpzBAcfCMQS8IY4+rm8FSz5aap/rFts0bTv5P4kAwoyvohlxLdkWqZWfR08s/
0bqcMrt/bWjL10ijghw8WW+DTlaNWnJdYJoI7aYL/H17TghVGOP6pvHT8k4newhdALfB4njTUFat
ar2aL+OJRwGQEbuh4YXJE/iInd/lPWz2NvD2kL6yVt3Eh31Y1FbAsG7KBDPaH1rGmxWrDotx5Nfm
TGGc6238D3mPaXE3E+HAoKq3cCf9Yak7S7oGONVhskAjImSgu9h/6u3hWI4lXJ1EAFInKP5wnreU
RL42iMolbAWRvPZbZgbD+0Akj9HlxpHprNpwhsCfpNlL55Z+Mr2Mb6tXxS9VUvKt4HXPqAG8NXjW
fbOBwynjOOQ+US0I54KbjzY4tIf6NLXE+E984pGR6KQUw5Iiejxi9K3udDatGT5EEZfaMMINGQw4
FI1zMMFfvGbsEV5+7iCkR0PXYagb915JNazav9DZzcPXCPHz+RKtbD1l/wtI9v2+X0uu5ZnWEtOu
jOv2B/El/PFdMKKUaWmoXVj3vznf2MSP4iQWf8jVK7fnfgLPNXspnLrlLpjDFE7vpptDa/y2WPS7
2boEOsG9IUf6rYa0EEDWz4R6x23wcyOdnTwhHYmjdasmE3bR2L46uGdfjFFcyqvz7y1PbJzrMRZ3
LcwjRz4M9ZGHagSs3jk1TEC200TnoRU7XUi6F5IRt+bY7wLX+H4QIgm1tKrQd2IY6KBxR77R8G2v
wmFLn5Qd3KHE3bH2vXmgTiXweDDR83v2oougxwhSMz/onjjl8QsS9pEMZVTg6T/J31kcQABL5J+U
wcIn3mbpxVbwbtnfNmjfzUE4NTo8s8SW7Vdpk8R5y/jFbQWXg7NKY3+vDU6bS7PJL9u08EpFQwVH
Hkbw3WoA8Ke+xbexGFiir5oQEwlnH9f2iOjMkH8dnp2WVWGMri5HVdHJjZzsZIhwX1x6booN9XIt
8JZL8CzPQ3oBo0BdSJTi3K4Ow1fbcSaldriFn/iGKK0oWB5hb/uJZnAgIfYJZO0UAnUOnBEkBCrb
jGd+iFQG4S7dmiZo1cljtMW1+rQiK5tdAI+oMnhDFKCwYHBfYwyWXC/XLHAwWNa1E2QX3N6mwMri
YATGo37tXXjHUsQChsSzpc6vq4Ne3SKk68FrkRDja1JPbpAfF+jgvo3Ka1IFx2VfHMflFNfpmRQn
B+Vy7pfY+F/lYk3yTdBgtbgSVrxdOhKiGPm3KkUvunCVXlpIp4hT5rqcMB0AhrrsBRZv0aj0UEJM
wagod+nqw+mwm3tCBPEJPKC5HiWsxf09MMpa8WTxxvcIOFEAStQNc44rvW4Kypk00OikGpDsZ8P+
AS8JeXkBmBMavUOqkNnpmTikNokZpEEQ/5T+eue2vzN6DGD61/8ZvhgjXqInmilIiB8A08DguVUW
7oJijXEhQt/X29BPZZHoSJarHJ5Vb1YF70q4MIAhfpPiJ0/dk16mfJx7G80f/9xvIPoNg0uD5ygg
5+n1Jead0MNHkQ1HbF97Bm9yVgXhW8tpWqQp8/vazPDr2HrB9QT40gKRpTO0rwBbxoqmK5eM+8vr
Bv1Rd3JFSoPG1VnTtTyXvsJbV3lByvcAlkr//yJ3w/WFY1MzKXfCKqeIASscOSCOa3zi3nzC8+nB
m3FXnOmzQgZ+BQF3AnEr+c695MLOZ9BPGkaRXuFHKsp00zpP8R3h19admi/vRoJs+8gP+Prjk7Hn
RGPsubd9kRJSpJRWqKmj+caMKWbrAOyHuz8h/IaPVf/ePbjBq3q1mbWxvPxLcdUciVTV4i+s54Ca
eT2rVZbXv2tNIYIvaGtKvr/acanzQloxOH8VUm3IBfT5frwSh+Ry/jegn9WplPpo98yvCr5/7j5E
NfqYfRhx9IUilpkrT3esbTsAKug67iPjRGrUYrZ9HWhQKRp5kIEazpfYZpBfmUTbNaAkQWwyoGmN
wBcGeozX/Mpn2x1F95TZWU1tAFfx8DC09WyNgIAHoWgIDihjtyKyLEg1sCYQq2Kv8HSJ85OAUPiO
SLOpZlCTNYEuw4r/npjWNWlUgVYsyYYiW9u9flp2rADPbUGrDuzTXrMheQQysbJ1XhBqbeqZ+xO5
2oDB37mTULrgOyck/svjVx/i1XO748FMSbK2afb0uhGUIXHg6p3BXazWXTxieEXgTVfS0ummRWVe
gLaUhTAK+QiFVgBYmW9TsfIpPNyHx+fgPfW7kJlexrsybnDpgOYtfbiXeowD6Y1IFpqV0zAuSN8l
6zSnoxKY0I3lg1vkTLHrvg6qrA2xY55n2Rh+SyZHMdcw2h7hBXSsTLV+GNZ0rd68mRmAt1gZXzuW
bgOm5L1rSPNRhMe9cdj1/cn+GNpoJnuLReG1hrz+TkR+UglE9jRVFbyPOZwi1SvacVYOGG3b5cNq
Y6LHY6E/SqUEMp8rPkbXcOroAx6h/z3ZkCN5NxUqEnfgeEltTho0L0yXIH8AsZg9ABymMmzLYnFa
zt7A49ZRoQugJ+KDMZfOJyH4nCDyIjdaXiJ61DKDSh8qbyf65BDZhmsSWvLMsSAZfSNb1FLq7F5j
4QE0oaQ52p8ic3QuIcFIsPGCTTFWkBcXxQwHYf05rocYsNr0x5kUjH0+uF46feH3YCAeDzcFlaE0
qXVhTQFSQvm2COuSgCVWbPZvmpHrp3ObySQH4Bw2ay81atbWnY1vmLNHZfUwSVHOYoJ44Jxovlte
3V0z8gxBBsybo9IOduSTUdqFx1qNJ0EufOusyta0e6sazJ1o7Qc+wAk6Pfr9EUwLZNBzDg0Vgv7+
XBDEf31QQnpowRuaUbeoLpCkEnbS5/Mi6AkMRO0A9Kuxxyos7oR8MIA6XWyNAGqgq8hzh/82oHKi
jZm4jU7WdYbXPMhgJcKUtqR1Hc4tMfZATd3pcPv4y0nWujGGBYei3i6QTGcwOc7JC2kW6CE0zaHq
ISsfjoN08DfzXIx3XEY/C5B5l49HSxaWZdPhFgcLH93mZ2Xt01NGIZYO02I/G+Z278xYqBDg5kFR
QJLy2DL1Q2oY/QnsXCzPBIESSoitrqdxG96xqT9Vm5QE3LwM0p5mMADPeR4fbCtbAMxGowg3GUfz
qlNkwlKLlcuWu4e5RUez2qQS0BgdBdYxFPepwW1c0qz9GkLCjwRGtIT0SrAyH8dwpIjhtgodQT4p
BZezMXbOgfxfmvPelVMIQQaykFKjM0zQY8r3RDCmhgqQQlHWVNBptfwOFfIc+rmtEzZuWeAgTzaj
glqsx+8RMx8gmBcikSTIgu3UBEl1p/Rw2Vu3YIY3V9E3rBZDRNcdV3/PzxBYauqB1lxI4+vfDoSO
5GNfzyQK+gnPy6l6hotvLUkqeCDmVBPSB/v4B71cAQOHORgakKtHoZppDuKvtcvXAeeGKbj+Oi83
PpwKCNmePL8UV9Yz4Vf/oH3xtNbxPeLEGhxHADWecm4zbULS87T3sMETM1KULILp8jiki4kA1IQd
/A0Kjktravd9H7M2GEFW49yxisJk33akH8hVcZ6LugWKwv3QhISn26V6mRdiYfeWvfm/lmiy7y4a
K+bDjqDfWhI1wSbkpxv7dRfN8HavEMuBU4ACi7Kc0tBEJ1M9YevYx/pQ2RRz0KKNdsWAG7tsp7Cv
QuneVkxRKJ25YNOjQgRIijblEY5mn817ZgxgaqsutKalcsyR9fzs2unR1q+5mwW4Lq5J+G7zim6N
WNlGiMe6AvZSzbhnhaOyEoaiq3DNjhhxNN/PPzuzhYOdUH5o/Fs2xQ0IU2+z+bdf1kuVjjk65dW0
I4ofTVJz56vQCDCTD1yMAfAM0LfbgXQgfznpANkwbGMOjcUkspQF8MwOMmetXh/g3pf2S4HlPlux
PC5OqfI2za4ps3HFqvEfa7Etzy+xWkjG00YBKxJ/ule9TwmdiDw+46o4lEdZigxPySo5mfennGVN
eDylXSKu3SYs+MZnPon7KxDBRbLUBgAxo62tohQzxaSXZ9m3Rk+axqrdvWC0O6bInt+xIvJw69Rk
Qa5aVrpH6YiRqBN8X5+yiVsNTNBUrfiWTN4BUydqai3UbB6oehoaiaaxIX+acx+NBumG3Nv6x8pp
52em+1BelGmmPFO5xw1VPpbkx721kq2S2FgHKiCU4j0vQ6SOlVjnSC0Y2gFtEJGFlfIjsulQcIyl
GaP/Fs1ZfhHn4isr1grczGzuPdy2cF/JbRXmvkM/Z0IrUQGKzrjyTQRblPM4JAKnKYMtHA1dwzKc
BKgeKTdXPYFE2xovUmP8TxnjWIzgNOMrRlFkAFGFw2oXf6HlQedHbJ3CLm4NyGxWW0yfuBspqkqY
bktxHXStADVNb5waWPb0HipDbu4oZClldqUqIbAhjcqOeK1Rcj1eB6LJ1m4LBQJGumH/3UA0PlgX
CvuVnaCEfCT0Fns+XZ7HWQQsCMS4o3s82Caim/PToA2T3vv1HJ3dRWlQW++w97MTL2jCK27fCFLA
Iybm8Hb27oXP3+6bL3WIWYWz41prZlNhNd07aKTamfxbeho6kt3ljaXrA9K7+AxeROQxaB7RbQQl
WSbc02wVJcrApnCiB+LmkDYLUkC+KS8xXAhgUdww6I6N9Bi65KY6SLhqKsa8XecI3vaTG4dwxdVl
apT63g2mxzOzXAOMk/FSetypmZqpeUh3p9gxHVoLtI6Ac16wBjqrTmbh+eD/ebmD6AUrVL27ceo3
JXUmTy3pbMUn4ng3fIkhUXRpR2PHRKpQJIxPU3H3Z42WIO+EsVrXsttCcYsa6wUdIcW7huh4i/H5
/5Xz/oXrEQv3kNVAgKOue3EI6O5H1Q7RVZcsWnuyi9wEQICyo0NVDSBhJ0HYfkkuo7krRwGmDxR6
AnV9pd6CO4HerkbpqVyxJEcbiZmMiI2Jb7r95WePFkyl1TRAVRx/EeAO5adioGYawgD+2X4Mt4XB
A6yRlKvkpOZjuTZr9mCjfX1cXg2BUpI6R9OUDp6Uk2HTwHxpoWK/fupr+ay3WGI1wcwUVvBJhYSZ
72bFLS8DWD1GFnvxz0mOuioA7HyqAsmoFwYkQPhSWMpwsvhHTqotAzEBMVDZSG6dpVQKhJCRUCI/
6smSs9nMy0+ld81a+NTgcB5oKRBttcqWyzZj6jnta52iXTxuQvtGBooh2i9H21RovUex8niZhjpp
FE4FofJmk4hsNfO2Xz2Aa9fi+XVMOeGpIBO3ggFbdLofLeo7NVCKTUF0pEU1w1tI08TAxPnM4rHC
7AdMfi1aVH7CjoVAjJMbNLqn0VGxzCP4Fh+1SoHuuqMDbXz+1Qqt94VamKU+UhZa5Z4a4LogMyXX
l1yXpTfO2ONXnGcfBPu7Sih7EOm2EqTBRKBchcyS0dBCsk1O5w9fU1weu+PCAt51s/g3y4mEqETJ
fYh2X882DS0REIwIio6A2aCXmjS7tXhVt2j8F2WfeXMe0XKK6SazJreGJYP8nrb3mGdvCdTqE6EX
Mua1EoAoVFDeiw/QHts9WoKnzz7tHTC0MxtbY/9i0ERkvfI35iIkiolfkpYjNs4Y/q0EYl+8iHZf
xQjEbmsCRdfBnTWviIgb+MTWPeoJ7tFn6Gyz14QAr9FytYtzvb3ipPycWOK/YlreW3uVBt2ozACL
3jBW1RMKpgINaNWodyWxlbfswk3SqL7xLIfgCll+7t80/2JuzBNgdu8MLbNvsqRSB7FTw9JKVpjZ
Vw2tNN/3Md0Rdgd2XrpZSa7QWlaJkSYv2QsRecBNZF7ahtGbT4IyG0m571uLFyGTsHxzmBZBENmW
k2IuWHeE4hlemv8Q6RLJYxgFwFeVQ3ZpfN7KDwDzG7QYWZhQVVlANzYUOcj6vGYmHJ1bHPXrjWQd
qoqwUkRLAa5ffV9EJ1GulxDIwgSzBwiFv23eP0D6oUE4nNPRtvl3coVgXfnZxoa5fl7iCxNgp7Qz
y8BHZ5m3p1sk89mlJBtTzIMTcyIXjGGSqP4HaRPw8RTVpIWjV/Iexqj1huB5uk1IZAohCv7uZfhf
TZJ9EfofGzCEvcviOnAyDTXmqOfZmispsKkVQC4xCX7jtlTrb3u5sIWWKukKGeF0R3fTAoEXg65m
NbvOBlDzdsbM15nbpz7D6278DqKMnMo+ZmGuOhtHQLSJeEIAeSEjZTalyEOF6G2m5UZz6Hw0j8Um
kYnZtnjgTtiF4qTTUG4ZsX1+wjJ+nD4rhzO27WGr1yS0cR4U/7CWiD103hFLB1sp/8GdnwtBYUD4
iD8L9i31Z80YzJUB9hEhjVPV5ES+fhxGefIteAsX6dVkYEM5x6s49lK+q+U1uo0q1rhoqLPzuxLk
63LuixdQJtsrL0Ig6r/Qr26WfRdIWTkAdjGC1FJY4TT/1axdOuUai2X2428nn4c9u2jpco45kd1y
vQ7Csfkgywjjd18tl6eWvaOwwc3P4WURM6Y2n2+AhwpiKxz2gmc19tG5IYmwSzZxIxLwfiwLZ8tj
V8pic1Tv48N5zHewsWCz8/mF6RJ17/SLKYOqSiRfOMs/k2vMK+9O99St5ARsfXaG8nd0uv+2dHIf
D986OYoPVOpevGG2JdxV0PSb8eU+BAbBlGqKXH91HNKdDpQWIs6n7ZWhmV3QEyd1Es/3hk3J4b91
HWwSxxPZcbudtrTvbGHZx43ZOE/UhJmriamgyBL/AGT5JzzXL79oeVK5VRlouuUWuSYWciuCikWG
l4JgYqJgfOzTS1fzfCDZCXZ+D5i6x1BmatVsca6YknaC3UlZm91fb0hDtLT1o2atiKzoMaIaFBsv
mi5tcTXwKeXSKbP6Hr5rtlgRTficBiCjbkxFDICGaM/XBC3mxmwZllKX3SityBKjDJyUPI4PgGjR
nxMo9VCzK0fb9cRTQrIr/mPYdUjAMsQw6I9dthe8XPdLL8lhJTyZOhfubykVjCDoXi5/RwEijCYZ
p9sQ9dgygEoJ4ROu/DVdgbYGaWJW1aw944pTEaafIz0caszcQgVFkYclad8uCt9Yn5EdoN/HHcp1
2XY+ZVPSCAJb+//+XL+1GPXoMxdqYFA0Tx71V+RJbi8qbvNy3OUfZ4oq+wG/xXTbBzRcFjvz3C7P
CGy39EC5Ncz38/3bwOtKCanxRRH3vV5RxrJG5y8OHhwaiP1q/49m/p2K/QBpdImw5GC1d5943PA0
3extWdaUAbt28Pc5uGFPpFNeP6n/7WBP20Y8PLty9Sszt+QjbgCVmPm84tHHPUGLYr55AHVKKDVp
Nftxe4ykYTpQ15ZBgRqp4pz62AQih8/3R7OgitI/hk5cJ5O3E1s0mlvbzN4vHqlstikjP/KrD7Pq
gSZiGXiDesKgBl5QAjMtvUU0/ywwu6WbA+xSrJTdGon8kXr0uVqk10XE9IqZzJ0Fua48vLsM9qWy
pHueZr3Hai9B1YTzGAO+v/p0EkycUOgZdJn6wd3e76aCvMLh2zV7a3q4jsiCM5l0v09z1KLnVcWV
f53fDecVnRnx+NkWOTgAHQC2uJyXkTVGAf0WD7wi5Kp2xTbdVq+Ay+kn0D2pmjq/D68Yr12ayYUI
YDPj8TvPh4MY9ZQhqW4APCSIdBn7ER7aCEmvg96a59bBoAIz/PHLNBLbe6+tQpJNPzNQ0X+HxHyx
MY2RT1gNUF5R5YyDafYAaps8IKjP8xNJGNB+WPIxuXNZdRAPaU1FeD0jbHkFYS8ej9ASRmluTihM
2JbHaNiw8C+ct5thNjqzChZlFKQ9Vt+dDrEIcpIOGu4ethaVrp0hdKqrLshP3EMx6QoLFCUgFkET
vQsIxGJGreeCt659ARStIoEs7nEjQMLdmWhpHUHJZn0UZpNA5kaa4M5+cg2CMyFgPfRgON+ch63I
hmXu3/7d/CuZtv5V0cf1O67P+nCOWwuR8qt3HD0uFUkot80JQxjf4WZehLmwFTupsZZLxbAlgM1g
VQOE3obsc2bxsL9ABV3gt46iZpd88q47sPYQWCvOZEZ5BTQMQ8j+8afgUxPTY8rYEWURxoGxyFih
W3tMLEqVah04AKKfF+UsaYUTZ6JFhm1jidE9erhjk2hmcyXHbY6ykcbQwrmvD2uPVNvTZ5J3zMCd
llD+SwX3yR8ubQi9vTzXHLaGZytTw0NU+WGfgyGVusgLyw7+Wqgv39kE7+Bbxz0yBoz2LkNunvSm
WX9mak9g85/QXKXWLx7Pmjkl50Cg30ABjhdmtloHD/+cNlvifD4vWXYeU89/wAkjuc6pDDprwZE6
tofWJFFDKvRhA31Yr4e7kaWiGU7WOAC0OvHfbUZXppKHgMKX9NeTdLVYYiXclh9blmBBwvCQAzFa
D6qvXwY5KGFLkzvsZikUz1Jmwx1an8CT000Plq3ynVFSWaeEsau65wboFFLqGUvMHTnPjkgNEwN9
j/b5I0N3Ip6nuvRHQgWMnNsKedNy4yeRrVUWXCeDIU2RG89ZBJ9huCPSEao57qZFZsvmvn3jl/bP
q7FA1bRs8fE9lyOSbfe7FKWY7RNwUEYMQSmqP0QqVB8Sc13F80t/jgls7wZ6pEdU6Zl6As2psyfD
b0qpy2Dshd4ToufVypBoTV3qHF+eLhvy77o+4KFETohZXsPsNMfYQBms0eRAIXe6leyRDdh+c8K+
YcvSrP58ZdHDmYjdSOyGMVKnpo5eAJWgcFhz8KyzqJqMT5051PExjEqbRuTyTTR0XV9SenmB97F6
1vR5vDS1wFWspzDFS9/Ip1R929IF3Z9dtSxSX8MMvEMjPrI6gBHmPAejnIjuWb3EdHSFrKwn7HfB
bDpm7CV0S0HfrRQCAHqqbg8JPLlBM3yIdT7nnEnvHED+9kQZGI+2iEBdLnzIPr8WchkD3CbmheEG
ku1iPJWIqfifQL4OM9GIhw1ayMlYfvNBugTD6V2bgH1ZA8iYSlckkb65MtbD+jq97b9n0Ocdxh3f
7w9W0UXDNbIOkKsegJ3q1A/AfHaph/Z9FATSXIwh7xropmAzDzyPAoPBZZ/Rw5Dm3EbJejEGhnZV
eDr/NtaLmkX4xEJwGXnk34viyvApMqfMrClpGbRVau+eE6yE60YUAI7CH367aqOC+fvt5Ug4Rwz4
TOtdfH5Lmz+d3ubkPR/h6+GQQMSBLUEyulACVjdzwgnJZg5RX0krf+tUl6frfFrStxDHELqSz4sw
JNjYp7DKkM750EbEt66ABZVlPHbx7yi0KPaa0r5RAr8sbU1G/RB+ZvUjyT7Av0oWJj9FOGI7UjNm
60VLCSN+QgoBIffhZMOY5r49nup7W3UxjqlgoIZsIafl8rS9GGpKrcyYmdFsLwas14gZhAqs8J2F
vmYY0LO5qIHeO0zVyCRKtXrQ0/Qu7G4cP2ku+3TV3bNEjqu0owxd8qe+xsQbaGN0UKhu7uj2PAnE
3uRqhLJMCaoEVX85v2jSSRyI11gZCQjwMFeFbAhCQoMfliRozwmpZeqV6AiJqrlCSZxk6UDwaOaY
KGL9pP/deZrqC4j1CNwFySF9TKnnRg5uxy8CVZmENvHImi/eBck9EGyfMoLuPBKWj3CqNlJ3Pwtl
cHyK0478/IgNxmoTTW0ZxsmseBm8EUUVIABRsFmbGYeFD2N5sKZTA6hZfxqjCN4qx5ocl1FgH1PZ
GWJFqD4F89ybC4h+0IJ7x3VqWwmHCqyFejqd+o6MWhfbyHz4F+fNRymQFzk1AF2xBX2u+8FO181F
pY1YN4xKDZv0htO1GQp7wmzSbG5RHv40F04uUlTHtGUt+dxK93Hc+VmxVNe8WXXYpih4eWDrIJgz
yoozbtXfFn5gpB0TMGxvKGACaAS6WoKhtfCbmsGMcXqQMz0kW9KHXVk+O6CjGYj8qUUoIXiJH/ZJ
lLF8hpkffUGmBfcy+PeypPg1f03Cktm9k33ydnUtIt4V3oMAO/gHIgLbQnZSQaGxU5HDSRZuOmuX
wsegr93nDaIpoDSrnDXYFsWIFQcbE8xxSpLvTkgIS6633ajeRvFO3ckYeRoJg0qpR+Cyn0tzOTmq
9Q0bBzrC+OqrTSUZf80VN4ma4YoXAu4FS5Zt/iVtLs7P2cDzFz22K2qxsSw22H2dMs+XnxxVSXM+
DL6w9+D/4dyXmfHwsnpkG1imqZL6Bx4sjTmjPf0XXjfF0oA4uOV6kCGGXqDO/5tHgW6kBYzorsVH
VQhkTa52WJRCWlbhLH6INBT86loA1yNJby240rJ/STzMIVHwW9AlZat0FrdAQKsHk0IxsDG5cKf5
kolbsCTHg15Op56lwjf7zBsBi8ULDFoWnTwtQDD19bCieD63t8C0zJSukdr8RihUKmxDzc4U629l
dGAUpUyQVRXDAHZSXc4Avky85zGviMRJIhxMrJQzve2rs5LSMSvcPWNTCqzMVwy28JJ1Q1Ypc4EO
FiGO1qD0Lp4b7RHi+vI4RMsXSZkzoHOIOKRrvoUs8XLQXp6qfGp91uvp8DZbys/Et6psCW2JfhgD
bADu4ibF+VUtJcM035e2iy1o8hcYo4ZVCaI9D5y2yIMaohneQrmIU5B57pIuNZHbSH6eNVboNYTT
6pzkCpFECE43SOvrnsTu4IBV+wVBLlhc74ap8ZxWehrHN4sZTw6PhrnTjSahu6BejctsUos44Fnk
xV4GzRW24VzSUlB2W+8OW7Y3LcveoNG1X+qE7fJtItNV6lTv/895ETevDfp0/xb6wQhZ6cC4i6/E
PkAVj66yICTMITTXXquYzaib9mvBNEd0BG7fQfe+e4jRFfXW9M16z/5PdqZi8N8Gyez3eu+Smg+G
VDFcmnT4YxZt4xYO2sCsS2EyH+0BJzleqXExZz+8iZjK25mWsYSRx7IUX3jr9xFKqKtefKDwARpc
gqtCJoh3K98fFzTMsy5RcpTtXClopNMQEW+94C1fRsW26+FXbASVfiv+siz6qpq+Q7VzK+rcy+5r
nPRvHO1+zTUDrGj3wk0vSOB9adrErerx+c8zh+/8jNICOWLPZRN3WTFiFkO6lnY9ROUO/iyhKjqU
QXuabSMkE3Zm5zQ4zye4gBqN6hKiJuRX4vh0xUqJ5OEdRhViQ1G1ubccDjM8pxblse8B5yodXt7a
PSHG0oVLQM/jpMKEN69MjEiwjAObu/i8duohnb7tvwEj84FDHDc3RPGr72rrI+SFUxxt35jCh++z
YJomd8a/pYsbYX8YoOuvvrWv5HgpxQRk0AB+yga4Bfx+PuLu76vIvT1VWOLTJWZrVH9/UAH7BhWp
bN+2LwgfOdqxRKwtV1VSFDNxBvtn7vZuL6ipjEYwmHYP3/YpiuJoL+qCUGEGFtcDv4ixtiMeVItZ
Ga54YF2MFc+rL18YGyh7g4BHLm1SzFSZ6ZdQ1DiLn2pYqowBESCORXLnjzHipbDvChk4A0P3voq1
vk95gONtm7rSmQ0dUCPOhqFOrO29nWAvAP7ekYaN2nfGuUFVMN4XOru5st647T7ymaRGNBhHEJxT
7yzYBrYwcKxzKNQxx33hqlpWleyOr6I8j8sqKygukd5Q8H/cwsoufBJ9os7YmVu1bhGbkGtG1dO7
Xp3PhlZBL9lfb0Tz/UP0SB58wYhZfuvJUlRep7X0uzmRS/I+3Au5BcaLC+hFQtHHAXerSeFmEllt
YHNp4TRMcsh+cqPsoi9ncwRLviIDKPmFZRr/pQdFoGeZp5f77T3PcnyyAbtmLvEoGVKyxb8qkVj8
wzTzhKUzO4r85p2aipzNHWzopVSZQNlac9X14tfrFBqcWXW73iFktIIcxjiL7ugQ8rbo3ejRb7/5
2pq5U/PDSWnhCN0oE8o+FZ2lZVkOguI67dgf2ZuQ3DwFz/yp0g73n8qruWNwWfin9xy24M8e5nTU
gT1uJon7XTeXPXF8tlBYFxiTG8NhoklKqmZUQIGPIQ+1buXvdReLtBjw2oWgbka3ZcpxkLf9aRsf
npFu5pghAcsOGzIb7e2Ne7zK6rv04ee6oUsuU9ovyvRkBLllBB8sq+JjldBWE5RsOfj/tQ39cY29
8jBy/9RL2ajfBc8Y4/ZOsZHfr/Yjbtg6q1XLilbKoLkGXLuGJlY1Aer9NNiitMdPiXdSAOI9p1WO
wbtZszY8MfhiSTlpv7gs2WYtkPb2HEj1FaP2J6KHuGdndwE1gMSoXu3MXO+DKdtAkWVc9mWtUfdf
RWQjAN/TxeP5K/t1TSkLyo0RoVwf2TXVLqng9Da6o8jE82C06yuZxw1nEuWJzbExNZ8hUJRALDAT
SsKZyQdreMGzLKvo9YTZ1uDYNZERDcOD9Idbo9q2mf/Tp5Q6qZH1VnGwYKgi/F7wzI26+Dhq98I8
SuoFBtXbRyJxigSnSExKPo282abLM5yp8EvMYsWjsszL5/5UslqcZrUBHaeQ01j4Kq5z9I7NoV6A
8xmpHWYgOAfdqLQKowhLYZoYy4i6e6m565pRt6iZRcbXf/TGbNtIdBsJh089fHkR3/zt3jnTd16K
eAOAehQ+T3Y6x/55tH4bRX/7xkr8eK2BcnwoJEoDyezDZxdLCJDyb9npm36Xl+xhDlIE/JXBbWgC
SYOIONfyZdHO9ebiUTq/GVQJMrtT91HZrS8SIIS42l1PzWpEoM/c4cpB7ggSBvWEayV4nRpi1Tdg
c8g8gCowXzxFhK7xcYzop7uBpRCW7OTl+SlNkhKn6QSyTfqxsML1hqvw8orOBM+k9RVtFe8fkxyA
Ni7mP9CEo3O8jU+zLKCDdBkRtnBOoJDz2+SGfaejJAHpF9hVlJ/cNyQYHSsHcF7vxrxU7zPrw9fs
UUu3MTmqz/dG2jS2dK86EIne4ssCqzauHuk9q8pCutDaVMTa8bP9ieYnZ8sT2bGoPvMQ8q4PauSD
k257XXw9DdGt8pPF6U9B7l+D/Q8PB7lUtUN7PQX34Cer/vLytZGsrevcebjq01cOD2LviiwARLEQ
991yuimiZeLit+3EXCME81JtIrNx/qRBHFWsCYcaUqPl/GTVFraAlnMnMLI3UeE0oYQuFqtaycZw
pb2+9ng8Xb1VzLWvGnfU7SBb/ADEmL0wOrpBQ8138/04BczAQQhGbN1YilnRANzehnUaXZY08L8p
ty1dUNL/FuE1sYWonQFTdWdOSNhgDEu2BA0GBFrpPciks+MMcTbUeKFaCoU/YVFcTG/WtCFQeNry
cSTakYna0iUmf/izJGpZ7ewH2GRtNnMEKP1Y/Huizhmqvrbv80uBjFDYaa81iep2oIVJIY3be1W+
EbKrHRzXpWiza2yCnqmY1bY4zCj5oHXsDYrhZBGJCzM+j+2E7zdtBZ5U1eCyeDDwJP7+betnIcwr
dMtLlr7HGTPgjEsYsRfBN3exjf3oyon9SaGAkboQ/WpqYg6lxV5/GImwOWeCjwYaocUDyfNhBnCE
rOLRytzRukM0OsRfFe7Z2SMPO354Lmt2tgWOTh+T2lKnvhkZ5aANgxkzA44UQaUfMxxwIW5cuzJD
uUU9ydWI27RGtMi8YO/hY4JGJie+cAbSgOtcZOCLbsFszMlYN4Z5XohbDuUp9TNQNQc766g5fAb0
+EVNZhQodEBT0tjrc+6Tobqtax9qc2xnqiM9Ecrq0zP5Ur++D8miSgdBmIBtcWWOx1aCIfUKexHc
6CyvvA91yFeut8BLan1FGBvemu3jX+XuZgVM/ljTuYF3KkjbdmOz/kvah36gHo/Nm59GhUY3Pcm2
w5Pl3c7oEL+xZVELg4AU3a4dho4YVbX5GQGmWxXDE+QVFupvirvKXF2FmFqYsSBTVJjIOPVR0Cn+
LoK8HRxpoHIL1bhwMVtXwZDp5Mb5eDFvPelbHgpi6GnRoVHnlBSpFE3Ly2+dMku6i9RGwX7aXk1q
TiFSoERc+fU/HNeM7pxjOcf8oseUp26PPUf7uii79oKz7cVpcdFbN5CgBXOs7NELESyl5vnYuOUA
/3X694byuu6/phOt544vIEcYC+/NHAHLGFq3gpL5Jw3wK/BK8npGL1V0Gt+KLXJYOV5S/2Q3+/GY
rVqJ5/V4zJajneiIk5JBVktshj8Cz4Phx+3rv7ntdfmVmQJcFoNnkteZ327Z4l5WQFLOvRz2Q7Qe
384WbuMIEvhlss67ydO2BEWxjrMfSOkKBVTDAH5EN/8KiBLI8LVApusLhYxZ59cAl8AzxAxzTTxB
bMf9PvFcNZO/VOAPALtQNV0qYD+SwtKtF6xKlVLOlYecnMmGdr92YUaHhM+4YVQRMSG3EtZMSwyO
JYItCk1WuYuGUu7AZGrDmD8nnVvdperEIXDXFDt23kSvnLUohWpxsH8Pqyf8fH0PxGS5X+JQvq2Y
c1oCXucH0D5kK6Iq2xErm6xax/ylmVDmHD38ps7ZhtqMFRR1MJtGUGJH38S/nOTZ+vLAveHdRMyW
64bxLuvvaWh5iUH0EDEon1HzyCIZo6/FyZq186y9mTPg3NA/J+KXJdHEmo51NS4IR+hJciz4yIyK
ZLjtwkmo65Eevf/cy4UzrHYh9Jw1Xhno9e71xH1LxyFNMQx0c6OtyAmcgHboNzZrQsjhDAqmyzsx
fquv43nNL98m0ugEpUxlCkO2NxOTILjLgRENu/8UoyWJEyz/yG/g4Bbu0ai47JIQuHpI2RAw9WdD
zqm0Ny0+5s7S+RPaKaX5fMmiHfzUjzy+U0NvlRLKxVzGvZjzZs3MXfCGys3mi2bD4LSl4gMFms/5
x2CTP/JcegB9NQdwbLYAai09lv/9VdvrjIN3zlXDqfG+yy0OgCDgfUDSRoMEa1Lkxwk2b4+evzZx
3ebpnTCgT2QS9fV8fDszgPbFW72GpYHvci11XXsbhJy3rr8RyElCwI918RehUROdjiBqbAul/Hs+
gaN8Kc6C4B6cQUYmnfFzFXuqv+eK76NCb0H75OPKRkUmTBHD194rfanGKfUiCgoZSUM5GVKclBHS
e4MsfyhZkt99s7RLZUTMTfUXqvuxCOMlgSHk6YheIVfTm43EtONYdrl39FWVV3IBN3CS+KwSPmHa
DrGKhtUqntjK3CZvGAuEl5ZDKpAO3V8+kcREbuPsvPpaQ+9/SCfR9mYP0KqKa96QgVlOU6X7lwSE
W2sbsPMEB6vG+Mt2sycFFtrrO1OzRDOBXCVVL6cpTA9I9dPA6JuNa4AcVv73VIiBXGQd3jyAXrdm
iNcE0GzGLzJS+ck/AfgD7L2luAL8zXyr4TXenO72iKlO2qYuKiVpckygIcpoKuDxnfC3hZChcMpN
n0+JhSzFe0AqGP90xEeDpOfgPz+UBFd8C5DDnCEwnC1kTxb8c997LsjJ9zgveAIFWheHBEOoDKJQ
VelYRhxp5JjRxNxhwiE8mgU9esTwRHZDo+zXH2Hvj1vyLKfXavIZyzNbM9yxS9cBg9GkEw5h+m8o
pa5bPKaZ+IJzpT3vhKcwGicYlifT6m3xKNcG56FRTA5e4Sr+MJjgBI7TppDMlK5+WdnhwTaPO2QO
eS00ZnayZ8Aj7QPYmAJa8QfI9qaKDqNeFk/d7vDaHri7SRs7uNIsmIwgIZmM/3D0uGJUnInCIfXM
fSJXt95i1015CAI+RC+hfxfstGI2SQRnxYVTDRQrX3eVujpU5mhUe5rxsuN14Qrzo/hDNZgetRI2
sZyP4hfz1Y0PpjlFC6jo+qsTic19nieznV1PbnqWHm5+l2SITX6RtLsY+XRhVxWd59YrvL5D8gLn
2Ug/HjjDZgMIzz6gZwJ288RLXb9ZADTgJOS4pPn+jAfYxDJQaRzAgUKCEWMq87MKbw59H+xELfgo
Pk8dUyYL0vPjEIW+NpH8SyqI4sVg8jd2MifVrIspBllYAp3Zgh4Gtb1ZGSAbK7KEJ6Lk8kw1tcMg
GsmKthjFL784VxcYSlztb5QcFyLRuJuth+vvH6vKtWwYwksuuoVJmUoWT9WKZbHYiZD/Hoio2Wao
XDlu0C/rouRly1PNENanDXMgAp9Wc/SxsEf9UuvQKd605fiboLE8+KOKehaxlSBn7LioaKGO8nMw
7Ok0dGSdF1G4PMMBaICPyEV5gnm7GVrKYjsDQqVYV4cYRCJIb3+5UzNS/C0ULQ1GCL9dqTFsbd1n
yHwmNzNt3WL/d1vpxfZxTb50bZceuXaxcV+ca9Y5nks6vFsehckjPUGB8GmA+vvi1+cv5wpvHWUY
LTyJrQNZkHCNsGx+nmdGN4DYDV4Dl+Vfvqow4u4rdS4q1B5f/0SLpQela2ZRPqJc54GC/I64+9qc
Gi7RdGysnqVBosn25e8T0+jWHZasSCFHCeYFR+Is0tKOiRXWIBJrelJARgDDHJjy+T6e6Fy4ZpN3
eZoQKvbWvAsli7AHpG6KyAnV2etGXWDijutUc7A7HIzuGI5I7Ql+41KJ2Vm1x48sKx3LafIkVHCw
Ucc/9OXN/4k7mlZSJahvxDnB5RlsKF3b/TTbY6KNlLGEEO4FEJLTbwNTywLDi0tNmAXP9J8ZLRHz
v5Skjc5S6vd5IY2RLtaDz2laJJgcsaON72JqJV5VAkdPQTaYdmdtiaLx79ZHeZZ0GsH2Yrab+iF3
bcuMnRgROZ41RCdo4nVJ+hqLT15y9AkPq1jBbdiqgL+Xz4+Hl3EtFaS4sic4HMXjhgiUD5xfgxcA
lh/g814FxP8xKojUKUqmi7SExI3V6tW+SA84NexGkLC0NRxKgYLZWpnSjFGEeZ/qNP/LY6sXtLRT
dWZVYiiU+d8TymkRwI2BHzL+Y61oG4+e66hwiRJ6Pmx/sm4JL3twgGCdv5wjt711a8MoiccBc0tm
FK8cIbdJ9UTpPm34QNZHLdnTQsDVCZj0L/1TWXsLYQYMzTQA25ANYXxxdm2kC8S+cQcbhhHJjeqL
wKkiYLtkjJa2S6aDgG54Bg3Gf4DGOfHbTG/tVUTCFTMcSqNJmwb5djU6AAlzRiswSa/2XyvWFnXE
g0pmBjwYs/XhRs1IZUWblHqRrxKE1fnJlZueYSa5YUMtp7qJO1t9xA44EHZ5gRGyoe9ETMhvWMei
qrJOOyYhCLoZiHb1hkEtyrApVwdjzal4UvGdYFudBwxHOaAkXLFAuZhIHSoYyD40AdYV73lfJOHY
Ety9FaUG0qpEw/EmJw8KNYEihG/d/lFtWf2pPlxs4jriAKG8NrC3aINZ7Y96JJnpN2v4FhCe/VXn
Cjwc9BPfwV4NbH91Cf+6yS3Tw5ZqjAB8r8TbdrIe/GvQus+LYOrrVeG3ACDpd9Ng6X1l4l988fGt
bO/5u7Skyw0gR2nqWIJzVJpOLWGpOTXlt68ZvCmHJsSAfTXwIHXut0U12dCn+TDoFtvijGPB3uHH
yirZfk0ircOJ16GpucdH/RILO9abGeNj7LoFySGH51F6p3SMQbvJWkvzbHywqCut/wg8C/aDQg5V
pBb+Am8kTXxc2kRvKgw26ksRDzfiOFCo0GoCrSFQytlC34NXH7QwwOcnqd4sMr7YKMq9nUetJQVQ
bdsYveepaStycNhZTU84FmpWWbj1CyUhDU8GfkBIFxL24HF/EsjNp5P8Gut3DNLdIqmtIfpNm7dZ
SJ2EqO1oXW5xpBJG/yFgltjJ7oucQmlMAyHDeSPiv7q272GzmfFIySJB91IelMxKAXJ3gz7sycYZ
feh0kcVlGl5tAzFjVEX5F5lwZVww5WPwGbi49wDnhlw6KTZsMR8EkbkY5wDAkarU37Zmt1ihKoJr
8SByAStQdUNrRUvjn0afMwa86HNRA2o2gkNSJgO/mjUEC8NogoJ3MMPMQSseLCK0dMaIMv4r6rjj
QgpKNChB6eskml2cm2Jy3HWVNdomNn+mOvJYLaC1BBpCsbPd4Ej+DYeFb/LtgtIVEG5449U4W+Ke
OaP5+UXHL/jEImZq6R/iGinCDSVrzm7+2x7185yDO0p5MhbsuGMQGcZaWnOOtD8D1EVTfDfC3EY8
/GExTTAK4oYiqBk/NaXRSuyT6WC8IgUnjTimSddRjzvkXW1crzF6R8iCYv545A0CjzKMNUMjMqeT
y0ZqYrJNK5BOSgptNlzoC5ltEX3eIEErhcsmuBvLrz+dEtZXPMNYc1xnHNPbUH3BVaR1H8V9BSpi
sT06UIzx3OhbkKr4NTIwwweyv+MbII7bq7yIuHxQR4IctxUzvlD9GR6WpkUx5s8jzSdnqBdnYNLo
OGHp1ckegoFcuoM/E/9+/mMjWC7BfmAufTV60isESHp0NCaWxhmUpPX52mopseMEBSYBj6anALmW
01ACrhU2gXxdhJJQ4ylbMXH7hJtB3+/MVa6YZKPygVD5ZcxiJH4JPH63AZDr0IznsTwX/5T/eJVC
dzU0RvmLoteya6z2XkmHGh4nMYMTJt+xqMz3LhAojqI/hCRTTI3KD3J0Hh8iFvi2xTCGq61N7mGr
78FjkXkyv54m+cxifc9Y1ybs/VeBS6nZYx/oqg+Gfqi87Mrrd8QxMZoKLytk6W/nag5aXli3W3yF
46tbkcUH75e6ZrO5KWRviEon8ICXmjvWOoQM3D9Z3xIkQ0x4Eif4psJPw9BmkBzAAmCCXZNHFpbq
ZM+4kEFKQ3+LmbPOlEofkqKgbx0+Q+n+f03uvH8v/BKTgAz8MpwNGRHcnyrjEqhCwlUQWd5jPYiK
ArNjUTb+bN99F7qPS8jxnAdFZHIl2cIojW8cRUrSKRB9f9j8MARMKk3USgznEO93vmknspRhHHPi
yFwypTP6+o2dqveRQIxDGKwXfESUBqejhRIOtFjI0zmy7YTICvnWYgvyV9SCvrPcAk3laA7rnDmn
IsKAzUQaVKpfpXocGCAAKh7sHRDuS2Ih+mowxy322OvIF73BYLpr+TtcEZHetrc/NfV8D9b45Fx7
HxGV1cw5+beYlXnP5nVB0xN2tlV8uwVMK+90tT+5Su2KDLY8yxf68zOdwTDiOz8PYQkaUpON5ICF
lnLDpqgzpiIQElzdha44wJnBO2uehrQNZBLXPUBP0GGWGp7sIHIX9iU3dfxIangClwXR+ylVpJYk
5dSBUoDNmu/96HXtO8nP/4v/O0k2cGPb9anYk5uS3cntSREskFcVB98J0jaCKa2Yo6R8IzW9yoQB
2u2eeBK8flC7nE56e33xXKrEl+1j2csFdIhxKwcBMl/npFA2oMtMPBwXCTXBH0vrGRf3OZuscrVO
iFh1APM92StsDZa8ZZxZlnVB2ZqVylso7CefgvqF80BU07N7exwog3F1EFTL4mzvxCt7zBd8JRFh
OfAdKeygWuU49pUte5wE+wBuXWO/nE3Ul21tv2SiOlIRm+XvfgRzfTgCaVYHBc6pd1pBCoYA6hBd
x4YG4iCjtRPKJb0ffaCNlMHwXqzVlf9hBxl9+oeZ+PBkXDfOqc4R4QSDn5FDiehJMbYuHawq3Qpw
Ojw43/YP8K0Bxa53PC3f+O9uhZMCXTt/1wSfjLhkZRFjgf0WYTkWBSZ3+SURWwwCDu3XznTfTrBw
SpObH4IDgrKeaMXrAlRQ6YrJ5xQMw4TRwbUcGUQBgIR1IlFwq+MB8w+riCwS6vjKROhHVQa/QAjn
V3Sqm5v+9wg0IzGbNu4VKHhWwUamMcdXqByahbNAK+UblULHhtkrWlmUIX9pknnBZqnjXmeL6uf9
lZWTSOVc1ppO136iyMqRvcBiywRmCICc+KXpLwIUFeedZ3W270JWDuf+IE0pv3uCFy1zzXQq1lNr
++3VzKLEA5Ros+Iqw03pjRj0T1ih/kHiH37viLnUyOeptlF2/rCFrXoVww2eeIoluAductnkRKOt
a7y6pUjf885EW4R9lyhn0zrQHuL7JIStb8RT015k3X+8ad3pF00L4f+hyHxSY8JffixOrkSWWFUz
5VNHaZ5/1CzU0yN+p9MVja4IBkvnu9PRfnghm8xuZ3qYYSlB3bzYw3/bnfCLvAbgRGUUwJRWTkuF
6/FsP+mBeigcaHSQevxcKdZtB81nsxA0PC8SYPnKPZ8e5iFuj/8bFOxKLnQxfymLc4VW0NW9N4KM
kgDzSdYDDRnxR5tLXjdkZ26yht7dIEXJ6pSv3NScb3pTptZWTUzowJP1RZbYATAVeGuMDlfFQaQ+
7sqtU+xU7MoOhCetluhBBjV8w/qCdAbSTlGMRGwHL04aQzY78XBmGXhvBfkvCvwMXx3zmBfJfnqN
RcuKFhAAqjBG0pCJ506rUV8NjMfHvFeZpHRsEUMt/4uin0Lv/XX2yo0WNeuGiJRsFuMbrzKRjvZt
AGU3Ccl41fsqLKAJ0iW7GZUoPHXV25VVDkrMr5Ww9GfWOOeXdWMTAL2nvoJQHF7Q/0Wb9Mmr1/5p
AA8C+3Vb8YB0D1+Z+ETaBK/3ly9iXuJ7AydwV1bOnTDw4b27JdiFVIGUkZoMxJ4bYoCIRpOW+vpG
oc7j/eCUJtxBAl4OtK1JD0Fa7Qx3xEBgX28YhcwwXQlr0b9Wd9aCIq4MggVy2PtgnZrF9HdfjWXc
9Qpy32kt08BfBRncO2X5ZCCp3zFrtuFOozWhEs6Cs8rbRCQ/lSWoONox6pWK9r2YpaJUqNc1qBNP
/IOTQimCAxYi753/HBNn7tK9muX4484qW2KQIO/m4bLw2kKJHjErVTDzYajYsinMG23XKpN/wGnj
2GrJCT1KPg24cRkKNR/1LxrMu6xgKetRRebi1/CUai5O9TGtZdkm2YW/HKbCGtAkGSf87Vgen1eZ
DP+MhFKn736lD38K5V/JdFPTDfQlhDhnhn1xd+GqFqnrVNsoLY2zNhGlKjx6KqkX9+wqkQgHa2mB
JjQDCoBFuwbnJjRc+en9J527sIKgZNcWGKjOpPR2Eeoio3kmuRt/Bb8fuEWwVtxkbk0PL8frsvkC
biie+p9somWQu9N6vHNRRtThv0E2m6CbWMXlN7K7jnHqmHtfPIGwGNSSJAcdNbL7VLO3xcA9TXeW
DMQFYey1P3sconDIsuhyJVH1ZLcD9LR2CAQJDW16HFPSaiXDc1TkOmGfHAAubVfRHDfEBr2/L98b
hFuCXgKj6KkYavwbUsveSinI+acY4FMDjqYbCtmuhBM9CysgwnDL75RCId2AJE0ED5pC9zZcRyL8
8NEPLz1NLkjUdj4III2JElxy4daGJtbVm9MQPWd6lzcRKbprhQ0BrQQH0qWKJTkR1M5k15QHi8mN
1D8Wy5wHoEwqFjRH/1Ylq+BNzVCH08tbwVX0CWXG1uOg6ZyU8dZD/oW/MOEuf55Lbybv4PdLiQmw
S2rn1KAX2QSF1oSKaZXDmGA0RZn4jiNnETG0tox2pay1zucRpRIgo0PlHBu1NOvBzS16MBrLv41a
0spMUav/mC0MbD5BpGdLQFPyZ344EVyeofgq/BWlQrhjgSMOma/Ec9ouVQKKrRWI77ZkxiUHo11U
BkR90VAEBnAFQ0/NoEit+IGpoS5ALH/mpQx1YPX0/mOAqxewBXEj7yxKicxMHAbv3J/euoi0n0Jn
FatGhL8YPxvuSMjDJIQpw3RTqCN1L3F1JV7itLkGOpU46qwC2NO80cagrOckSQk24OvHSviWidmE
G/qmo+bKdulb+LOlqxj2BTEJ9jyaVrUGZKX/6IYpI9uPhYWW1QB/02Km1/u2xDDjlxmZsyu0HS+N
cShsvbJqoORkaAk5hjWx6zytIVYvYlmUUZct4pgS/hGLgPMnir8Zjyp0DeiisRGoRbCY2uIyqeCa
EpXQO2ApgLRfLVS1cRfiTAMlBDR857aqlzDrJCK6GiRKCK0C3p8pPaTZohlXQIgpPnX9sZbgQdTM
kWJNpDJfwSwo0TbguQHwHBKxauvM1yl/ndaaUzoH/y/DmzbIc6E5bNVHcyZXeKW0R+ihfDXER6d7
VhaJHQDPlKDur3J4z3GjibBTcjmTmbKIa91xZo2mavLc649OVqUrNxR+sj4MixrTWzpc1ZhwYabw
3k2OU5AvHWHKs1HY++/ZpHZTI/HPW7Rx7dSYmjjmOmU3ftQYg9B8HdDcjy9nLgYvSDUzo+ty+jHw
s0czd1jU07JuAz518vhPDEnRRSDma+1nIKXdlz/2hHZTCu317kEezXUO1uWbcgl8X9V9DsJsODEA
vFnrdRymMbYkcpZmttmLz2aUQGreIrMXqIngQ4qWy2oPh60kBF4dn4TXnUXt9pBdHHali3w+AOPd
oi1HYevjq72sZWa22i/jh9uFWXCLJNc4q2EzISH2qrELxqQDRhATnbtMAlSysEYOUhzvohRUoOXv
JPSUZ47VP+rxUkI8tb7jaIwQuU2nfhBsFRRCvqYSBmBrIqJl3pih3IH6wAeZ4B/JlQFz+U0A3fId
vTFCvCtKOvSBK+yf3YA+66njI2QyNPn1gikxq16SP5Y8bQlDr04e5s8FmxSIMni8fL/P22PBJ7NE
aGy/o633KU4FtSpB9l4hWpXXzwwPdA6vOne7mFcur8FtAfKSNNgq/woy6KPx+FxetzZFRDgvSAzt
mVGckesyFc8hCeI9jUa7kwTNmPJ2bU5+Hrs2sgP+NnhRhHZhJxEjsbk5wEKdeRMWbUL3qU7b4WKn
ATy2xE0NL3u3OmKW2Z2SoYeJgsM5D5Y7vQWKZeIZeSECGkqKp4ovk4BxubC1qrO35Mn5bpL/XXs1
vP7FcLlQB0gthDzMd0xg8WPHNSwPsUz9L9dow4CizPY9Encw+5PzqTlHedowfZEj7LveLxkWXCWM
mJ0Rgs+Qg0ZJpiVwdPiUVOI+TVL+CX/00nRtFfP+Pk1p0WG36fF2UOef2wQWV/mva0ASkgXww8gZ
RRLgkuHlXo0+Y44tuCrkmcI39h1k+RRCUDUDuoQvtpniwzVT6hFmTCBB4Ccy3/Ddb/uBeKl2vYv7
lwGLWPTxQavsuUaNsVJ+JZp2qwFspO07tBWRcPz1xrUOC1a47BTk02t8KTj/KYO/78cw24yqssCH
EGEztCHptEssAMHxhqQXFwcyLuXerGNGAPoi8WjV8g4mmNg/Y4oo4fbMaEKnY+5+5zbaJ+TOHx+S
B6kiG0A5008qSdjYMa1ZP1WFCXbiF/TZON1nNviPJ3+/6IqtKpLHTuPEYvYfk9F+EI/OwVNmEO7F
GJkanz+ZbQCcAyMUxGS/kHiwW5XzBPgH61gMtMsJfsN08UOAdwrZZQ9qWTpNZJ33zlt8tEgpnpnR
sKAZH61LoyyMuzoVkNhgeHktwYPhXGvCiPm6jot0stAqRhex12ivKKN58q+SdCBCEOhJibaWIsye
y8s8eXrnvfUmvEiYDH3pgZu8YaexteSUVgJt/dhGkotVgT8bnbVg14Ccm0mtE11DWNCNxwvICxYA
fthOfU2Puf2pnSUTvMh4q40q3g8Y4t7pmAUf5r83sY3TulDxcoz4yku5wvXhamjlA7P2EfTAf7SZ
0Psmt061V6506YjrdVtZlb/SPDKnxHUuIFr7iRNlSw34ollHfgAqcPZeGMdt4h36kmaAYHVAUi1T
8rEfSD69jjCbX8mKDbR8MRBiyZU+Hi2YdqA69AIegQ1s0+OGFyJ/VP3HVsNKGOVSd8n+PGmUOw2k
NvbtANNe9tLpTF5F+omdpHsvFM077GBSvm2dudCPvCV0rpKtHLttV2YL95ivy4gfZkWXQDbWY8OF
zgn+DypuuHAJ7mnWNWf7iM8JGs9fA7aZS7y0QUcO3oHJjNwU7ailhcKSTaSaMcAwXSH2WXYEjmSK
P82KLmWDQFCyebhNeRnbdSEWL4WRcdN/Nz5RQlH6gy8npn2vqxb/Og5FGyQsTYPe2UC7/Pzrg56G
pOyTu3aOpFkPggXWZZ+wmDTJQWgLcH1eyEQlMy661u9zYJrCnKjSXg0u8gcWZ5FOduqwoHHGmyG6
H3nwwXiB+sWycp88EPciDNIC3sGET5BZzpnAgnVsaqlTjfbMh5Z+iQyc/Trq8MdQt0cRA5qhN4Vh
vY422dJpy0ydkvraC3tjTQkOIVgo5N8VwMxEST39Jv+oyfocNlF8oB/kHCLRzTPscHpHS42ftcn2
YD3WYMI3T1nEcBEpa15k3PuFbWBm6zs2PrMSNhWEmzSINHvtOTpvM0bzZDe1/lbFkLwZLQd+MqGA
Q0rnRQf0N8GfFg1Y4Pct/THkujTfR6+pNGlZDuDHgXG7/ZZ5T0sOvIuNEaFUKDxsy2cuiMgT89gM
LS9qEdEvxrx1+ebqsGHo/9F4igDi1N/guxNA7wFspHwOAoYlnf4nFKuh3XnP3ooF+rvCrzRJKqVy
pnvNHDKUAM4yqIGrQIcO4aXZvm8ByqTOG5Sm+p+Nyli4BGZw01t2MGPO5QYjepveuaZ3ZmmMBoWa
suK3lFCe5nBHzJrtMJq7U8at5WQny/98POfJsZHvjq2mSqu6XcqLZFn6QOiJEo0Qhp0LJmLDULsK
trp0t0a96zptm4wvXZmkURf3EPpnIwoPvndRXSnLGcAxzFdOd1xRxYbp4E2I5kGAHDxBFxHNwMej
NkNjUMKsSY7cBJKvNWM6q2aWYjrdWgjUgHYRs1tzGam1nBS2zZue/DgvP/6RPwOMH4Kcj7MlPLr+
6OxkoHk7m1t1tZ3U6CQpSh7sAfqjSopfbOyoJ+8xEhylA0fgXXsF30wWZaDZTATHsvN4SUeLA/94
1LCxe2KpqkEznZoNoIQciglKnLbm3loQxDEPVk0lNc21CPD4rqFn6KC5lMAi2Zi+8GdvCviNz3AI
eEyoziIE1LjpdDwqWhe4A9Q7O/z5xG8Zv/LlxvNmnLsrgiC2n8W73HN3ApGIgLS+jR74Jpea5X3T
8/AZ4Pg5Kz7Rw6ueZZSQrecNzL+URktnA67eimuEorxauvL00oQ2G3mvthi9edP9bFa0uV8tkdFt
RudypEvA4sG5AgtLFfk6DgHIV9Fa4djUS1myimb0f8H6uK/yOnLogZl3AEm65gb0qTQvvT/7rsim
/0UZNkxphzyIV22bTJ6zL3ZWfIGEyGZ3uMlN8uAyncDgP1CR6qGUxOm7Avaiq3LGWVq/lk2W92hY
kJTwAObX+m8E7iyTnnc0kl73A3DaoH/ZZCAi39AHhbvhOZ4AXSVaCjjGK2RS2Bp+mYqDfQYuZL21
b3Xly0lcwcwFMAhVX31+bPAPHJkRyETFei8+YHNloXo7c7uxkWAQ/mHfARN08AbpnJFGT9wfEOFw
RqeiPEZ7lw/Bo82bkL8MAvYVxyRNMrk0YkTaRBuGmQHAlE0YmOw5QCrYYZgJnwbKwLalGrWJPGxD
TjvbEpjflceSiUyCWK2RjZn1UykCeX5tBM0HbJDXzIG9lgFD0zioCH5PzMYv8CnLAUhAImLa5rEQ
yT1e9hQJ5YzOt/umUJrN5K+un8Rn+zgHKfu33wULnZYipbL+YbYQVhyyda0oh9OmbWvSdTF3d46J
f74lgiTqNLrOtEbXuz/g7BL0WsTDYW+zulK0kz0GQTkl57GfP4RwrSzx2gF+ivVX14/94bN7xZ8A
EuAxoaea4MnKLN9yNDfsuCqvUIQ2281D79n63KXVl0sBbphLTiXGZ3B/22dnKhReo57G3Sd8js7A
OjYL2OCkWimuyGbYEW8150+/cf5lpz2TTs05HquDG1fup69Il7DJluvZayVtsdY2ll228FepPRCX
lWo+PPW+24VuzJ9Pl6Eckmlz9mlD3rIpgSAOnqtyzddwXHwi/y3Yj4KyjWXyV1fVrKu7QrtQKbsG
E+HdeKwv9AJyIov/6UGAIHcMCI8b4tfDLsxTiySX+vnsvEetAdV8bF75GVExHNtbm5UGXAonBbEx
eX7vHn2P7V3Xa9diT/Ca97/knuX2CQ2Fc27uH/atp+GQtMbjHkg3u/oT8f4BXC6kEho/Q6N+dc0+
2jnUNyCmcl3640CdUbFU4oV8tJbdRUP1bQMcQhElGQ4AYdfADIyyed5CqkXp04/Hbj3Cf0A6+krg
E7rEg6y0koojDwdg9AlNB5VjkEUDyVhlMOf1mvVtiEzPCKPwhsvLrm+VdWT4WAJesNOUgBrrQMXb
APFnKbzyEoIVEc9iAwc6wAPufDx3kYoZW9TS1/Pps5XfvLrb22X9eNc5Cnl3JATu/OcGEiwXZoVl
K0rq4rkYpi0bzQmsEg1IOois0IMfQmoYh52ufqs2XmeVMKK8YiygZkW3bgb3+Ax384RR8Z62oJlk
yG+9J51RWxPOhIY1U1gvBsqapImSwt4lyyFdMJNrw+iYw0RjzSHTPEtPjw0AUwnC9nFHkz61hdam
aV/GE4SrxU3yuuQd60N90qjuLq0Sr2xuR/AxqowFEIgbQeUWILTWbuoVwe+T9nf6v2C5Dpv5g+6X
qBwMEuiUTVNH1s722BKkQIo/HlSLZHwFiEMNGFx3KSs+eQFJn/v7cCL2VqzbPGvkWoYnOlBaUaMc
dWtKR2qugM8z2De0edGlGrXyTAk0mBU1CkEC9h8QmY/E0B4L+0QJx/Q1NzXCc4T/y5mLoMzY/bMc
08vPV4HO2+dJqdgy8JPRyoG8NQAcF7pU6JAHq3g8lrzL8wBW0rfP4iNKSbreXTN5EcJp4WHYy202
MO2flOmtDlrD12ZMc3bMvmM5REux7hfZpZ8T2X9tGm5mA+UOie/q9nQpiCGgmZ9CbYGBoH/IsNgz
9D3PWQJGs4dr7myOz1mkPzxqBbX7+moip59bdQsHQY23wmAzBdGJrSl65nq7F0ILSnr46yAUdU7L
XQWvH3P8OasHKT+tnWswZlhKnh8qbJpLZruAGigx0KKcxloCg9R+/quQZ9nH6LMoLdDIEw3Ig3Cl
EDBFDyap+fS3K9fKRiuR6/y8FoSjQIjx9ltJEYEvn0BZyidgeIZrsA51GnQkPPDQFPsawj26tUef
ocnfS8Ot/nrcCpX7bad3QESd+S/PjnuvyQoFD7v6iFXxcHoWnM/CqSf3gRBI/Ry6l1CzFxbZyg3Q
qvsWELIloZmvJqudfnjkkQrH9U9YZgftyUN4r0ENISU/C1ErSwFQH3S1Uaek4CfvMpNaT5hZ1JkT
D6JjjW3HK3PmKzGMHyYXVKO76JSNpet0BYzzFvXiQAaV7dtp2dS9FEQgOPiaqJMD9KzoB0XVULTi
6JE2ekQdXaQMnZUI+p2+QPtaGO+iZAAPuBuOiSxmUDGevZ4zjFLcS/m/gza4rld9q+BBEv/Hi0Gb
6E9zlu0CdMN/PDGPm1KZAOqzqPMiKykzJjBf12nWe+rpbThlXZt40LBC3Z2OOelCUmuLWYMoOur+
8wWFVFqsaEtq4aXoklpIRa5koh/CG5liQPsCE92/tRevsF44U472rAvL0iUHxPXfimvhKx6VSxKv
kgau0F6G6TS69dQ15qW9Im1NkWymMMo84sZQ4xJ0Ys7plHM2YjxXkON9B+rBBTq2sMsGqrFjxGX9
iU6Eappft+ah5ss2Bj5dB1hhgMs8Vi/6jgfLSXH3C73Z0LH7ScB+I7yNWb3mZ4BshYdZpESHsZPj
EnH9GR9fiwlzMh8TWaN3+PyLm1FLKeWAMENr80Fktt8DBbvLVikDFNB0Z/aO58y3O6zdot8awQz8
KRXxCy30WhMLLyODqRgpSHKSOL85AOaohJmL9nbK9e+mEbmNlI+OmsSw34DXm+lBDyCTMe84D57Y
xMCkYJ3J7W7K+fOz00SjjhpgAkElo/c5vUF1PH390IiLV/SnXa1yTr7xeoeMWJUwDXEdbJgu9Ewt
H59IUmptn+QG4nCNzdCUoXEysdo+RuOrh3sceKm3UfR7tqvJIcc6PcINoUv5x+BKp5w+YDjTbb+1
gCap6BshdlJpeaEiYf1tiigY19JTyeaNuuPzkzN+RuRvgmSAIhMFEPdOK0arwDwbJW8fTQmqa5XL
zUUGfKHLctHnuLhtC+YawndN2CoAUEhymbpsKNGGaeHSimbbdtl9dkwPrektCFT6W2IpQRWX1cZU
9GDXoP5HQS5fOKAx4lONGGsd6tZHRajSTtZeg7Ykpt8HGumkLBzXE2DzAv0D2r3HC8VVxl7WfiuI
cedFwr0E8qS2gg2pfqzAHWNFDryjUK11HhArQZzObnTA1AsBJVNbhFiue9X+qjVYZq4th6v6hGF+
U3oeJHbAnu8WUiQ5xt9jMrxxulHjFP4DYRGW0VNf9lviWDs/AoEvca0YzVXehNOCZ1YfPvb7NKxI
6rj1kpJ+QRc5jk15HnNkkUIHMUIZF5OgVh1hkl6R/lXKc6Ioc5je5P/zRJSm0EujxhpgIQVwAyaN
ByYexqK5gyn0p0X+rHMtqW7B3UX4YxyoVokerIP6AOOrBL9/O2q7bSgnIvYnzsekq8I6RUyaU561
YDajPJ/xu797VylKQ2AzVrmnFpF3TGa73BQVVrDhyaes7vyJpwfMGGbRwFbPx0TkTtJef8xWGhW9
sUNABsmxXDEzdAThjjzO/r7/81NxbiVzRFN99JiXJSxDdlDgPZHA5RyNKn9Y80mX2EZ7Pip+LOPh
LzyAaTy6XEklJ/6LaEo3PCCbX8cI6I8PRlxa4T4Gt4BQcgEnYiewSmpa0E5iZs5+NMPm8FFzlpDo
aN+f7eYvh8meX3T42L9hSPMg2lrqmi8Gy8AYRTWTrmGJfaod9QmhW2rQ2NoMQyV+lMwpR50qTHOM
fZexAoJRsG+cMERwJK+jgIMH3QgI/sCqTN01hc63NzAswI2Yla0CIG3qx9jV/N/Vwlr4LuRWu0zX
pjkaIDTAuS7bXXvRRz6CW88c/I+oyiJsldJu1gMFVZ0CvGyLrI1aQ+etkI86Ig/0Bnk+pV9amCS8
DmKuPsDXMlGA/am0ZwDJL4qFUm/3//9bj0JM5dINsEUeH9gIHF1Zib1rMrFnnsqS6IBxWG0152Oo
3xXlgvQ3dfsxp/dYP9CKo2IoO9gsK9G60F3ywTV1Y5hI17RIxC74ibacKX8/aC5WHTLTpf6/4JD4
iygTQykkm47TBlE1Ti6D3TIEQkZjXJuHY8xalsDGxAMUw7Q//+Cve4s822GuqSaXLMZ812L/5D06
M5eo+UMBnxcsGLq8UPSDe+rrg2rdh0nc6sZVIScYaBSjNzjoD3iXWPC9Gp1yTzON3jRPDtXtuxkU
mg/oS0RS2YNmUJJr/6JHVDIkAzN38DqDFH2soTgsdXDJN3FQJaqKk46AZK+qNlqfrS9TcZTrnpNX
JyaDTPrqtjDFQCOMZ7WpNABBleCXLvCyVMHigNGbA1pBFHI8DtEwPeQfsyErxhyQt00RAPG3EK4Z
eTguAfY1JqzXdzx/o2+ovTcEifo96EsOVMFGdLLSs3ctU0vR4eid33i9juaFq5Hu8BjwaSrXb6vN
IUBWI3QOuleXskaeOmYTG4F0+rRiJHn6H1qtN1BBCu9ufbByN1o7k+5shgJAWHhPr+x+MF1o/mfv
afYqmu4Kp/cFazF/KO58WbYHs4TTXlydNmbEWXbh5RG+H0hFJrI5oN3UsazorSykJCfNLwEgKUn+
E4b/CU2ivxprCbIloaIDPfIumL1P6eSa1PyVFC0+M79n6Hek32YQvhCnH5crp1tq9oK+GU/HWCnv
cSbYkv7g+rPI5dzm8jD+B7LE+6XF2ISaxCSFVgP1tt4mf5leGQ85FFtio8SN4KygfY78WdTy8sTp
DhjB09hTm47TirdJpPQBulk0t/OFbUZ6mTvu7u7a90zpxNmjIP4b5mCf2lN1FJwJ4vln/7GL5uJz
24uJfel7ioj/W2OghCPkqWkBMro08tMxUCSiW98bNp+J26nlG2DrpIufw+xXSQ2KeVTKU101G9nO
PVtSQott2VAVG/TlQKn058ABc+5tGUHPbDNMmj9MkHbIfDGFpdIocAmI7jLCsxe4o1pzWu7NOrPj
qIQu037nGx/lB4VExpeOZftwWC0sI4anfDg8Icr5qBP2H014SrUr3+b6R0LWiVmyi22MfbSHQSUG
EsyXXi7ljdN5F1ycIbgR0VSCGunPrIUFjpDL+NFoK71lQ0IbrdZ2eu5gzp352M6G2YFI5zb1tLy5
nTd3Ni7vgU7mlJMtwCLoSpQHCaosENFCShP3Y6/EW/NdPFRXypemhpCzMxY+sdu6XEpBIx8EVzYO
1iY5tRvbg+jGiGUwGczpBTVEgYqJj/Qu1KwWjqieoBhQJJWPX2IrSDHhVHwpZRlso1wCTFyBQMj1
FYXO+7FVjgVmtriVgwzXDShe7h5SB9b5uYmLXYqMmgQD3nexQhuu4gjFuBjaYbQgX8IdwTFJVCeM
dhHzIwiQbUpe1Z8VNyH7/WPDuYxN4lu+2XQaHk07x3QJUE7ry4RoNo5AFp2ieqAdHIQaUsbtR2t9
YH6+/5C4H3rdOVWoaEGA4frv4Pqyuo7ZVb3Tp37ONEAizQL8xaEcEK9I5XM39ytFxPKS6XScZsoU
4PNguu3nuHPgSIKe6mu3MMp8jbM7hXj/XGA6P2ATEDGoDsqci5HJPbeQkzfJjEINahas2Ukq9XyG
t0EJIXxRAIWAHwAYvH6MJvaM0on8l/CPQM1VS42fG20iDDFareiY9Np9CrG3x+2gox0WcH74ChWd
l43YgQZbo/6fhqF89YfIKMdsSvZIdVGAYVXRSdefg1vPHuSMFj08ZsGyKa2AP7ug1wjzDfc998SM
WwgcwZFPTk2C2HAwCTuTO5AtO+yoILbTf60U5j8CaurKhOm+FlXWBI82kO+qqq4JPtU3k7KpKaIB
B7eJ7pwZE/1ErwEuvtB1ZbMZSjxCxvrbKc3esXyMOTQcT+WWkS/XeU1lvTeT2MMGdfAp5TluHEbb
KPSItruhJRvD1hApNpCPRrjg2tXPXNYaF1ERXKYuw4tcQ3EHrMQU+0LW27wI1+urgsmgD8Sl/lrC
naDDPWpZhcprcitTtNrJf/m2BLNnMViVsTjEmrTq+BYuqTtxp4Z3HeabzvyI+2KXx//GPgejdYKi
FoeJA8FE+UjlETJnd7ZtZ0RLsHVziONFitxKrAaNDJDRjsJgrtB8MDcZJ3lucpyyD8D5H+fO9XSx
xB45UUsn/xPmopU/jKy0kt6jc+sRf/CGWkAjMCPGTplwKr6LlzKAjdNBRMSPC0NqEaIpb2VkI+YY
Ww5eUts1AdTlnDUfgEjAqiVwJ0h/BOp1dRLCheA5TXqssR+6CGyk6jCnOfRatMk+Yh1aa0AWiYFW
bebaYQA6U7pxfFROjA/xKrh9dIdMJzs8ZjT+2OQRKeJrKZur5+dpdfdSNBvXBdTlTn7vbl56y0Qa
8t+Q/6+h//EXvMZsdCLL8PdK5bxoUtNe1L1KZPWPax7r6ZZ/+OrN20uCrr5gw86shlShMmoyK60o
WAe5mlTdilCapIZdfubY3Rb2/BD7pulZOsdcGUqsllwdk1Ubvf+ATuh8y4ruUzqjE9WrxHYGmPNH
9mpChm6A1SKfVdaNdiw71M1VGcOGCuNmSLuU4gh/VmoEhRCIXqm6aYU2qsGfejCPGf7njgOTnszQ
CSJiAuGqOdXtOsemHMzNeaCXLiLFRf8aVRHqtQTwZoy31sKpWHKepims3cXKUWWeLas9AH/fULzR
0aBg8fKp0wpzKwRmu7YKsZdnqjeUq5AzB6GX6nJvS/WvotJ1tdXfTwjQTtjwscev0FWU9EpZcQxH
LMtZt+mgloaoUTQwugP8ZpgcK1ab+uPLxCynBHl4WdJYXEQabRLLdOc26VKk1GD8tsh7/Ln3Xc1z
mAkV7xYkarRzQIQZ8l8QfB/JOwQy/6Ioc3peaGCy6ALx7QYXWOgu789RNo3vH39BH1X0AZuiiSkS
/OzqHnuep/QkjFqFySCik8PyJuhIWwEP6E2f6NPT4vvp0DaQssNlHppGI00bR8VBjqytNuw2uuuR
6dYEZRSoWR4fnP6s5NV8sI2xmEh+bPTArNJPWxZOTHiLti7clqC9Thckh9bATE3Fbi08VcjhbhLj
A7iUJ/XKqZ9fKlRVqt7S+XiIIrm+zD3RWn18MELC7AUUeQZnQf7Q4UD4oq5dlyHxSa7hzpvG1GZM
ZaWt++ubbWaDEi6rlHPlyQkidCE/rgE7+Izdr1chK+9Gf6XbygmGfz38bV2DL9Un/oraRD29sIuU
49VQ+wYaUdiTqXvfOz6mnMltx/f7eHCMhLfS2G4ssHbN0Lq17vtfHsB7o8JITu6ECtK0otn1gZoP
VSrqMp7GnKJtAcqyrJ81Judtn9qV1MNzjjFU3Nivt1TJwoXBj6xeNvp5a6SWxga3lowbPCDGNBWL
ChXHDgmb1c5m2kDHb91KHkZF6JrhfmDawT9U6C5vTK0tUvr696n/spdTqigWzDH3Qi+zQrp7sCE4
EiUQwaLpzFbgfHvzz4afskpaRmvMiZtiefTDH7AX90m72kkpSf/6D281srS8Vb+nXH6riGDtL70O
NnCJEK7jRxE9Mydy4yjHFzfjz2M0W4VHCwXpiEF9tDKO9NNUV6zLiPRpUAolXplvIVKChaqk5COY
lLfP1YQ8J70ewZ+ECeNoQs1ErbTPKZe7OADvsi2G+hyy1DE/T3O2lKBu8bQTGFrx4tzvZ9zxvmE7
7NeCGv/uRIYsZkWc81Ecv6cF+JJndrumlW4aZM/trySO0/RWn3EvIpa0bD4NzoxWA0d1l0b92fOF
J7sgsKbU5Zmvpo1Wfonx3D6BaI7sopndWo0LITZp7HAPVAZQoAC5DZESXGO0uciER68Vnl24fO0g
fiOCjluiop50QdeyVKyW0WYf7KrjkfA1mL47IfT/ydNjyO0pJVpw61AOhkTh6CdJWkHX/p/Orpvz
XAbf/qCpoFcz5AP19vfVuv6HoHg5FMDXnGPM2NkBtKdYimsDLiUoV+5Mpc0+82oaxWh4BbmBGnT7
P9k/qI4XCr+D4Q5/AejxOSFxMTL0fU+fLk2PcDtF1lu4FSPqaWPGUtMBSKlP5Hg6u80evJrxzpza
lS8e7Pl4dUtiLajVEAoywKrjLa+otaUNY/MHML8hM1D6S/RZ0pv2ijFdJ9htjciffFrlAiIwU91W
N8Rb4k1E3pG0RsHb9ruRAfWvNPbQYOcLMM0YsDqp8fMfuSdRkHRerVK7N6M8Bu1lXmNgbLTxJ246
2Qqyo/91OWtyU/OPs+iXdLTqGgfju8OXis5vKHjXJMA1DIPXxt2elMiWicLaqTyTY7ZRBtY5hbdQ
XG8q6R/Lg/oNxFkMqQEzDBDP5H/Gu+Vyj20+Q3khYl1T/dT+PabBT7X3/mDahkI55ZIRm+0cXhVG
Pnp5SlZHIh2KQAmzRfUqzmtf0XM7OHDv0nuN7NY0WJczCFLnPaPxDk8HrKgstpna34tazL8ZAQp9
yeThussAvHNGGxN2yUlijzVPejl9vkLYLnUPyGlKwGM5mkcFn/EJeG+DW6YMI2m8kgt/5F3Jo16k
EOl4kaA+YUqNVJztUm5xagr1fX9t5tVDV4eWLsEKSRN5dAwugy7uFX7g0joazDWu0GOQnLnpmSGf
2WPkO2+xlMd5g+MiEJUiVw2lFGP0K6JbjuqcyCxBxBjS3PqWxQAI/RjIlWJYQjHXeLXNlf3nerl4
H0V1EoPXKoFon6lI5DOhPaTNZIy4UP9r/AXF6f12+sQ2Q/ADN0Z3pTCH7DT4seTmvw2jMr93KSxN
8sqYoKn03CjgbKMg/aZZX1g0qLsul/Z4z4so4PxkVqIyqdt1BFX4NsXy5BKxUOtomEOkf8gxf9N4
LwHGEVvWWkJKq/KrsM2bT5nJRDNokEVcxZrYy8c5tPkB9g4wJd+8ppJlo8L0+JxfKsrkP7cnDT2B
Bzl/Wi0rTM7Uo7To11bxoRrn+hj425WYYohvzgRYZ1dhPVWNBSxRzNbwEgU8vw1bwsEPEOzcQ6MA
CD8SHYkxLwcl11daVuw5nr9336H4Kzt6UR9nDYCGgLQ5O9lcRVzyTL3GW44++qE/Ft4Jpg36zCx5
la1sKbzef/IhCPdYyN+wJfzBeOUMnN2dvxhTSzhxczSC3HvShno6oQFV6/gTpMnqUqKFiLw0x94r
FQ9kuHr4JN5E37mhEfm77ubUe285zE1UO+ekDI2NdDe2o/Smm9fPNT8qyI/8TedEZ8DlrxhLlr1P
BWrOI5nSffc5h3qmI7VpQlwEw6iE08qJ7dHrvF3kXme9qh59szald11vnV71oNz8j2Imu7y5XLek
+EoY3fLCbPgjkNyJcUNmn4RnxRABteHV83Oxv6oY3qQdU0rrNhUQypDI4MELZPECzcGEqA7fwjxA
rQwvVqyeW4/7oYv2a1bYsesBBAGcw47EkcyEAH3bdY3PvCy6rOd5+jivK7LwhRmgQ+ZlkXvHrsnB
+m+2PG+LHSI0MwLpo2nnRZAoO0wJkUGySWYNEHTJV5Ws0zerGjsrf7DQdSHYKc9BxdCSg1iu3dVe
aYPMiR0WUx/EvtLv9ObGwoyZYyInTMfAHEoO9GGsxYzAwGzkCLBuNeuDphX8zfFPcredlG3wVIgy
rsmOjCBGDX2zt02H3q1R62rC9flMgYEs2WFItyrQ+xeACZEuQuYungUq2fpGnoUqW5bKF2cmSuLQ
lRDLqydqins/SRb/zE4UY8Vn24TQusBa8mgdFptWReCDtQ5msSM47cPkDqQblthzsyamiNk9imOs
tNcFd+a97axEJ+4H3/wA3vQlLHXtFlsM+QkcmrPfh9xZjPu8H8/vnXeaKKzJlbMxBeSJOk7i/440
RfNl1W+AYS2PUN21jCYmFvVpQlO78WaiiUuPOoJOTkENoRdy+zg7T88OS1NKibrzdCvXX4dMl+P5
dF7CNNLz5Ovohpw8OV3w5TlqsdqUu3kj1D1VlUM2WgM8oh6IIw5jYjp4DXtsauoFeHo/IU8EHlVQ
Kxn8q/oqf+UZjJ8c/oYmMzbr/ma5xr6ebx1mhYvVcWW4qb9xrMx12gXPzJmxonmo8CEkX/vN3x3B
8Bj+XnOWCm+xzT57CicUHIJ0T56+TijbOqNYgXXV2GvqAsruesyuNuyEYISQQFQpoCTlKZe72NPi
PDqZF2RR3FigwbP+hYF3fEfft2LohwMEnVn7I3Ebld+b1rVI15ecBb3J1j0W1h9Ssju4mMtVegUl
ivGts7nJSOMGphA9Rj6XlvnsTpgXVPC4KlSDMQ9pT7uue/sd0jN5JIkaRSzSddRVgp1L/K2qTFWt
2GwopkM0TVZs62mpdxi6lOTPbsH9xnYqkhY88mUAK00gIAlqk4M5MoktfJsMACGvH+e1GY/m2+Zb
fwUTqViYkOK99mZ44cYLkCFhCRgjyy8td5iNGy/SP/ONR783z+ePsPV7hQb39x801igDU2uv1hwz
F2pKLp8itIz2MKvnjimdNg+u2rMsJbEvIp5Jdjh0AiENPD5vxSy64GZibaftrXOMzO6NLVwIvd5a
8u4UEk6B4oIAFkD6/HIY2kItpCvWA5Cq8S1wyX35eBwBI4wXkT9MIMp18tRXgnIa/+xlE//OnEh9
eniwQ1AQUc7f4nyg7Np61YO4HnbDbUoWHpgFvqAhKPFuJpLWTiigPK4YF4bNJoUVWS8Kkx057r2N
fxT0+eFzvKyHflh8C2srE0btlxjVLxr8ZeRRdWbC/9WwmPuV0OuuA+h51y3RvsD+wzI5cBFZZ0g0
jawJybO3kk4I6fLvfxCokx97uw7wnKpjdIUjY2AHPolEtaT7Kl0hMJTIT29dFpjVf9MpCPTktDRI
MaKu+oFDQujdQsyEwlF7f36JNC3WNSIjZSuDEgT0KwmNj4x+ydfaoFoYwxRQrC6/LsRQjJ+v2HAx
etSXv+WTVGc9G6XTDdJoc8P89WKGnxDDCLHvI73RmlI2wDEpcNB/frKAcyirNBzSDK1WB3qfEK3e
atPtxPqV2lwfXDjl83sCD67IcQKGNwkiFeic76qqBj1OZxkyRF1EcyKFAdZMUdEL1BI3JcZI51um
uMp7bQwT6R0iQTO8tRJ/kCV49BIRhMHsE2Nb05T5Fd2S1Q1tVnbMiFVwUVy4h58/1rpMK0ruWqVD
4fZIuZlFviKxjx/l1IRrVBMAyQbxehuii4uMFT6LXeSuAvtH+Fyp6Jb1ehHTK7huBBeaw1WgUK6H
oPpL2Mhscxnx9+vsOvUztQUtXFyORh4NaDypQvQCcjVU5YYrKDbCLJQIXuBnBfXtr5YPMGhnXv6v
pUxcmjO4gJSroNanNKWiknI9vQ4sTbsJtuXZ5++nS0XD6NaK6ocFZf7iDgAZ7RwvaGoHiuxW9UgC
4KxftmgylidpQWaomzLQ9kSc8mHAO7JA2h/S6GDiN8h7aBqRlxLaAIk68Zz3LJdv8j5Y6LxOx+rR
W/j5vRmHEqq3cf9rdbsdEpaappeeLuhSbD41LYSmDhBobky7tbx0OxPBszz6KjFZOxRpLGrk7/bq
6XXif0/GO4mCB8h9rfhSGav+DxRxZEO596TJ/2UTxe7aj754qY4xfBLOPzGTOSIoW/2IBXWE5xqL
AHfF/eo2uBVuJP78hs1YjklsCrOeM22Fq3ezilIX5LA9iuVRm6DANSXkZQFCJLf/wYhM5h/b8FmM
i8RSFxZOZjji3DiwCQNZb3r3llFUIT4uYyIECC1OQFiqFUo5bOSTdMGiiQT8EE34qd1ieye1QAjN
dARCFGlctf7F8JMZYLvtphLhTLGZYlEzIycdTrl0cfAiTkvNxLVDgsM4RwX6DO/G9we1T9WJ3cUR
G9nPvoqTE1AKB1u6foMcsDtvxeBH6C6eHjatjoxBbkxgyhw6+Zh/Je+3v66Wl+XvFEAt/HpBkUsu
SbA3YIDgK6sYF+0ibCudoBYPLudTMyxf2yP+86asZi0poCKVqAf7PU3EoPvSfa40XerjytACpJ47
Jb8AOyMDW4cL9pB/Egqaka4+0x4xPgpIfMwzTMZW1cTEFAVQ3vhZtFfKwDarzWtfr0WoR/RSa9zj
IUYFzmQuOQTdCH5pYIQRY2QsjhUKPqRJ5SQOHW8idv/ENWCFpubVXodChJNO+EFJN+LVhAPWo6Yo
ezBV7DjK4gRm8Hn3ecxkrczM4tOCHv//ozwCnM4JGzEBBpUZQ3tcTyUYPqPUh5rsv7ZPJRRoaBZd
XWxZ+JxzKkhEFb6U7XbjgXthnugYDHuEdsAhtlgBjPrBAzi+LgW22xJYP07qIPvcWL0MLJ/oYr6g
/jP8iNfmG+1euDV5zr2SuiC3zFtTg+v+eEvyeIb6Aw5EhsxhLEoI3t9MVj185MynLyOKq7jn5szW
NfYMivns08Cg/VGAU25rC76x1xKRWMSfRtNRXVt96LljBcLd8gvV1uyUaXAJrn5syjsLtJhEb0u3
3jxH/aVimu49hv8xRoo+kixI0edaCkAiVvJLMjWDjpgSU5mYOgHIAn+a/jqHRVxXr71ZrPBm8h2j
11ISzhZT5G0iVvm2YsT8cuZasARPtNzClPFwDWjege1//M5x/uSzB37NKHOmXpkR5wUDbfxBBtk4
4XmBvKc1VQ7w45B+wrRAhvm0s2fqUrAx9H6pMZa/aEj3obtA6HyN1GwBo6XxAu6kg2LFTnu+Lhmu
J4hoEt/V2nH+VsWtxeSFSze+OmgPSlJqGRdukjZ6P7TMBzVquQnigR1gelDgHY5Jh4FjibBtItb+
LrEnoxfqZKtbyL1I6iLPvaTqZTXpkZFfoNlFp5KqbqM55Ncuw9Af68fKDNpxt0UqYhDCoR3q8QOi
t3YLXQme8jatBNQlQe7QM1n3kwnEZuXtmgefK5mx78N218vCuJaMUyd6Mn8zliyScfSfihUNMpeL
9NVsQpWw06iF6N25RuyYq0VQBbWrnn1lLT0+rDmpibsEkP5PZ51WulqIwzkChHTrcHJ8lUmg0SxY
Ae6XVGBKX9DH2fEuyvx/X8rq90CRhpXP1VDpT9XhcosrDYtH0Q+o0tvUI/+YeQnllP2+fNGjp7S8
TOvcDJP9GihNUDVT4mQfG6sRhAW73ynwLiTYzLIAFdyZfrDVAQZu4yNtnHatXYIngc8F4/LwdRIq
2KaosF0n5otMc7aL1TyB0InTykASJkWp60PP/5rAolUxeMmb0Yi9NdBRTScwVgoVhwvgxi1oinEU
6p3jRcrHbCfwTlo5Lgwoug3LHYXuCjQCzpZiNs2VXJ7AJyRKMfPCczX9uTCnxYCajpXWKeI9QWVu
s0xmmbi+V0U4y0DSsS6klc9rGSQW3RQcTvcAjZxQwKh4r4lxUL4LsHdxUIY7tI7yA8V8TORPzGNN
8wgA1yqq7WLUY3NmunXvPbvvwhLthIi/s/MGWF42hz/ZoYL0HhEWQ18kYli3ry62s1k5uyRGLzWe
1/YQEQQOvUlfvtgSQhphgX3Qn7+oFDseVyKYPglZExSJVF4TjuD0mmMJK1mGYAa0gIJF8HpgUwXR
HfugM8HlEqL5Z6aHsEJ+FLYx4qKih7j6FWw/iT0Y+MGe81trDyNlxgKgh5aIK3RXWK8CLKMgHalR
UnYjJ318x7bQW7Ir2CG/Oaigjr2Eb+ezyWX1ouzTaaZm7t1metR8DrhFrvqxt8OsdI181hpoxpgC
9dyhpbS1HHAr2NfXvf/N4KRIZmgz3uZlfobQ4cjuPI5SSamNPYy91Doaa2hMlPrfxLK4di9yFt+U
bCf3Oxq4OR7Ym5OWgbRfVodFSqtjW2y1gslpBGco6VjB4ij9gOL3261tmO+Ty++45pbZ/hoH67vy
3OtxRGBo50AD4evr75ofz+LDwaTdCOPe2vt2oJR1C20oF1bdvLBUC3Cvkbj7pr4fRqX3RfbSRVIM
Z1fTIoJaTI7MKp0IsjZ85Gb36vS7ZKXjrwWno9wfLvFf4mPKAsbFKIrlLxdWSXqEC38DfEGsl0/f
vjvD9kM7Q859geiCkeeB0gh6EchhlgEcTLEQF/XYSG6VjNMgZcmJuyjA5OJLSR1xTD170uS2hKcV
Zf994mIiys+DTrDCk9RUMOpZzLLa6oddv38uZ9dtugde4UoSK79ZucH/RD0TAQPbcKvx9mJtTQqV
/K7LHjauKPKKNYCrfiaT0KiAbDM/IhOSVCxTs+eTfujR4E5oLSOkao5k+rZtJOhEJFDU+7CmOLLV
EER7JcdGSivljm9GLsG50xLxhByDxncYMr3EeAa3KuQWKxclIOhiocO4EdOpJLOlRpSvdjdDEDBE
KbA+01LkGsjWey/+XKCJOMvoscFKoiGa1hLuVmjOrSgM+dfc817waKfThbOS0xCLs9EJ49l2L0pg
V/bpPZIEyD+KRp8m7UYw3QKv+um/+FsF++xGz7d+tA+DfYUTxf/YAghWMJUbRz9UQsAzOC5Eu6bt
YfDpd7TwSjeSln4z5r/1klzRfwwtlglhXevOwOItlCWcq9aGdZU3505NLraRg5g9G8W/CGm1Hoza
TpsLkSzIk2BsfEC8ru5K3B/gK8g/REgOP7FcBe3Y+qYaKYSrIBUunOsmkh+MANLLXUdV7fjdBpYk
TVCMQXxJGz9RE3IukTlK9sf3FY4RP3pVe2dZuvytySjkQAq5uX1wVbO19FV9DW078TEF94OHKLHj
HmGWBVdu7wp21OrY30MubkkEPINDdZ6gsc5mmgPZEdGXHSK15ArZALOmMgJ/QrIyD4ZgfzWpHTkX
5j8/xUaPm6jF7XwtUlocoi8PPksrfXrQSUiS5uwosaRSy1G7OW8wkEvjZmPU8DVc76MyXh4aANsW
BS4EJi7c2ZP2g6XP5exB0zo0o2C5gQi/Ne24e5FfsTUJ1SpN3+IEg0mnTTNdvPtlhDG29KccgC40
f5gLgp01tT4IgV6nQ5FdC4pNOmdCJTgxPLRnHzjV3B+0t6nd9QO5SoBc3ib/THD9IhOMiPC7oKQN
X/u5aGjQfOoOu8AjBu0mieS178SIGR/sCUeS3rhGTdRI6+gg+HdBpLjk/GG+aqtrY9KYgepH5e0u
5td6xgQVAivMofr4GZhpO2Lwrj/pf1fle8MPeotMrgMIHpzL56LYbQf4SRCxEJTedrxJzJSY2mwr
VuSJinhRryFwOh4LdY4PpvfqEHHyEx6sQWaNABBCIFTNXBiHRiDoe0CgXX7F64W6B0/Hg4kFkh/j
TPNM8Vh6mDJp/QgEwbbOdMeganPmoDNafFl+7UbHIcpV2zj3jCzeKDETrEQk0IoN1Vb6GdQK6c/U
jHzkn06i0ay8ohPFeu7rpbFVVWH3QLcwugs/3QgfkTrnauEOI4iNut3djktFx09NaSyUOT4iCYb7
J+NyDZiomv4S4H/mSsC/z64itQllLopn1mNdg4ZDznDEL/GTYe/DBHnqJtGHX6YUr1+nIHVAmxf+
3YGNLpgR79gDdPaVyZGmbAebmOo9Bky2MaImyao/ccKP3TUQQwUiEvHnBjrSbP5MvbgCbaai6dhN
egaX85TzFlU3hnB6KRD+32ko4Kwkx6ih+ICI1f4XiBDfdC2uBsmCRKAH7ooIAGkFDQfPRmyjaoMF
QQZehOSAQovHmDHukgYjIQna4Be8ISn6B98+UG1+OsFV+d7BCCDODkNd2oHcXFAk/6AVw8XC9OA1
lVbRJjkYGJHlWIfpjF33K8ZObQgsF8IGGM2Cmw3yZ9idVbGsUZ9SV5cNOFTswvfMNzHk3TOUMu3d
wlMC0w77V/f4
`protect end_protected
